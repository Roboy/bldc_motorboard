// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 21:12:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    inout PIN_6;
    inout PIN_5;
    inout PIN_4;
    output PIN_3;
    output PIN_24;
    output PIN_23;
    output PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    inout PIN_12;
    inout PIN_11;
    inout PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__51094;
    wire N__51093;
    wire N__51092;
    wire N__51085;
    wire N__51084;
    wire N__51083;
    wire N__51076;
    wire N__51075;
    wire N__51074;
    wire N__51067;
    wire N__51066;
    wire N__51065;
    wire N__51058;
    wire N__51057;
    wire N__51056;
    wire N__51049;
    wire N__51048;
    wire N__51047;
    wire N__51040;
    wire N__51039;
    wire N__51038;
    wire N__51031;
    wire N__51030;
    wire N__51029;
    wire N__51022;
    wire N__51021;
    wire N__51020;
    wire N__51013;
    wire N__51012;
    wire N__51011;
    wire N__51004;
    wire N__51003;
    wire N__51002;
    wire N__50995;
    wire N__50994;
    wire N__50993;
    wire N__50986;
    wire N__50985;
    wire N__50984;
    wire N__50977;
    wire N__50976;
    wire N__50975;
    wire N__50968;
    wire N__50967;
    wire N__50966;
    wire N__50949;
    wire N__50946;
    wire N__50945;
    wire N__50942;
    wire N__50939;
    wire N__50936;
    wire N__50933;
    wire N__50928;
    wire N__50925;
    wire N__50924;
    wire N__50923;
    wire N__50918;
    wire N__50915;
    wire N__50914;
    wire N__50911;
    wire N__50910;
    wire N__50905;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50886;
    wire N__50885;
    wire N__50882;
    wire N__50881;
    wire N__50878;
    wire N__50875;
    wire N__50872;
    wire N__50871;
    wire N__50870;
    wire N__50869;
    wire N__50868;
    wire N__50865;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50851;
    wire N__50848;
    wire N__50839;
    wire N__50832;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50822;
    wire N__50821;
    wire N__50820;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50798;
    wire N__50793;
    wire N__50790;
    wire N__50789;
    wire N__50786;
    wire N__50779;
    wire N__50776;
    wire N__50773;
    wire N__50770;
    wire N__50763;
    wire N__50760;
    wire N__50757;
    wire N__50756;
    wire N__50753;
    wire N__50750;
    wire N__50747;
    wire N__50744;
    wire N__50743;
    wire N__50742;
    wire N__50739;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50712;
    wire N__50711;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50703;
    wire N__50702;
    wire N__50699;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50676;
    wire N__50673;
    wire N__50672;
    wire N__50671;
    wire N__50668;
    wire N__50665;
    wire N__50664;
    wire N__50661;
    wire N__50656;
    wire N__50655;
    wire N__50652;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50625;
    wire N__50622;
    wire N__50621;
    wire N__50620;
    wire N__50617;
    wire N__50614;
    wire N__50613;
    wire N__50610;
    wire N__50607;
    wire N__50604;
    wire N__50601;
    wire N__50594;
    wire N__50589;
    wire N__50586;
    wire N__50585;
    wire N__50582;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50572;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50560;
    wire N__50553;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50540;
    wire N__50537;
    wire N__50534;
    wire N__50529;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50506;
    wire N__50505;
    wire N__50504;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50489;
    wire N__50484;
    wire N__50475;
    wire N__50474;
    wire N__50473;
    wire N__50470;
    wire N__50469;
    wire N__50468;
    wire N__50467;
    wire N__50466;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50455;
    wire N__50454;
    wire N__50453;
    wire N__50452;
    wire N__50451;
    wire N__50450;
    wire N__50449;
    wire N__50448;
    wire N__50447;
    wire N__50446;
    wire N__50445;
    wire N__50444;
    wire N__50441;
    wire N__50438;
    wire N__50437;
    wire N__50436;
    wire N__50435;
    wire N__50434;
    wire N__50433;
    wire N__50432;
    wire N__50431;
    wire N__50430;
    wire N__50429;
    wire N__50428;
    wire N__50427;
    wire N__50426;
    wire N__50425;
    wire N__50424;
    wire N__50423;
    wire N__50420;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50400;
    wire N__50399;
    wire N__50398;
    wire N__50395;
    wire N__50392;
    wire N__50389;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50364;
    wire N__50361;
    wire N__50360;
    wire N__50359;
    wire N__50358;
    wire N__50357;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50351;
    wire N__50350;
    wire N__50345;
    wire N__50342;
    wire N__50339;
    wire N__50336;
    wire N__50327;
    wire N__50324;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50313;
    wire N__50310;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50294;
    wire N__50291;
    wire N__50288;
    wire N__50285;
    wire N__50282;
    wire N__50277;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50247;
    wire N__50246;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50229;
    wire N__50226;
    wire N__50219;
    wire N__50216;
    wire N__50201;
    wire N__50198;
    wire N__50195;
    wire N__50188;
    wire N__50179;
    wire N__50170;
    wire N__50165;
    wire N__50152;
    wire N__50151;
    wire N__50150;
    wire N__50149;
    wire N__50148;
    wire N__50147;
    wire N__50146;
    wire N__50145;
    wire N__50144;
    wire N__50143;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50136;
    wire N__50135;
    wire N__50134;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50130;
    wire N__50129;
    wire N__50128;
    wire N__50127;
    wire N__50126;
    wire N__50125;
    wire N__50124;
    wire N__50123;
    wire N__50122;
    wire N__50121;
    wire N__50120;
    wire N__50119;
    wire N__50118;
    wire N__50115;
    wire N__50112;
    wire N__50109;
    wire N__50100;
    wire N__50091;
    wire N__50076;
    wire N__50059;
    wire N__50048;
    wire N__50033;
    wire N__50018;
    wire N__50001;
    wire N__49988;
    wire N__49973;
    wire N__49958;
    wire N__49945;
    wire N__49914;
    wire N__49911;
    wire N__49908;
    wire N__49907;
    wire N__49904;
    wire N__49901;
    wire N__49898;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49871;
    wire N__49870;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49864;
    wire N__49863;
    wire N__49862;
    wire N__49861;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49857;
    wire N__49856;
    wire N__49855;
    wire N__49854;
    wire N__49853;
    wire N__49852;
    wire N__49851;
    wire N__49850;
    wire N__49849;
    wire N__49848;
    wire N__49847;
    wire N__49846;
    wire N__49845;
    wire N__49844;
    wire N__49843;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49823;
    wire N__49822;
    wire N__49821;
    wire N__49820;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49813;
    wire N__49812;
    wire N__49811;
    wire N__49810;
    wire N__49809;
    wire N__49808;
    wire N__49807;
    wire N__49806;
    wire N__49805;
    wire N__49804;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49800;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49794;
    wire N__49793;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49788;
    wire N__49787;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49764;
    wire N__49763;
    wire N__49762;
    wire N__49761;
    wire N__49760;
    wire N__49759;
    wire N__49758;
    wire N__49757;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49748;
    wire N__49747;
    wire N__49746;
    wire N__49745;
    wire N__49744;
    wire N__49743;
    wire N__49742;
    wire N__49741;
    wire N__49740;
    wire N__49739;
    wire N__49738;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49731;
    wire N__49730;
    wire N__49729;
    wire N__49728;
    wire N__49727;
    wire N__49726;
    wire N__49725;
    wire N__49724;
    wire N__49723;
    wire N__49722;
    wire N__49721;
    wire N__49720;
    wire N__49719;
    wire N__49718;
    wire N__49717;
    wire N__49716;
    wire N__49715;
    wire N__49714;
    wire N__49713;
    wire N__49712;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49706;
    wire N__49705;
    wire N__49704;
    wire N__49703;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49694;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49689;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49683;
    wire N__49682;
    wire N__49681;
    wire N__49680;
    wire N__49679;
    wire N__49678;
    wire N__49677;
    wire N__49676;
    wire N__49675;
    wire N__49674;
    wire N__49673;
    wire N__49672;
    wire N__49671;
    wire N__49670;
    wire N__49669;
    wire N__49668;
    wire N__49667;
    wire N__49666;
    wire N__49665;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49131;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49100;
    wire N__49099;
    wire N__49098;
    wire N__49097;
    wire N__49096;
    wire N__49095;
    wire N__49094;
    wire N__49087;
    wire N__49080;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49071;
    wire N__49064;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49050;
    wire N__49049;
    wire N__49048;
    wire N__49047;
    wire N__49046;
    wire N__49045;
    wire N__49042;
    wire N__49035;
    wire N__49028;
    wire N__49027;
    wire N__49022;
    wire N__49015;
    wire N__49008;
    wire N__49005;
    wire N__49002;
    wire N__48999;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48987;
    wire N__48986;
    wire N__48979;
    wire N__48976;
    wire N__48969;
    wire N__48966;
    wire N__48961;
    wire N__48954;
    wire N__48951;
    wire N__48950;
    wire N__48949;
    wire N__48948;
    wire N__48947;
    wire N__48944;
    wire N__48941;
    wire N__48938;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48928;
    wire N__48927;
    wire N__48926;
    wire N__48925;
    wire N__48924;
    wire N__48923;
    wire N__48918;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48891;
    wire N__48888;
    wire N__48883;
    wire N__48880;
    wire N__48875;
    wire N__48872;
    wire N__48867;
    wire N__48864;
    wire N__48857;
    wire N__48852;
    wire N__48849;
    wire N__48840;
    wire N__48837;
    wire N__48834;
    wire N__48831;
    wire N__48828;
    wire N__48825;
    wire N__48824;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48816;
    wire N__48813;
    wire N__48812;
    wire N__48811;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48796;
    wire N__48793;
    wire N__48790;
    wire N__48787;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48774;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48737;
    wire N__48734;
    wire N__48731;
    wire N__48726;
    wire N__48717;
    wire N__48714;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48704;
    wire N__48703;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48697;
    wire N__48696;
    wire N__48695;
    wire N__48694;
    wire N__48693;
    wire N__48692;
    wire N__48691;
    wire N__48690;
    wire N__48689;
    wire N__48688;
    wire N__48687;
    wire N__48686;
    wire N__48685;
    wire N__48684;
    wire N__48683;
    wire N__48682;
    wire N__48681;
    wire N__48680;
    wire N__48679;
    wire N__48678;
    wire N__48675;
    wire N__48672;
    wire N__48669;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48653;
    wire N__48650;
    wire N__48649;
    wire N__48648;
    wire N__48645;
    wire N__48642;
    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48635;
    wire N__48632;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48622;
    wire N__48621;
    wire N__48620;
    wire N__48619;
    wire N__48618;
    wire N__48613;
    wire N__48610;
    wire N__48609;
    wire N__48608;
    wire N__48607;
    wire N__48606;
    wire N__48605;
    wire N__48604;
    wire N__48603;
    wire N__48602;
    wire N__48599;
    wire N__48596;
    wire N__48595;
    wire N__48592;
    wire N__48591;
    wire N__48586;
    wire N__48579;
    wire N__48574;
    wire N__48571;
    wire N__48570;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48558;
    wire N__48557;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48539;
    wire N__48532;
    wire N__48525;
    wire N__48524;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48510;
    wire N__48505;
    wire N__48502;
    wire N__48497;
    wire N__48492;
    wire N__48491;
    wire N__48490;
    wire N__48489;
    wire N__48488;
    wire N__48487;
    wire N__48484;
    wire N__48483;
    wire N__48482;
    wire N__48481;
    wire N__48480;
    wire N__48475;
    wire N__48470;
    wire N__48459;
    wire N__48454;
    wire N__48449;
    wire N__48446;
    wire N__48441;
    wire N__48438;
    wire N__48429;
    wire N__48424;
    wire N__48415;
    wire N__48412;
    wire N__48407;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48399;
    wire N__48390;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48378;
    wire N__48373;
    wire N__48372;
    wire N__48367;
    wire N__48362;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48321;
    wire N__48316;
    wire N__48311;
    wire N__48308;
    wire N__48303;
    wire N__48300;
    wire N__48295;
    wire N__48292;
    wire N__48287;
    wire N__48286;
    wire N__48283;
    wire N__48278;
    wire N__48273;
    wire N__48266;
    wire N__48259;
    wire N__48252;
    wire N__48249;
    wire N__48246;
    wire N__48243;
    wire N__48236;
    wire N__48233;
    wire N__48222;
    wire N__48221;
    wire N__48220;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48193;
    wire N__48190;
    wire N__48187;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48171;
    wire N__48170;
    wire N__48169;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48161;
    wire N__48158;
    wire N__48157;
    wire N__48154;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48139;
    wire N__48138;
    wire N__48135;
    wire N__48130;
    wire N__48127;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48084;
    wire N__48081;
    wire N__48080;
    wire N__48079;
    wire N__48078;
    wire N__48077;
    wire N__48076;
    wire N__48075;
    wire N__48072;
    wire N__48071;
    wire N__48070;
    wire N__48065;
    wire N__48062;
    wire N__48057;
    wire N__48054;
    wire N__48051;
    wire N__48046;
    wire N__48043;
    wire N__48036;
    wire N__48035;
    wire N__48034;
    wire N__48033;
    wire N__48032;
    wire N__48031;
    wire N__48030;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48018;
    wire N__48017;
    wire N__48012;
    wire N__48009;
    wire N__48004;
    wire N__47999;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47977;
    wire N__47972;
    wire N__47969;
    wire N__47966;
    wire N__47961;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47944;
    wire N__47941;
    wire N__47938;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47915;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47875;
    wire N__47872;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47859;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47842;
    wire N__47839;
    wire N__47834;
    wire N__47831;
    wire N__47826;
    wire N__47821;
    wire N__47814;
    wire N__47811;
    wire N__47810;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47754;
    wire N__47751;
    wire N__47746;
    wire N__47741;
    wire N__47736;
    wire N__47735;
    wire N__47734;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47723;
    wire N__47720;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47691;
    wire N__47690;
    wire N__47689;
    wire N__47688;
    wire N__47687;
    wire N__47686;
    wire N__47685;
    wire N__47682;
    wire N__47681;
    wire N__47680;
    wire N__47679;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47673;
    wire N__47672;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47655;
    wire N__47652;
    wire N__47647;
    wire N__47646;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47634;
    wire N__47633;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47611;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47603;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47578;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47554;
    wire N__47551;
    wire N__47550;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47519;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47495;
    wire N__47492;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47471;
    wire N__47466;
    wire N__47463;
    wire N__47458;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47407;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47395;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47381;
    wire N__47380;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47365;
    wire N__47362;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47332;
    wire N__47329;
    wire N__47324;
    wire N__47321;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47313;
    wire N__47308;
    wire N__47299;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47273;
    wire N__47264;
    wire N__47261;
    wire N__47260;
    wire N__47259;
    wire N__47258;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47249;
    wire N__47246;
    wire N__47243;
    wire N__47238;
    wire N__47237;
    wire N__47236;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47210;
    wire N__47205;
    wire N__47202;
    wire N__47197;
    wire N__47192;
    wire N__47183;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47167;
    wire N__47162;
    wire N__47145;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47130;
    wire N__47129;
    wire N__47128;
    wire N__47127;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47121;
    wire N__47120;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47116;
    wire N__47115;
    wire N__47112;
    wire N__47111;
    wire N__47108;
    wire N__47105;
    wire N__47102;
    wire N__47097;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47085;
    wire N__47082;
    wire N__47081;
    wire N__47080;
    wire N__47077;
    wire N__47074;
    wire N__47073;
    wire N__47072;
    wire N__47071;
    wire N__47070;
    wire N__47067;
    wire N__47066;
    wire N__47065;
    wire N__47064;
    wire N__47063;
    wire N__47060;
    wire N__47059;
    wire N__47058;
    wire N__47055;
    wire N__47050;
    wire N__47047;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47027;
    wire N__47024;
    wire N__47019;
    wire N__47016;
    wire N__47011;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46995;
    wire N__46990;
    wire N__46987;
    wire N__46978;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46968;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46945;
    wire N__46940;
    wire N__46933;
    wire N__46922;
    wire N__46919;
    wire N__46914;
    wire N__46899;
    wire N__46896;
    wire N__46891;
    wire N__46884;
    wire N__46879;
    wire N__46874;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46821;
    wire N__46818;
    wire N__46815;
    wire N__46814;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46792;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46778;
    wire N__46775;
    wire N__46772;
    wire N__46769;
    wire N__46762;
    wire N__46757;
    wire N__46752;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46738;
    wire N__46735;
    wire N__46730;
    wire N__46719;
    wire N__46716;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46708;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46682;
    wire N__46679;
    wire N__46676;
    wire N__46671;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46655;
    wire N__46654;
    wire N__46649;
    wire N__46646;
    wire N__46645;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46637;
    wire N__46634;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46615;
    wire N__46608;
    wire N__46605;
    wire N__46604;
    wire N__46599;
    wire N__46596;
    wire N__46595;
    wire N__46594;
    wire N__46591;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46575;
    wire N__46572;
    wire N__46563;
    wire N__46562;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46535;
    wire N__46534;
    wire N__46533;
    wire N__46530;
    wire N__46527;
    wire N__46524;
    wire N__46521;
    wire N__46520;
    wire N__46517;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46488;
    wire N__46487;
    wire N__46486;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46475;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46467;
    wire N__46464;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46429;
    wire N__46416;
    wire N__46415;
    wire N__46412;
    wire N__46411;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46401;
    wire N__46398;
    wire N__46397;
    wire N__46394;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46382;
    wire N__46379;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46356;
    wire N__46353;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46345;
    wire N__46342;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46320;
    wire N__46317;
    wire N__46308;
    wire N__46305;
    wire N__46304;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46287;
    wire N__46284;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46263;
    wire N__46262;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46235;
    wire N__46234;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46222;
    wire N__46219;
    wire N__46212;
    wire N__46211;
    wire N__46210;
    wire N__46207;
    wire N__46206;
    wire N__46205;
    wire N__46202;
    wire N__46201;
    wire N__46198;
    wire N__46197;
    wire N__46196;
    wire N__46195;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46188;
    wire N__46187;
    wire N__46186;
    wire N__46185;
    wire N__46184;
    wire N__46181;
    wire N__46170;
    wire N__46167;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46163;
    wire N__46162;
    wire N__46161;
    wire N__46160;
    wire N__46159;
    wire N__46158;
    wire N__46157;
    wire N__46152;
    wire N__46151;
    wire N__46150;
    wire N__46145;
    wire N__46140;
    wire N__46139;
    wire N__46136;
    wire N__46127;
    wire N__46124;
    wire N__46123;
    wire N__46122;
    wire N__46121;
    wire N__46120;
    wire N__46119;
    wire N__46118;
    wire N__46117;
    wire N__46116;
    wire N__46113;
    wire N__46106;
    wire N__46101;
    wire N__46096;
    wire N__46093;
    wire N__46092;
    wire N__46091;
    wire N__46090;
    wire N__46089;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46077;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46065;
    wire N__46064;
    wire N__46061;
    wire N__46056;
    wire N__46053;
    wire N__46046;
    wire N__46039;
    wire N__46034;
    wire N__46027;
    wire N__46018;
    wire N__46017;
    wire N__46014;
    wire N__46007;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45968;
    wire N__45963;
    wire N__45956;
    wire N__45953;
    wire N__45952;
    wire N__45949;
    wire N__45944;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45926;
    wire N__45921;
    wire N__45916;
    wire N__45913;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45889;
    wire N__45886;
    wire N__45881;
    wire N__45878;
    wire N__45861;
    wire N__45858;
    wire N__45857;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45819;
    wire N__45816;
    wire N__45815;
    wire N__45814;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45791;
    wire N__45790;
    wire N__45789;
    wire N__45786;
    wire N__45781;
    wire N__45778;
    wire N__45773;
    wire N__45770;
    wire N__45767;
    wire N__45766;
    wire N__45763;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45739;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45684;
    wire N__45683;
    wire N__45682;
    wire N__45679;
    wire N__45674;
    wire N__45669;
    wire N__45668;
    wire N__45667;
    wire N__45664;
    wire N__45659;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45651;
    wire N__45650;
    wire N__45647;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45627;
    wire N__45626;
    wire N__45625;
    wire N__45622;
    wire N__45621;
    wire N__45618;
    wire N__45615;
    wire N__45614;
    wire N__45613;
    wire N__45610;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45576;
    wire N__45575;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45507;
    wire N__45506;
    wire N__45503;
    wire N__45500;
    wire N__45497;
    wire N__45494;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45444;
    wire N__45439;
    wire N__45436;
    wire N__45435;
    wire N__45432;
    wire N__45427;
    wire N__45424;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45410;
    wire N__45407;
    wire N__45404;
    wire N__45403;
    wire N__45398;
    wire N__45395;
    wire N__45394;
    wire N__45391;
    wire N__45386;
    wire N__45381;
    wire N__45380;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45288;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45278;
    wire N__45275;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45249;
    wire N__45248;
    wire N__45245;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45234;
    wire N__45233;
    wire N__45230;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45214;
    wire N__45207;
    wire N__45206;
    wire N__45203;
    wire N__45202;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45185;
    wire N__45182;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45167;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45147;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45116;
    wire N__45115;
    wire N__45108;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45093;
    wire N__45092;
    wire N__45089;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45079;
    wire N__45078;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45065;
    wire N__45062;
    wire N__45055;
    wire N__45052;
    wire N__45045;
    wire N__45042;
    wire N__45041;
    wire N__45040;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45022;
    wire N__45015;
    wire N__45014;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45003;
    wire N__44998;
    wire N__44995;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44968;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44933;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44888;
    wire N__44885;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44866;
    wire N__44859;
    wire N__44858;
    wire N__44857;
    wire N__44854;
    wire N__44853;
    wire N__44852;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44810;
    wire N__44807;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44754;
    wire N__44753;
    wire N__44750;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44742;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44732;
    wire N__44727;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44696;
    wire N__44691;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44683;
    wire N__44678;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44668;
    wire N__44661;
    wire N__44660;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44649;
    wire N__44646;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44625;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44615;
    wire N__44614;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44594;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44582;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44439;
    wire N__44438;
    wire N__44437;
    wire N__44434;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44419;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44375;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44326;
    wire N__44325;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44310;
    wire N__44309;
    wire N__44304;
    wire N__44299;
    wire N__44296;
    wire N__44291;
    wire N__44286;
    wire N__44285;
    wire N__44284;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44268;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44244;
    wire N__44241;
    wire N__44232;
    wire N__44231;
    wire N__44230;
    wire N__44229;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44189;
    wire N__44186;
    wire N__44181;
    wire N__44172;
    wire N__44171;
    wire N__44168;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44150;
    wire N__44147;
    wire N__44144;
    wire N__44141;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44112;
    wire N__44103;
    wire N__44100;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44057;
    wire N__44054;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43979;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43959;
    wire N__43958;
    wire N__43955;
    wire N__43954;
    wire N__43951;
    wire N__43950;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43845;
    wire N__43842;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43797;
    wire N__43794;
    wire N__43789;
    wire N__43786;
    wire N__43781;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43760;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43734;
    wire N__43731;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43710;
    wire N__43709;
    wire N__43708;
    wire N__43703;
    wire N__43700;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43685;
    wire N__43680;
    wire N__43679;
    wire N__43676;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43662;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43656;
    wire N__43655;
    wire N__43650;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43614;
    wire N__43611;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43603;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43591;
    wire N__43584;
    wire N__43583;
    wire N__43580;
    wire N__43579;
    wire N__43576;
    wire N__43575;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43545;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43533;
    wire N__43530;
    wire N__43529;
    wire N__43528;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43479;
    wire N__43478;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43463;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43437;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43424;
    wire N__43423;
    wire N__43420;
    wire N__43419;
    wire N__43418;
    wire N__43417;
    wire N__43414;
    wire N__43413;
    wire N__43412;
    wire N__43411;
    wire N__43410;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43395;
    wire N__43394;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43383;
    wire N__43382;
    wire N__43377;
    wire N__43376;
    wire N__43373;
    wire N__43372;
    wire N__43369;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43347;
    wire N__43346;
    wire N__43343;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43320;
    wire N__43319;
    wire N__43318;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43308;
    wire N__43301;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43282;
    wire N__43279;
    wire N__43274;
    wire N__43271;
    wire N__43270;
    wire N__43269;
    wire N__43266;
    wire N__43265;
    wire N__43264;
    wire N__43261;
    wire N__43260;
    wire N__43259;
    wire N__43254;
    wire N__43249;
    wire N__43244;
    wire N__43239;
    wire N__43230;
    wire N__43227;
    wire N__43222;
    wire N__43217;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43152;
    wire N__43149;
    wire N__43148;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43052;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42977;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42957;
    wire N__42952;
    wire N__42949;
    wire N__42942;
    wire N__42941;
    wire N__42938;
    wire N__42937;
    wire N__42934;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42906;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42873;
    wire N__42872;
    wire N__42871;
    wire N__42870;
    wire N__42869;
    wire N__42868;
    wire N__42867;
    wire N__42866;
    wire N__42865;
    wire N__42864;
    wire N__42863;
    wire N__42862;
    wire N__42861;
    wire N__42860;
    wire N__42859;
    wire N__42858;
    wire N__42857;
    wire N__42852;
    wire N__42843;
    wire N__42836;
    wire N__42831;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42823;
    wire N__42822;
    wire N__42821;
    wire N__42820;
    wire N__42819;
    wire N__42818;
    wire N__42817;
    wire N__42816;
    wire N__42815;
    wire N__42814;
    wire N__42813;
    wire N__42812;
    wire N__42811;
    wire N__42810;
    wire N__42809;
    wire N__42808;
    wire N__42805;
    wire N__42804;
    wire N__42803;
    wire N__42802;
    wire N__42801;
    wire N__42800;
    wire N__42799;
    wire N__42798;
    wire N__42797;
    wire N__42792;
    wire N__42789;
    wire N__42782;
    wire N__42781;
    wire N__42780;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42758;
    wire N__42749;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42718;
    wire N__42713;
    wire N__42712;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42694;
    wire N__42691;
    wire N__42686;
    wire N__42683;
    wire N__42670;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42636;
    wire N__42627;
    wire N__42622;
    wire N__42619;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42601;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42525;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42513;
    wire N__42512;
    wire N__42509;
    wire N__42506;
    wire N__42503;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42493;
    wire N__42490;
    wire N__42489;
    wire N__42486;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42469;
    wire N__42466;
    wire N__42461;
    wire N__42456;
    wire N__42453;
    wire N__42448;
    wire N__42443;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42276;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42266;
    wire N__42265;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42241;
    wire N__42234;
    wire N__42231;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42223;
    wire N__42220;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42208;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42173;
    wire N__42170;
    wire N__42167;
    wire N__42166;
    wire N__42165;
    wire N__42160;
    wire N__42155;
    wire N__42150;
    wire N__42149;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42092;
    wire N__42091;
    wire N__42088;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42054;
    wire N__42053;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42043;
    wire N__42040;
    wire N__42039;
    wire N__42036;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41954;
    wire N__41951;
    wire N__41950;
    wire N__41947;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41883;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41868;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41860;
    wire N__41859;
    wire N__41854;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41836;
    wire N__41833;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41816;
    wire N__41815;
    wire N__41812;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41782;
    wire N__41779;
    wire N__41774;
    wire N__41771;
    wire N__41766;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41760;
    wire N__41755;
    wire N__41752;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41731;
    wire N__41724;
    wire N__41723;
    wire N__41722;
    wire N__41719;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41704;
    wire N__41703;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41686;
    wire N__41679;
    wire N__41678;
    wire N__41675;
    wire N__41674;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41632;
    wire N__41625;
    wire N__41624;
    wire N__41621;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41593;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41564;
    wire N__41561;
    wire N__41556;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41530;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41479;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41454;
    wire N__41453;
    wire N__41452;
    wire N__41451;
    wire N__41448;
    wire N__41447;
    wire N__41446;
    wire N__41443;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41415;
    wire N__41414;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41406;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41383;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41366;
    wire N__41365;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41324;
    wire N__41323;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41301;
    wire N__41298;
    wire N__41289;
    wire N__41288;
    wire N__41285;
    wire N__41284;
    wire N__41281;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41263;
    wire N__41262;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41229;
    wire N__41228;
    wire N__41227;
    wire N__41224;
    wire N__41219;
    wire N__41218;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41200;
    wire N__41197;
    wire N__41190;
    wire N__41189;
    wire N__41186;
    wire N__41185;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41154;
    wire N__41151;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41090;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41082;
    wire N__41079;
    wire N__41078;
    wire N__41077;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41059;
    wire N__41056;
    wire N__41051;
    wire N__41044;
    wire N__41037;
    wire N__41036;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41004;
    wire N__41001;
    wire N__40992;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40950;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40942;
    wire N__40941;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40929;
    wire N__40928;
    wire N__40925;
    wire N__40918;
    wire N__40915;
    wire N__40910;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40892;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40877;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40845;
    wire N__40844;
    wire N__40841;
    wire N__40840;
    wire N__40839;
    wire N__40836;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40787;
    wire N__40786;
    wire N__40783;
    wire N__40778;
    wire N__40777;
    wire N__40776;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40761;
    wire N__40752;
    wire N__40751;
    wire N__40750;
    wire N__40747;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40689;
    wire N__40688;
    wire N__40685;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40657;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40589;
    wire N__40588;
    wire N__40587;
    wire N__40582;
    wire N__40577;
    wire N__40576;
    wire N__40571;
    wire N__40568;
    wire N__40565;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40550;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40536;
    wire N__40535;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40516;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40468;
    wire N__40463;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40437;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40407;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40389;
    wire N__40386;
    wire N__40381;
    wire N__40378;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40323;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40311;
    wire N__40310;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40286;
    wire N__40281;
    wire N__40278;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40245;
    wire N__40244;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40226;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40194;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40148;
    wire N__40147;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40131;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40101;
    wire N__40098;
    wire N__40097;
    wire N__40096;
    wire N__40093;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40051;
    wire N__40044;
    wire N__40041;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39986;
    wire N__39985;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39973;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39942;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39931;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39919;
    wire N__39916;
    wire N__39909;
    wire N__39908;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39837;
    wire N__39836;
    wire N__39835;
    wire N__39834;
    wire N__39831;
    wire N__39826;
    wire N__39823;
    wire N__39822;
    wire N__39821;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39792;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39774;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39756;
    wire N__39755;
    wire N__39752;
    wire N__39751;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39743;
    wire N__39742;
    wire N__39741;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39705;
    wire N__39704;
    wire N__39701;
    wire N__39700;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39669;
    wire N__39666;
    wire N__39661;
    wire N__39654;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39636;
    wire N__39633;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39625;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39576;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39558;
    wire N__39555;
    wire N__39554;
    wire N__39553;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39539;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39525;
    wire N__39520;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39503;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39492;
    wire N__39489;
    wire N__39484;
    wire N__39481;
    wire N__39478;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39460;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39424;
    wire N__39419;
    wire N__39416;
    wire N__39415;
    wire N__39412;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39394;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39343;
    wire N__39342;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39326;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39306;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39291;
    wire N__39288;
    wire N__39287;
    wire N__39284;
    wire N__39283;
    wire N__39282;
    wire N__39279;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39265;
    wire N__39262;
    wire N__39257;
    wire N__39252;
    wire N__39249;
    wire N__39244;
    wire N__39237;
    wire N__39234;
    wire N__39233;
    wire N__39232;
    wire N__39231;
    wire N__39230;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39208;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39148;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39136;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39111;
    wire N__39108;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39090;
    wire N__39087;
    wire N__39086;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39071;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39056;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38985;
    wire N__38982;
    wire N__38981;
    wire N__38980;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38940;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38910;
    wire N__38907;
    wire N__38906;
    wire N__38905;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38880;
    wire N__38877;
    wire N__38872;
    wire N__38865;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38850;
    wire N__38847;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38839;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38790;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38720;
    wire N__38719;
    wire N__38716;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38702;
    wire N__38699;
    wire N__38694;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38673;
    wire N__38664;
    wire N__38661;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38650;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38612;
    wire N__38609;
    wire N__38604;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38549;
    wire N__38546;
    wire N__38543;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38519;
    wire N__38508;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38463;
    wire N__38460;
    wire N__38459;
    wire N__38454;
    wire N__38451;
    wire N__38450;
    wire N__38449;
    wire N__38446;
    wire N__38445;
    wire N__38442;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38392;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38381;
    wire N__38378;
    wire N__38375;
    wire N__38370;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38340;
    wire N__38337;
    wire N__38336;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38321;
    wire N__38320;
    wire N__38317;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38289;
    wire N__38280;
    wire N__38277;
    wire N__38276;
    wire N__38275;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38228;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38190;
    wire N__38187;
    wire N__38186;
    wire N__38183;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38133;
    wire N__38130;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38112;
    wire N__38109;
    wire N__38108;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38091;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38083;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38065;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37859;
    wire N__37858;
    wire N__37855;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37843;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37831;
    wire N__37828;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37771;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37743;
    wire N__37742;
    wire N__37741;
    wire N__37740;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37710;
    wire N__37707;
    wire N__37702;
    wire N__37699;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37679;
    wire N__37676;
    wire N__37675;
    wire N__37672;
    wire N__37671;
    wire N__37668;
    wire N__37663;
    wire N__37660;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37626;
    wire N__37623;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37545;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37537;
    wire N__37536;
    wire N__37535;
    wire N__37534;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37469;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37443;
    wire N__37442;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37434;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37419;
    wire N__37412;
    wire N__37407;
    wire N__37404;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37390;
    wire N__37389;
    wire N__37388;
    wire N__37383;
    wire N__37378;
    wire N__37375;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37336;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37284;
    wire N__37283;
    wire N__37282;
    wire N__37279;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37261;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37235;
    wire N__37232;
    wire N__37221;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37213;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37193;
    wire N__37188;
    wire N__37187;
    wire N__37184;
    wire N__37183;
    wire N__37180;
    wire N__37179;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37140;
    wire N__37139;
    wire N__37138;
    wire N__37135;
    wire N__37130;
    wire N__37129;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37101;
    wire N__37098;
    wire N__37097;
    wire N__37094;
    wire N__37093;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37071;
    wire N__37070;
    wire N__37067;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37052;
    wire N__37047;
    wire N__37044;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37036;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36993;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36972;
    wire N__36969;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36938;
    wire N__36937;
    wire N__36934;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36912;
    wire N__36909;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36854;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36831;
    wire N__36830;
    wire N__36829;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36794;
    wire N__36791;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36754;
    wire N__36747;
    wire N__36746;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36735;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36717;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36709;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36689;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36646;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36630;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36624;
    wire N__36623;
    wire N__36620;
    wire N__36615;
    wire N__36610;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36540;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36525;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36428;
    wire N__36427;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36407;
    wire N__36402;
    wire N__36399;
    wire N__36398;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36315;
    wire N__36314;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36228;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36220;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36185;
    wire N__36184;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36153;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36138;
    wire N__36135;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36071;
    wire N__36070;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36019;
    wire N__36012;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35988;
    wire N__35985;
    wire N__35984;
    wire N__35981;
    wire N__35980;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35968;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35900;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35894;
    wire N__35889;
    wire N__35884;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35854;
    wire N__35853;
    wire N__35852;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35830;
    wire N__35823;
    wire N__35822;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35810;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35665;
    wire N__35664;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35656;
    wire N__35649;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35639;
    wire N__35638;
    wire N__35633;
    wire N__35630;
    wire N__35625;
    wire N__35620;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35603;
    wire N__35600;
    wire N__35593;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35577;
    wire N__35576;
    wire N__35575;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35547;
    wire N__35546;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35516;
    wire N__35513;
    wire N__35512;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35486;
    wire N__35477;
    wire N__35472;
    wire N__35471;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35463;
    wire N__35462;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35441;
    wire N__35438;
    wire N__35433;
    wire N__35430;
    wire N__35423;
    wire N__35420;
    wire N__35415;
    wire N__35412;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35364;
    wire N__35359;
    wire N__35352;
    wire N__35351;
    wire N__35348;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35337;
    wire N__35334;
    wire N__35329;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35304;
    wire N__35301;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35249;
    wire N__35248;
    wire N__35247;
    wire N__35246;
    wire N__35245;
    wire N__35240;
    wire N__35237;
    wire N__35236;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35213;
    wire N__35208;
    wire N__35203;
    wire N__35196;
    wire N__35195;
    wire N__35194;
    wire N__35193;
    wire N__35192;
    wire N__35191;
    wire N__35190;
    wire N__35187;
    wire N__35180;
    wire N__35177;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35157;
    wire N__35154;
    wire N__35145;
    wire N__35144;
    wire N__35141;
    wire N__35134;
    wire N__35127;
    wire N__35120;
    wire N__35117;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35081;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35073;
    wire N__35072;
    wire N__35071;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35055;
    wire N__35050;
    wire N__35049;
    wire N__35046;
    wire N__35041;
    wire N__35038;
    wire N__35033;
    wire N__35030;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34913;
    wire N__34912;
    wire N__34911;
    wire N__34910;
    wire N__34905;
    wire N__34900;
    wire N__34897;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34877;
    wire N__34876;
    wire N__34873;
    wire N__34872;
    wire N__34871;
    wire N__34870;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34862;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34856;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34844;
    wire N__34839;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34784;
    wire N__34775;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34763;
    wire N__34760;
    wire N__34753;
    wire N__34746;
    wire N__34743;
    wire N__34728;
    wire N__34725;
    wire N__34724;
    wire N__34723;
    wire N__34720;
    wire N__34715;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34691;
    wire N__34688;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34674;
    wire N__34669;
    wire N__34666;
    wire N__34661;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34646;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34613;
    wire N__34608;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34569;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34525;
    wire N__34520;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34499;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34405;
    wire N__34400;
    wire N__34395;
    wire N__34394;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34343;
    wire N__34342;
    wire N__34341;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34333;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34273;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34247;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34230;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34213;
    wire N__34212;
    wire N__34211;
    wire N__34210;
    wire N__34209;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34186;
    wire N__34185;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34179;
    wire N__34172;
    wire N__34165;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34143;
    wire N__34132;
    wire N__34129;
    wire N__34128;
    wire N__34127;
    wire N__34126;
    wire N__34123;
    wire N__34118;
    wire N__34113;
    wire N__34106;
    wire N__34101;
    wire N__34098;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34080;
    wire N__34073;
    wire N__34050;
    wire N__34049;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34013;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33938;
    wire N__33937;
    wire N__33936;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33918;
    wire N__33915;
    wire N__33914;
    wire N__33911;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33895;
    wire N__33892;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33882;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33866;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33854;
    wire N__33853;
    wire N__33852;
    wire N__33851;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33835;
    wire N__33834;
    wire N__33831;
    wire N__33826;
    wire N__33823;
    wire N__33818;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33795;
    wire N__33794;
    wire N__33791;
    wire N__33790;
    wire N__33789;
    wire N__33788;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33772;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33752;
    wire N__33749;
    wire N__33748;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33707;
    wire N__33706;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33668;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33645;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33618;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33603;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33573;
    wire N__33570;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33558;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33543;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33497;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33471;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33450;
    wire N__33447;
    wire N__33446;
    wire N__33445;
    wire N__33442;
    wire N__33437;
    wire N__33432;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33383;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33345;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33333;
    wire N__33332;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33324;
    wire N__33321;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33284;
    wire N__33283;
    wire N__33282;
    wire N__33281;
    wire N__33278;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33264;
    wire N__33263;
    wire N__33260;
    wire N__33259;
    wire N__33256;
    wire N__33255;
    wire N__33250;
    wire N__33241;
    wire N__33238;
    wire N__33237;
    wire N__33230;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33180;
    wire N__33179;
    wire N__33178;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33170;
    wire N__33169;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33146;
    wire N__33143;
    wire N__33142;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33113;
    wire N__33108;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33090;
    wire N__33089;
    wire N__33088;
    wire N__33087;
    wire N__33084;
    wire N__33083;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33062;
    wire N__33061;
    wire N__33060;
    wire N__33059;
    wire N__33058;
    wire N__33057;
    wire N__33052;
    wire N__33041;
    wire N__33038;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32934;
    wire N__32933;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32907;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32901;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32877;
    wire N__32874;
    wire N__32867;
    wire N__32862;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32839;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32682;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32618;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32585;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32542;
    wire N__32535;
    wire N__32532;
    wire N__32531;
    wire N__32530;
    wire N__32529;
    wire N__32526;
    wire N__32525;
    wire N__32524;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32493;
    wire N__32490;
    wire N__32485;
    wire N__32484;
    wire N__32481;
    wire N__32474;
    wire N__32469;
    wire N__32466;
    wire N__32457;
    wire N__32454;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32439;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32424;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32357;
    wire N__32354;
    wire N__32353;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32294;
    wire N__32293;
    wire N__32288;
    wire N__32285;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32258;
    wire N__32257;
    wire N__32256;
    wire N__32253;
    wire N__32246;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32165;
    wire N__32164;
    wire N__32161;
    wire N__32156;
    wire N__32153;
    wire N__32148;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32132;
    wire N__32131;
    wire N__32130;
    wire N__32129;
    wire N__32126;
    wire N__32121;
    wire N__32120;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32076;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32064;
    wire N__32061;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32046;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32020;
    wire N__32019;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32003;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31938;
    wire N__31935;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31856;
    wire N__31855;
    wire N__31854;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31809;
    wire N__31806;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31784;
    wire N__31781;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31599;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31587;
    wire N__31586;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31487;
    wire N__31486;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31474;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31460;
    wire N__31459;
    wire N__31456;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31441;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31398;
    wire N__31397;
    wire N__31396;
    wire N__31395;
    wire N__31392;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31380;
    wire N__31379;
    wire N__31374;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31350;
    wire N__31349;
    wire N__31348;
    wire N__31347;
    wire N__31346;
    wire N__31345;
    wire N__31344;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31327;
    wire N__31326;
    wire N__31325;
    wire N__31322;
    wire N__31315;
    wire N__31308;
    wire N__31305;
    wire N__31296;
    wire N__31295;
    wire N__31294;
    wire N__31293;
    wire N__31292;
    wire N__31291;
    wire N__31290;
    wire N__31289;
    wire N__31286;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31261;
    wire N__31258;
    wire N__31253;
    wire N__31252;
    wire N__31247;
    wire N__31242;
    wire N__31239;
    wire N__31232;
    wire N__31229;
    wire N__31218;
    wire N__31217;
    wire N__31216;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31208;
    wire N__31207;
    wire N__31202;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31170;
    wire N__31169;
    wire N__31168;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31154;
    wire N__31153;
    wire N__31152;
    wire N__31151;
    wire N__31150;
    wire N__31149;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31137;
    wire N__31134;
    wire N__31129;
    wire N__31126;
    wire N__31121;
    wire N__31110;
    wire N__31109;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31035;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31020;
    wire N__31017;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31005;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30982;
    wire N__30979;
    wire N__30968;
    wire N__30961;
    wire N__30954;
    wire N__30953;
    wire N__30952;
    wire N__30951;
    wire N__30950;
    wire N__30949;
    wire N__30948;
    wire N__30943;
    wire N__30932;
    wire N__30927;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30876;
    wire N__30875;
    wire N__30870;
    wire N__30867;
    wire N__30866;
    wire N__30863;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30834;
    wire N__30831;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30774;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30744;
    wire N__30739;
    wire N__30726;
    wire N__30725;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30643;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30600;
    wire N__30599;
    wire N__30592;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30555;
    wire N__30554;
    wire N__30553;
    wire N__30552;
    wire N__30551;
    wire N__30548;
    wire N__30547;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30520;
    wire N__30519;
    wire N__30518;
    wire N__30517;
    wire N__30512;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30492;
    wire N__30489;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30449;
    wire N__30444;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30435;
    wire N__30434;
    wire N__30431;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30417;
    wire N__30416;
    wire N__30407;
    wire N__30404;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30372;
    wire N__30369;
    wire N__30368;
    wire N__30367;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30356;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30344;
    wire N__30341;
    wire N__30340;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30317;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30213;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30162;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30150;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30114;
    wire N__30113;
    wire N__30112;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30108;
    wire N__30105;
    wire N__30100;
    wire N__30097;
    wire N__30090;
    wire N__30083;
    wire N__30072;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30068;
    wire N__30067;
    wire N__30066;
    wire N__30061;
    wire N__30058;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30046;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30036;
    wire N__30035;
    wire N__30034;
    wire N__30031;
    wire N__30026;
    wire N__30023;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30011;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__29997;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29979;
    wire N__29974;
    wire N__29967;
    wire N__29962;
    wire N__29957;
    wire N__29950;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29927;
    wire N__29926;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29918;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29850;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29828;
    wire N__29825;
    wire N__29818;
    wire N__29815;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29664;
    wire N__29661;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29646;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29631;
    wire N__29628;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29616;
    wire N__29613;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29601;
    wire N__29598;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29586;
    wire N__29583;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29558;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29546;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29483;
    wire N__29480;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29450;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29354;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29257;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29186;
    wire N__29181;
    wire N__29178;
    wire N__29177;
    wire N__29174;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29159;
    wire N__29154;
    wire N__29151;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29138;
    wire N__29135;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29022;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28988;
    wire N__28987;
    wire N__28986;
    wire N__28985;
    wire N__28984;
    wire N__28983;
    wire N__28982;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28961;
    wire N__28958;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28938;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28925;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28905;
    wire N__28900;
    wire N__28893;
    wire N__28892;
    wire N__28887;
    wire N__28884;
    wire N__28883;
    wire N__28882;
    wire N__28879;
    wire N__28874;
    wire N__28869;
    wire N__28868;
    wire N__28863;
    wire N__28862;
    wire N__28861;
    wire N__28860;
    wire N__28859;
    wire N__28858;
    wire N__28855;
    wire N__28850;
    wire N__28843;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28805;
    wire N__28804;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28793;
    wire N__28792;
    wire N__28791;
    wire N__28788;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28767;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28698;
    wire N__28697;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28659;
    wire N__28656;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28646;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28479;
    wire N__28476;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28464;
    wire N__28461;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28421;
    wire N__28418;
    wire N__28417;
    wire N__28414;
    wire N__28409;
    wire N__28404;
    wire N__28401;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28389;
    wire N__28386;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28371;
    wire N__28368;
    wire N__28367;
    wire N__28366;
    wire N__28363;
    wire N__28358;
    wire N__28353;
    wire N__28350;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28338;
    wire N__28335;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28323;
    wire N__28320;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28253;
    wire N__28252;
    wire N__28251;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28224;
    wire N__28223;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28200;
    wire N__28199;
    wire N__28198;
    wire N__28197;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28154;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28139;
    wire N__28138;
    wire N__28137;
    wire N__28136;
    wire N__28135;
    wire N__28132;
    wire N__28127;
    wire N__28124;
    wire N__28123;
    wire N__28120;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28106;
    wire N__28103;
    wire N__28102;
    wire N__28095;
    wire N__28090;
    wire N__28087;
    wire N__28086;
    wire N__28083;
    wire N__28082;
    wire N__28077;
    wire N__28070;
    wire N__28063;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28042;
    wire N__28037;
    wire N__28034;
    wire N__28023;
    wire N__28022;
    wire N__28021;
    wire N__28020;
    wire N__28015;
    wire N__28012;
    wire N__28011;
    wire N__28010;
    wire N__28007;
    wire N__28006;
    wire N__28005;
    wire N__28000;
    wire N__27999;
    wire N__27994;
    wire N__27993;
    wire N__27990;
    wire N__27985;
    wire N__27982;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27948;
    wire N__27947;
    wire N__27946;
    wire N__27945;
    wire N__27944;
    wire N__27943;
    wire N__27942;
    wire N__27941;
    wire N__27940;
    wire N__27939;
    wire N__27938;
    wire N__27935;
    wire N__27930;
    wire N__27927;
    wire N__27926;
    wire N__27921;
    wire N__27920;
    wire N__27911;
    wire N__27908;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27866;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27846;
    wire N__27845;
    wire N__27842;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27823;
    wire N__27810;
    wire N__27809;
    wire N__27808;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27797;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27763;
    wire N__27758;
    wire N__27753;
    wire N__27752;
    wire N__27749;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27729;
    wire N__27728;
    wire N__27727;
    wire N__27722;
    wire N__27719;
    wire N__27714;
    wire N__27713;
    wire N__27712;
    wire N__27711;
    wire N__27704;
    wire N__27701;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27689;
    wire N__27688;
    wire N__27685;
    wire N__27680;
    wire N__27675;
    wire N__27674;
    wire N__27673;
    wire N__27670;
    wire N__27665;
    wire N__27660;
    wire N__27659;
    wire N__27658;
    wire N__27655;
    wire N__27650;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27623;
    wire N__27622;
    wire N__27621;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27604;
    wire N__27599;
    wire N__27596;
    wire N__27591;
    wire N__27588;
    wire N__27587;
    wire N__27586;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27561;
    wire N__27556;
    wire N__27549;
    wire N__27548;
    wire N__27547;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27474;
    wire N__27469;
    wire N__27456;
    wire N__27455;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27436;
    wire N__27435;
    wire N__27434;
    wire N__27431;
    wire N__27430;
    wire N__27429;
    wire N__27428;
    wire N__27423;
    wire N__27416;
    wire N__27411;
    wire N__27410;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27372;
    wire N__27371;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27297;
    wire N__27294;
    wire N__27293;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27258;
    wire N__27255;
    wire N__27254;
    wire N__27253;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27241;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27218;
    wire N__27217;
    wire N__27216;
    wire N__27213;
    wire N__27212;
    wire N__27211;
    wire N__27206;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27156;
    wire N__27155;
    wire N__27152;
    wire N__27151;
    wire N__27150;
    wire N__27145;
    wire N__27140;
    wire N__27135;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27121;
    wire N__27116;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27080;
    wire N__27075;
    wire N__27066;
    wire N__27063;
    wire N__27062;
    wire N__27061;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27039;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27031;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27016;
    wire N__27009;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__27001;
    wire N__27000;
    wire N__26997;
    wire N__26992;
    wire N__26989;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26967;
    wire N__26964;
    wire N__26959;
    wire N__26958;
    wire N__26957;
    wire N__26956;
    wire N__26955;
    wire N__26954;
    wire N__26951;
    wire N__26946;
    wire N__26943;
    wire N__26938;
    wire N__26933;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26903;
    wire N__26902;
    wire N__26901;
    wire N__26896;
    wire N__26891;
    wire N__26886;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26871;
    wire N__26870;
    wire N__26867;
    wire N__26866;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26837;
    wire N__26834;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26807;
    wire N__26804;
    wire N__26803;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26783;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26705;
    wire N__26704;
    wire N__26703;
    wire N__26700;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26684;
    wire N__26681;
    wire N__26676;
    wire N__26673;
    wire N__26664;
    wire N__26661;
    wire N__26660;
    wire N__26659;
    wire N__26656;
    wire N__26651;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26633;
    wire N__26630;
    wire N__26629;
    wire N__26628;
    wire N__26625;
    wire N__26624;
    wire N__26621;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26585;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26571;
    wire N__26568;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26550;
    wire N__26549;
    wire N__26546;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26529;
    wire N__26528;
    wire N__26527;
    wire N__26524;
    wire N__26523;
    wire N__26520;
    wire N__26515;
    wire N__26512;
    wire N__26505;
    wire N__26502;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26496;
    wire N__26495;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26475;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26460;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26439;
    wire N__26436;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26424;
    wire N__26423;
    wire N__26422;
    wire N__26421;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26403;
    wire N__26394;
    wire N__26393;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26378;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26343;
    wire N__26340;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26307;
    wire N__26304;
    wire N__26303;
    wire N__26302;
    wire N__26299;
    wire N__26298;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26226;
    wire N__26223;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26175;
    wire N__26174;
    wire N__26171;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26142;
    wire N__26141;
    wire N__26136;
    wire N__26133;
    wire N__26132;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26112;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26097;
    wire N__26094;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26067;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26052;
    wire N__26043;
    wire N__26042;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26025;
    wire N__26022;
    wire N__26013;
    wire N__26012;
    wire N__26009;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__26003;
    wire N__26002;
    wire N__25999;
    wire N__25998;
    wire N__25995;
    wire N__25994;
    wire N__25991;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25966;
    wire N__25953;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25937;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25917;
    wire N__25914;
    wire N__25913;
    wire N__25910;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25902;
    wire N__25901;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25883;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25865;
    wire N__25864;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25841;
    wire N__25830;
    wire N__25827;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25785;
    wire N__25784;
    wire N__25783;
    wire N__25782;
    wire N__25781;
    wire N__25780;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25729;
    wire N__25716;
    wire N__25715;
    wire N__25714;
    wire N__25713;
    wire N__25712;
    wire N__25711;
    wire N__25710;
    wire N__25707;
    wire N__25706;
    wire N__25705;
    wire N__25704;
    wire N__25703;
    wire N__25702;
    wire N__25701;
    wire N__25700;
    wire N__25689;
    wire N__25686;
    wire N__25679;
    wire N__25678;
    wire N__25677;
    wire N__25674;
    wire N__25673;
    wire N__25672;
    wire N__25671;
    wire N__25670;
    wire N__25663;
    wire N__25660;
    wire N__25659;
    wire N__25652;
    wire N__25649;
    wire N__25648;
    wire N__25647;
    wire N__25642;
    wire N__25635;
    wire N__25632;
    wire N__25627;
    wire N__25626;
    wire N__25623;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25607;
    wire N__25602;
    wire N__25599;
    wire N__25598;
    wire N__25597;
    wire N__25596;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25571;
    wire N__25568;
    wire N__25557;
    wire N__25556;
    wire N__25555;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25544;
    wire N__25543;
    wire N__25540;
    wire N__25533;
    wire N__25528;
    wire N__25523;
    wire N__25516;
    wire N__25507;
    wire N__25494;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25476;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25443;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25416;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25335;
    wire N__25332;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25288;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25207;
    wire N__25200;
    wire N__25199;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25185;
    wire N__25184;
    wire N__25183;
    wire N__25182;
    wire N__25179;
    wire N__25172;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25124;
    wire N__25123;
    wire N__25116;
    wire N__25115;
    wire N__25114;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25095;
    wire N__25086;
    wire N__25081;
    wire N__25074;
    wire N__25073;
    wire N__25070;
    wire N__25069;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25057;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25053;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25033;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24977;
    wire N__24974;
    wire N__24969;
    wire N__24966;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24956;
    wire N__24953;
    wire N__24948;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24938;
    wire N__24935;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24824;
    wire N__24823;
    wire N__24818;
    wire N__24815;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24700;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24673;
    wire N__24670;
    wire N__24665;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24644;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24633;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24626;
    wire N__24625;
    wire N__24624;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24617;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24586;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24569;
    wire N__24568;
    wire N__24567;
    wire N__24566;
    wire N__24565;
    wire N__24562;
    wire N__24549;
    wire N__24546;
    wire N__24537;
    wire N__24534;
    wire N__24533;
    wire N__24530;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24503;
    wire N__24502;
    wire N__24501;
    wire N__24500;
    wire N__24499;
    wire N__24498;
    wire N__24495;
    wire N__24490;
    wire N__24485;
    wire N__24482;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24448;
    wire N__24447;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24428;
    wire N__24425;
    wire N__24418;
    wire N__24415;
    wire N__24410;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24379;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24215;
    wire N__24214;
    wire N__24213;
    wire N__24208;
    wire N__24203;
    wire N__24198;
    wire N__24197;
    wire N__24196;
    wire N__24195;
    wire N__24192;
    wire N__24185;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24166;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24101;
    wire N__24098;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24081;
    wire N__24080;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23998;
    wire N__23995;
    wire N__23990;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23956;
    wire N__23949;
    wire N__23948;
    wire N__23943;
    wire N__23940;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23932;
    wire N__23927;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23915;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23911;
    wire N__23910;
    wire N__23909;
    wire N__23908;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23901;
    wire N__23898;
    wire N__23897;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23881;
    wire N__23878;
    wire N__23877;
    wire N__23876;
    wire N__23875;
    wire N__23872;
    wire N__23871;
    wire N__23868;
    wire N__23867;
    wire N__23864;
    wire N__23863;
    wire N__23860;
    wire N__23859;
    wire N__23858;
    wire N__23857;
    wire N__23856;
    wire N__23855;
    wire N__23854;
    wire N__23853;
    wire N__23846;
    wire N__23835;
    wire N__23824;
    wire N__23817;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23767;
    wire N__23764;
    wire N__23753;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23729;
    wire N__23718;
    wire N__23715;
    wire N__23714;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23694;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23636;
    wire N__23635;
    wire N__23634;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23626;
    wire N__23625;
    wire N__23622;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23587;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23575;
    wire N__23570;
    wire N__23567;
    wire N__23556;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23538;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23523;
    wire N__23520;
    wire N__23519;
    wire N__23516;
    wire N__23515;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23503;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23466;
    wire N__23463;
    wire N__23462;
    wire N__23461;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23446;
    wire N__23445;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23404;
    wire N__23403;
    wire N__23402;
    wire N__23401;
    wire N__23398;
    wire N__23393;
    wire N__23388;
    wire N__23381;
    wire N__23378;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23361;
    wire N__23360;
    wire N__23357;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23295;
    wire N__23294;
    wire N__23291;
    wire N__23290;
    wire N__23285;
    wire N__23282;
    wire N__23277;
    wire N__23274;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23251;
    wire N__23240;
    wire N__23231;
    wire N__23226;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23210;
    wire N__23207;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23180;
    wire N__23179;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23158;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23146;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23132;
    wire N__23131;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23109;
    wire N__23108;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23084;
    wire N__23083;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23040;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23013;
    wire N__23012;
    wire N__23011;
    wire N__23010;
    wire N__23007;
    wire N__23002;
    wire N__22999;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22985;
    wire N__22982;
    wire N__22981;
    wire N__22978;
    wire N__22977;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22965;
    wire N__22962;
    wire N__22953;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22931;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22854;
    wire N__22851;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22836;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22747;
    wire N__22742;
    wire N__22739;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22631;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22619;
    wire N__22618;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22568;
    wire N__22567;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22556;
    wire N__22547;
    wire N__22544;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22505;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22500;
    wire N__22499;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22495;
    wire N__22494;
    wire N__22493;
    wire N__22488;
    wire N__22481;
    wire N__22472;
    wire N__22463;
    wire N__22460;
    wire N__22453;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22384;
    wire N__22383;
    wire N__22378;
    wire N__22373;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22336;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22313;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22253;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22204;
    wire N__22201;
    wire N__22196;
    wire N__22193;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22158;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22045;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22026;
    wire N__22023;
    wire N__22018;
    wire N__22015;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21958;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21916;
    wire N__21915;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21904;
    wire N__21903;
    wire N__21902;
    wire N__21899;
    wire N__21898;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21883;
    wire N__21882;
    wire N__21881;
    wire N__21876;
    wire N__21871;
    wire N__21870;
    wire N__21863;
    wire N__21860;
    wire N__21847;
    wire N__21834;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21814;
    wire N__21813;
    wire N__21812;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21802;
    wire N__21797;
    wire N__21794;
    wire N__21789;
    wire N__21788;
    wire N__21781;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21763;
    wire N__21760;
    wire N__21747;
    wire N__21746;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21730;
    wire N__21725;
    wire N__21720;
    wire N__21717;
    wire N__21716;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21701;
    wire N__21700;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21679;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21669;
    wire N__21666;
    wire N__21665;
    wire N__21664;
    wire N__21663;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21647;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21623;
    wire N__21620;
    wire N__21611;
    wire N__21598;
    wire N__21595;
    wire N__21582;
    wire N__21579;
    wire N__21572;
    wire N__21567;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21535;
    wire N__21532;
    wire N__21531;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21512;
    wire N__21511;
    wire N__21510;
    wire N__21509;
    wire N__21508;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21486;
    wire N__21473;
    wire N__21460;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21452;
    wire N__21451;
    wire N__21450;
    wire N__21449;
    wire N__21448;
    wire N__21439;
    wire N__21436;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21412;
    wire N__21409;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21373;
    wire N__21372;
    wire N__21371;
    wire N__21370;
    wire N__21367;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21349;
    wire N__21342;
    wire N__21335;
    wire N__21332;
    wire N__21323;
    wire N__21318;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21292;
    wire N__21291;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21276;
    wire N__21273;
    wire N__21272;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21255;
    wire N__21254;
    wire N__21253;
    wire N__21252;
    wire N__21247;
    wire N__21244;
    wire N__21239;
    wire N__21234;
    wire N__21229;
    wire N__21224;
    wire N__21219;
    wire N__21204;
    wire N__21203;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21178;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21158;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21140;
    wire N__21137;
    wire N__21132;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21093;
    wire N__21090;
    wire N__21085;
    wire N__21082;
    wire N__21077;
    wire N__21074;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21047;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21004;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20975;
    wire N__20972;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20936;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20820;
    wire N__20817;
    wire N__20816;
    wire N__20815;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20803;
    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20782;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20740;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20717;
    wire N__20716;
    wire N__20713;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20650;
    wire N__20645;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20595;
    wire N__20592;
    wire N__20591;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20579;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20550;
    wire N__20547;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20454;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20392;
    wire N__20387;
    wire N__20382;
    wire N__20379;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20327;
    wire N__20322;
    wire N__20319;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20234;
    wire N__20233;
    wire N__20230;
    wire N__20229;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20125;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20102;
    wire N__20101;
    wire N__20100;
    wire N__20099;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20024;
    wire N__20021;
    wire N__20020;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19992;
    wire N__19991;
    wire N__19990;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19970;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19853;
    wire N__19852;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19805;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19747;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19577;
    wire N__19574;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19566;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19513;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19408;
    wire N__19407;
    wire N__19402;
    wire N__19397;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19367;
    wire N__19366;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19322;
    wire N__19319;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19137;
    wire N__19136;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19129;
    wire N__19120;
    wire N__19119;
    wire N__19104;
    wire N__19089;
    wire N__19088;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19075;
    wire N__19072;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19053;
    wire N__19050;
    wire N__19041;
    wire N__19040;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19005;
    wire N__19004;
    wire N__19003;
    wire N__19002;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18958;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18941;
    wire N__18940;
    wire N__18937;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18925;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18913;
    wire N__18906;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18731;
    wire N__18730;
    wire N__18727;
    wire N__18722;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18704;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18698;
    wire N__18689;
    wire N__18684;
    wire N__18683;
    wire N__18680;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18653;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18599;
    wire N__18598;
    wire N__18597;
    wire N__18596;
    wire N__18591;
    wire N__18590;
    wire N__18587;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18571;
    wire N__18566;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18530;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18506;
    wire N__18503;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18486;
    wire N__18485;
    wire N__18484;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18464;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18452;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18426;
    wire N__18425;
    wire N__18424;
    wire N__18423;
    wire N__18422;
    wire N__18421;
    wire N__18406;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18384;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18380;
    wire N__18379;
    wire N__18378;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18353;
    wire N__18350;
    wire N__18345;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18173;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18161;
    wire N__18160;
    wire N__18157;
    wire N__18156;
    wire N__18153;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18082;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18066;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18052;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18044;
    wire N__18043;
    wire N__18042;
    wire N__18041;
    wire N__18040;
    wire N__18037;
    wire N__18036;
    wire N__18033;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18015;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17979;
    wire N__17966;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17936;
    wire N__17933;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17916;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17900;
    wire N__17897;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17876;
    wire N__17873;
    wire N__17872;
    wire N__17867;
    wire N__17864;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17726;
    wire N__17721;
    wire N__17718;
    wire N__17717;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17690;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17670;
    wire N__17667;
    wire N__17666;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17636;
    wire N__17633;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17603;
    wire N__17600;
    wire N__17599;
    wire N__17594;
    wire N__17591;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17576;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17553;
    wire N__17550;
    wire N__17549;
    wire N__17546;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17522;
    wire N__17521;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17309;
    wire N__17308;
    wire N__17305;
    wire N__17300;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17264;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17225;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17210;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire \c0.n4_adj_2271_cascade_ ;
    wire \c0.n2_adj_2341 ;
    wire \c0.n2_adj_2341_cascade_ ;
    wire \c0.n10425 ;
    wire \c0.n10465 ;
    wire n10429_cascade_;
    wire n12965;
    wire n242;
    wire n12965_cascade_;
    wire n10429;
    wire n8_adj_2541;
    wire n18_adj_2539;
    wire n21_adj_2538_cascade_;
    wire n15_adj_2540;
    wire \c0.n17263 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n17265 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n17267 ;
    wire \c0.n17269 ;
    wire \c0.n17303 ;
    wire \c0.n17271 ;
    wire \c0.n17713_cascade_ ;
    wire \c0.n8_adj_2234 ;
    wire \c0.n17281 ;
    wire \c0.n17259 ;
    wire \c0.n17261 ;
    wire \c0.n13900 ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n8_adj_2257 ;
    wire \c0.n8_adj_2258 ;
    wire \c0.n39_cascade_ ;
    wire \c0.n48_adj_2383_cascade_ ;
    wire \c0.n40 ;
    wire \c0.n41 ;
    wire \c0.n43_adj_2384 ;
    wire \c0.n3_adj_2281 ;
    wire \c0.n3_adj_2322 ;
    wire \c0.n3_adj_2311 ;
    wire \c0.n3_adj_2307 ;
    wire \c0.n42 ;
    wire \c0.n3_adj_2299 ;
    wire \c0.n3_adj_2293 ;
    wire \c0.n3_adj_2297 ;
    wire \c0.n3_adj_2326 ;
    wire \c0.n3_adj_2313 ;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n49_cascade_ ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.n50_adj_2353 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.n47 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.n48 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.n17275 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n8_adj_2252 ;
    wire \c0.n8_adj_2246 ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.n17277 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.n17283 ;
    wire n17694_cascade_;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n17279 ;
    wire FRAME_MATCHER_state_31_N_1406_0_cascade_;
    wire n1166_cascade_;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n10497_cascade_ ;
    wire \c0.n17713 ;
    wire \c0.n17239 ;
    wire n15;
    wire n1437;
    wire n8_adj_2498;
    wire \c0.n6_adj_2265_cascade_ ;
    wire \c0.n18907 ;
    wire n13_adj_2469_cascade_;
    wire n7;
    wire \c0.n3_adj_2301 ;
    wire \c0.n232_cascade_ ;
    wire \c0.n6_adj_2364 ;
    wire n237;
    wire n237_cascade_;
    wire n22_adj_2465;
    wire \c0.n3_adj_2309 ;
    wire \c0.n10353_cascade_ ;
    wire \c0.n3_adj_2345 ;
    wire \c0.n3_adj_2343 ;
    wire \c0.n3 ;
    wire \c0.n3_adj_2295 ;
    wire \c0.n3_adj_2291 ;
    wire \c0.n3_adj_2289 ;
    wire \c0.n3_adj_2283 ;
    wire \c0.n3_adj_2279 ;
    wire \c0.n3_adj_2303 ;
    wire PIN_2_c_1;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n8_adj_2245 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.n17293 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n8_adj_2247 ;
    wire \c0.n10497 ;
    wire \c0.n2_adj_2315 ;
    wire \c0.n8_adj_2273_cascade_ ;
    wire \c0.n8_adj_2273 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n17273 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n17299 ;
    wire \c0.n45 ;
    wire \c0.n46_adj_2356 ;
    wire \c0.n56 ;
    wire \c0.n10513_cascade_ ;
    wire FRAME_MATCHER_i_31__N_1275;
    wire \c0.n6033_cascade_ ;
    wire \c0.n2126_cascade_ ;
    wire \c0.n27 ;
    wire \c0.n23_cascade_ ;
    wire \c0.n30_cascade_ ;
    wire \c0.n50_cascade_ ;
    wire n13849;
    wire \c0.n19_adj_2351 ;
    wire \c0.n10346 ;
    wire \c0.n17_cascade_ ;
    wire \c0.n25_adj_2352 ;
    wire \c0.n17962_cascade_ ;
    wire \c0.n4_adj_2226 ;
    wire \c0.n9575_cascade_ ;
    wire n12999;
    wire \c0.n232 ;
    wire n12999_cascade_;
    wire n18;
    wire \c0.n9575 ;
    wire n12966;
    wire n15118;
    wire FRAME_MATCHER_i_31__N_1273;
    wire \c0.n16685_cascade_ ;
    wire \c0.n6_adj_2267 ;
    wire FRAME_MATCHER_i_31__N_1270;
    wire \c0.n7528 ;
    wire \c0.n46 ;
    wire \c0.n3_adj_2332 ;
    wire \c0.n3_adj_2330 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_0 ;
    wire bfn_4_11_0_;
    wire \c0.n27_adj_2426 ;
    wire \c0.n16486 ;
    wire \c0.n115 ;
    wire \c0.n29 ;
    wire \c0.n16487 ;
    wire \c0.n16488 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_4 ;
    wire \c0.n16489 ;
    wire \c0.n16490 ;
    wire \c0.n16491 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_7 ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_7 ;
    wire \c0.n16492 ;
    wire \c0.n16493 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_8 ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_8 ;
    wire bfn_4_12_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1310_9 ;
    wire \c0.n16494 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_10 ;
    wire \c0.n16495 ;
    wire \c0.n16496 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_12 ;
    wire \c0.n16497 ;
    wire \c0.n16498 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_14 ;
    wire \c0.n16499 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_15 ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_15 ;
    wire \c0.n16500 ;
    wire \c0.n16501 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_16 ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_16 ;
    wire bfn_4_13_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1310_17 ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_17 ;
    wire \c0.n16502 ;
    wire \c0.n16503 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_19 ;
    wire \c0.n16504 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_20 ;
    wire \c0.n16505 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_21 ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_21 ;
    wire \c0.n16506 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_22 ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_22 ;
    wire \c0.n16507 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_23 ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_23 ;
    wire \c0.n16508 ;
    wire \c0.n16509 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_24 ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_24 ;
    wire bfn_4_14_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1310_25 ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_25 ;
    wire \c0.n16510 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_26 ;
    wire \c0.n16511 ;
    wire \c0.n16512 ;
    wire \c0.n16513 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_29 ;
    wire \c0.n16514 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_30 ;
    wire \c0.n16515 ;
    wire \c0.n16516 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_31 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_9 ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire \c0.n3_adj_2328 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_6 ;
    wire \c0.n3_adj_2334 ;
    wire \control.n18909 ;
    wire \c0.n8_adj_2254 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.n8_adj_2250 ;
    wire \c0.n4_adj_2271 ;
    wire \c0.n8_adj_2249 ;
    wire \c0.n4_adj_2349 ;
    wire \c0.n8_adj_2244 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n30_adj_2355_cascade_ ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n51 ;
    wire \c0.n10613_cascade_ ;
    wire \c0.n22_adj_2346 ;
    wire data_in_frame_5_6;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.n2126 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.n2137_adj_2237 ;
    wire \c0.n2137_adj_2237_cascade_ ;
    wire data_in_frame_2_0;
    wire data_in_frame_2_5;
    wire n16802_cascade_;
    wire \c0.n10569_cascade_ ;
    wire data_in_frame_0_1;
    wire \c0.rx.r_Rx_Data_R ;
    wire n11058_cascade_;
    wire \c0.FRAME_MATCHER_i_31_N_1310_3 ;
    wire \c0.n1502 ;
    wire \c0.n1502_cascade_ ;
    wire \c0.n10522 ;
    wire \c0.n4_adj_2266 ;
    wire \c0.n13033_cascade_ ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_30 ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_29 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_28 ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_19 ;
    wire FRAME_MATCHER_i_31;
    wire \c0.FRAME_MATCHER_i_31_N_1310_31 ;
    wire n63_adj_2534_cascade_;
    wire \c0.FRAME_MATCHER_i_31_N_1310_18 ;
    wire \c0.n63_adj_2262_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_5 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_5 ;
    wire \c0.n3_adj_2336 ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire \c0.n10_adj_2378 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_4 ;
    wire \c0.n7199 ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire \c0.n10353 ;
    wire \c0.n3_adj_2338 ;
    wire n63;
    wire \c0.n63_adj_2262 ;
    wire n63_adj_2534;
    wire \c0.n113 ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_14 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_13 ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_10 ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_6 ;
    wire \c0.n109 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_11 ;
    wire \c0.n3_adj_2324 ;
    wire \c0.n26_adj_2379_cascade_ ;
    wire \c0.n44_adj_2382 ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_11 ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_20 ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_12 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_27 ;
    wire \c0.n13033 ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_26 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_27 ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire \c0.n3_adj_2287 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_3 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.n3_adj_2340 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_28 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.n3_adj_2285 ;
    wire n18043;
    wire n18044;
    wire LED_c;
    wire PIN_3_c_2;
    wire \c0.n4_adj_2225 ;
    wire tx2_o;
    wire tx2_enable;
    wire \c0.n4_adj_2216 ;
    wire \c0.data_in_frame_3_3 ;
    wire data_in_frame_2_2;
    wire \c0.n18_adj_2417 ;
    wire data_in_frame_2_1;
    wire \c0.n21_adj_2421 ;
    wire \c0.n24_adj_2418 ;
    wire \c0.n23_adj_2420_cascade_ ;
    wire n16797_cascade_;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.rx.n129_cascade_ ;
    wire \c0.data_in_frame_3_7 ;
    wire data_in_frame_6_1;
    wire data_in_frame_6_7;
    wire \c0.n17813 ;
    wire \c0.n10761 ;
    wire data_in_frame_0_0;
    wire \c0.n10761_cascade_ ;
    wire \c0.data_in_frame_1_5 ;
    wire \c0.n17733_cascade_ ;
    wire data_in_frame_6_0;
    wire \c0.n17735 ;
    wire \c0.data_in_frame_1_6 ;
    wire \c0.n17733 ;
    wire \c0.n10569 ;
    wire data_in_frame_6_3;
    wire \c0.n17734_cascade_ ;
    wire \c0.data_in_frame_1_7 ;
    wire \c0.n19_adj_2400 ;
    wire \c0.n18_adj_2398 ;
    wire \c0.n18000_cascade_ ;
    wire data_in_frame_5_2;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire \c0.rx.n12963 ;
    wire n120_cascade_;
    wire data_in_frame_2_3;
    wire data_in_frame_0_4;
    wire data_in_frame_0_5;
    wire data_in_frame_2_6;
    wire \c0.n15_adj_2416 ;
    wire \c0.n2138 ;
    wire \c0.n22_adj_2419 ;
    wire data_in_frame_5_7;
    wire data_in_frame_2_7;
    wire \c0.rx.n17702_cascade_ ;
    wire \c0.rx.n17702 ;
    wire \c0.rx.n17704_cascade_ ;
    wire n11058;
    wire n16802;
    wire \c0.n18002_cascade_ ;
    wire \c0.n10498 ;
    wire \c0.rx.n10988_cascade_ ;
    wire \c0.rx.n12624_cascade_ ;
    wire data_in_0_2;
    wire \c0.n20_adj_2371_cascade_ ;
    wire \c0.n10516 ;
    wire \c0.n10516_cascade_ ;
    wire \c0.n10367 ;
    wire data_in_0_5;
    wire \c0.n10367_cascade_ ;
    wire \c0.n15_adj_2389 ;
    wire data_in_1_4;
    wire data_in_0_4;
    wire data_in_3_4;
    wire \c0.n14_adj_2388 ;
    wire \c0.n18631 ;
    wire data_in_1_5;
    wire data_in_2_4;
    wire \c0.n18_adj_2370 ;
    wire \c0.n13_adj_2380 ;
    wire \c0.rx.n10988 ;
    wire \c0.n18006_cascade_ ;
    wire \c0.n14_adj_2375 ;
    wire data_in_2_7;
    wire data_in_2_5;
    wire rx_data_7;
    wire bfn_6_13_0_;
    wire \c0.rx.n16532 ;
    wire \c0.rx.n16533 ;
    wire \c0.rx.n16534 ;
    wire \c0.rx.n16535 ;
    wire \c0.rx.n16536 ;
    wire \c0.rx.n16537 ;
    wire \c0.rx.n16538 ;
    wire \c0.rx.n12819 ;
    wire \c0.n18225_cascade_ ;
    wire \c0.rx.n5 ;
    wire \c0.rx.n57 ;
    wire \c0.rx.n15905_cascade_ ;
    wire \c0.rx.n6_cascade_ ;
    wire \c0.rx.n12 ;
    wire \c0.rx.n12_cascade_ ;
    wire \c0.rx.n11082 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_18 ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire \c0.n3_adj_2305 ;
    wire n1166;
    wire \c0.FRAME_MATCHER_i_31_N_1278_13 ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.n3_adj_2317 ;
    wire n26;
    wire bfn_6_21_0_;
    wire n25;
    wire n16609;
    wire n24;
    wire n16610;
    wire n23;
    wire n16611;
    wire n22_adj_2481;
    wire n16612;
    wire n21;
    wire n16613;
    wire n20;
    wire n16614;
    wire n19;
    wire n16615;
    wire n16616;
    wire n18_adj_2480;
    wire bfn_6_22_0_;
    wire n17;
    wire n16617;
    wire n16;
    wire n16618;
    wire n15_adj_2479;
    wire n16619;
    wire n14_adj_2478;
    wire n16620;
    wire n13;
    wire n16621;
    wire n12;
    wire n16622;
    wire n11;
    wire n16623;
    wire n16624;
    wire n10_adj_2467;
    wire bfn_6_23_0_;
    wire n9;
    wire n16625;
    wire n8;
    wire n16626;
    wire n7_adj_2476;
    wire n16627;
    wire n6;
    wire n16628;
    wire blink_counter_21;
    wire n16629;
    wire blink_counter_22;
    wire n16630;
    wire blink_counter_23;
    wire n16631;
    wire n16632;
    wire blink_counter_24;
    wire bfn_6_24_0_;
    wire n16633;
    wire blink_counter_25;
    wire \control.n11 ;
    wire PIN_1_c_0;
    wire \c0.n13808_cascade_ ;
    wire \c0.n14064_cascade_ ;
    wire \c0.n4_adj_2203 ;
    wire \c0.n4_adj_2201 ;
    wire n17694;
    wire \c0.n43 ;
    wire \c0.n4_adj_2199 ;
    wire bfn_7_3_0_;
    wire \c0.n18253 ;
    wire \c0.n16479 ;
    wire \c0.n18314 ;
    wire \c0.n16480 ;
    wire \c0.n18315 ;
    wire \c0.n16481 ;
    wire \c0.n16482 ;
    wire \c0.byte_transmit_counter2_5 ;
    wire \c0.n18316 ;
    wire \c0.n16483 ;
    wire \c0.byte_transmit_counter2_6 ;
    wire \c0.n18317 ;
    wire \c0.n16484 ;
    wire \c0.byte_transmit_counter2_7 ;
    wire \c0.tx2_transmit_N_1996 ;
    wire \c0.n16485 ;
    wire \c0.n18318 ;
    wire \c0.n18100_cascade_ ;
    wire \c0.n18103_cascade_ ;
    wire \c0.n2122 ;
    wire data_in_frame_6_5;
    wire \c0.n16994 ;
    wire \c0.data_in_frame_3_2 ;
    wire data_in_frame_6_6;
    wire data_in_frame_5_1;
    wire data_in_frame_6_2;
    wire n16797;
    wire data_in_frame_5_4;
    wire n158;
    wire n12600;
    wire rx_data_3;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire \c0.rx.n129 ;
    wire data_in_frame_5_3;
    wire \c0.data_in_frame_1_2 ;
    wire data_in_frame_5_5;
    wire \c0.data_in_frame_1_3 ;
    wire \c0.n16981_cascade_ ;
    wire \c0.n20_adj_2397 ;
    wire \c0.n20_adj_2350 ;
    wire \c0.n2128 ;
    wire data_in_frame_6_4;
    wire data_in_frame_5_0;
    wire \c0.n2128_cascade_ ;
    wire \c0.n22_adj_2392 ;
    wire data_in_frame_0_2;
    wire data_in_frame_0_3;
    wire \c0.n2120 ;
    wire \c0.n2124 ;
    wire \c0.data_in_frame_3_4 ;
    wire \c0.n2120_cascade_ ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.n19_adj_2415 ;
    wire \c0.data_in_frame_1_0 ;
    wire \c0.data_in_frame_1_1 ;
    wire data_in_frame_0_7;
    wire \c0.data_in_frame_1_4 ;
    wire \c0.n17721_cascade_ ;
    wire data_in_frame_0_6;
    wire \c0.n10_adj_2390 ;
    wire rx_data_4;
    wire n120;
    wire data_in_frame_2_4;
    wire \c0.rx.n18729_cascade_ ;
    wire \c0.rx.n18732_cascade_ ;
    wire \c0.rx.n11 ;
    wire n12582;
    wire n135_adj_2463;
    wire n4_adj_2471_cascade_;
    wire data_in_1_0;
    wire \c0.rx.n110 ;
    wire rx_data_2;
    wire \c0.rx.r_SM_Main_2_N_2088_2_cascade_ ;
    wire \c0.rx.n161 ;
    wire rx_data_0;
    wire data_in_3_2;
    wire data_in_0_6;
    wire data_in_3_6;
    wire \c0.n8_adj_2385 ;
    wire \c0.n15_adj_2372 ;
    wire data_in_1_2;
    wire data_in_0_7;
    wire \c0.rx.r_Bit_Index_0 ;
    wire n151;
    wire n151_cascade_;
    wire data_in_2_2;
    wire \c0.n18008 ;
    wire \c0.n8_adj_2369_cascade_ ;
    wire \c0.n10493 ;
    wire data_in_2_6;
    wire data_in_1_6;
    wire \c0.rx.n18304 ;
    wire rx_data_5;
    wire data_in_3_5;
    wire rx_data_1;
    wire data_in_3_0;
    wire data_in_2_0;
    wire data_in_1_7;
    wire \c0.n13693 ;
    wire \c0.rx.r_SM_Main_2_N_2088_2 ;
    wire \c0.rx.n11041_cascade_ ;
    wire \c0.rx.r_Bit_Index_2 ;
    wire \c0.rx.n167 ;
    wire n12527;
    wire data_in_0_0;
    wire data_in_3_7;
    wire \c0.n6_adj_2368 ;
    wire data_in_1_3;
    wire data_in_0_3;
    wire data_in_0_1;
    wire \c0.rx.n18196 ;
    wire \c0.rx.n18194 ;
    wire \c0.rx.n12552_cascade_ ;
    wire rx_data_6;
    wire \c0.rx.r_Bit_Index_1 ;
    wire \c0.rx.r_SM_Main_2 ;
    wire n164_adj_2464;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n17990_cascade_ ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.n18024_cascade_ ;
    wire \c0.rx.n12828 ;
    wire \c0.rx.n12828_cascade_ ;
    wire \c0.rx.n18303 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n15902 ;
    wire \c0.rx.r_Clock_Count_0 ;
    wire \c0.rx.n18211 ;
    wire \c0.rx.r_SM_Main_1 ;
    wire r_Rx_Data;
    wire \c0.rx.r_SM_Main_0 ;
    wire \c0.rx.n4 ;
    wire \c0.tx.n54_cascade_ ;
    wire \c0.tx.n10 ;
    wire \c0.tx.n54 ;
    wire \c0.tx.n47_cascade_ ;
    wire \c0.tx.r_Clock_Count_0 ;
    wire bfn_7_15_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n16524 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n16525 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n16526 ;
    wire \c0.tx.r_Clock_Count_4 ;
    wire \c0.tx.n16527 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire \c0.tx.n16528 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.n16529 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.n16530 ;
    wire \c0.tx.n16531 ;
    wire bfn_7_16_0_;
    wire \c0.tx.r_Clock_Count_8 ;
    wire \c0.tx.n11297 ;
    wire \control.n8 ;
    wire \control.PHASES_5_N_2152_1_cascade_ ;
    wire \control.n10356 ;
    wire \c0.n18801_cascade_ ;
    wire \c0.n18804 ;
    wire \c0.n18843 ;
    wire \c0.n18846_cascade_ ;
    wire \c0.n22_adj_2239 ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire \c0.n18675_cascade_ ;
    wire \c0.n18678_cascade_ ;
    wire \c0.n18741_cascade_ ;
    wire \c0.n22_adj_2242 ;
    wire \c0.n18744_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire n17689_cascade_;
    wire \c0.n18684 ;
    wire \c0.n18072 ;
    wire \c0.tx2.n14_cascade_ ;
    wire \c0.n18284_cascade_ ;
    wire \c0.n27_adj_2405 ;
    wire \c0.n29_adj_2408 ;
    wire \c0.n12704_cascade_ ;
    wire \c0.n18287 ;
    wire n612;
    wire \c0.n18289_cascade_ ;
    wire \c0.n18831 ;
    wire \c0.n18079_cascade_ ;
    wire \c0.n17725 ;
    wire \c0.n16863 ;
    wire \c0.n16982 ;
    wire \c0.n17722 ;
    wire \c0.n28_adj_2403 ;
    wire \c0.n6033 ;
    wire \c0.n18085_cascade_ ;
    wire \c0.n4494 ;
    wire \c0.n28 ;
    wire \c0.n12704 ;
    wire \c0.n18082 ;
    wire \c0.n18270 ;
    wire \c0.n6035 ;
    wire bfn_9_6_0_;
    wire \c0.tx2.n16539 ;
    wire \c0.tx2.n16540 ;
    wire \c0.tx2.n16541 ;
    wire \c0.tx2.n16542 ;
    wire \c0.tx2.n16543 ;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire \c0.tx2.n16544 ;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire \c0.tx2.n16545 ;
    wire \c0.tx2.n16546 ;
    wire bfn_9_7_0_;
    wire \c0.tx2.r_Clock_Count_8 ;
    wire \c0.tx2.n11312 ;
    wire bfn_9_8_0_;
    wire \c0.n16517 ;
    wire \c0.n16518 ;
    wire \c0.n16519 ;
    wire \c0.n16520 ;
    wire \c0.n16521 ;
    wire \c0.n16522 ;
    wire \c0.n16523 ;
    wire \c0.n18254 ;
    wire \c0.n4_adj_2231 ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.n73 ;
    wire \c0.n44 ;
    wire tx_enable;
    wire \c0.tx_active_prev ;
    wire data_in_1_1;
    wire n3_adj_2525_cascade_;
    wire tx_o;
    wire \c0.tx.n17697 ;
    wire data_out_1_7;
    wire \c0.tx.n11030_cascade_ ;
    wire \c0.tx.n18041 ;
    wire \c0.tx.o_Tx_Serial_N_2062 ;
    wire n18750;
    wire n10_adj_2532_cascade_;
    wire r_Tx_Data_6;
    wire \c0.tx.n17984 ;
    wire n10_adj_2537_cascade_;
    wire n10_adj_2535_cascade_;
    wire r_Tx_Data_7;
    wire \c0.n18188 ;
    wire n5155;
    wire \c0.n18354 ;
    wire n18756;
    wire \c0.data_out_3_6 ;
    wire data_out_3_7;
    wire data_out_2_7;
    wire \c0.n2_adj_2229 ;
    wire n2837_cascade_;
    wire data_out_0_5;
    wire \control.n12_cascade_ ;
    wire \control.n10 ;
    wire bfn_9_23_0_;
    wire \control.n9_adj_2459 ;
    wire \control.n16647 ;
    wire \control.pwm_delay_2 ;
    wire \control.n16648 ;
    wire \control.pwm_delay_3 ;
    wire \control.n16649 ;
    wire \control.pwm_delay_4 ;
    wire \control.n16650 ;
    wire \control.pwm_delay_5 ;
    wire \control.n16651 ;
    wire \control.pwm_delay_6 ;
    wire \control.n16652 ;
    wire \control.pwm_delay_7 ;
    wire \control.n16653 ;
    wire \control.n16654 ;
    wire \control.pwm_delay_8 ;
    wire bfn_9_24_0_;
    wire \control.n16655 ;
    wire \c0.n18888_cascade_ ;
    wire \c0.n18789_cascade_ ;
    wire \c0.n18792_cascade_ ;
    wire \c0.n22_adj_2270 ;
    wire \c0.n18885 ;
    wire \c0.n10861_cascade_ ;
    wire \c0.n18798 ;
    wire \c0.n10893_cascade_ ;
    wire data_out_frame2_17_1;
    wire \c0.n5_adj_2435_cascade_ ;
    wire \c0.n6_adj_2223 ;
    wire \c0.n18687_cascade_ ;
    wire \c0.n18690 ;
    wire \c0.n5_adj_2197 ;
    wire \c0.n6 ;
    wire \c0.n6_adj_2354 ;
    wire \c0.n18855 ;
    wire tx2_active;
    wire \c0.n14064 ;
    wire \c0.n12359_cascade_ ;
    wire \c0.n6_adj_2443_cascade_ ;
    wire \c0.n10513 ;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n10958 ;
    wire \c0.r_SM_Main_2_N_2034_0_adj_2213 ;
    wire n6707;
    wire \c0.tx2.n12769 ;
    wire r_SM_Main_2_N_2031_1;
    wire r_SM_Main_2_N_2031_1_cascade_;
    wire n18014_cascade_;
    wire \c0.n18362 ;
    wire \c0.n12359 ;
    wire FRAME_MATCHER_i_31__N_1272;
    wire \c0.n4_adj_2204 ;
    wire \c0.tx2.n13800 ;
    wire r_SM_Main_1;
    wire r_SM_Main_0;
    wire n3;
    wire \c0.tx2.n18164 ;
    wire \c0.tx2.n18163 ;
    wire \c0.tx2.n18062 ;
    wire \c0.tx2.n18717_cascade_ ;
    wire \c0.tx2.o_Tx_Serial_N_2062 ;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire \c0.tx2.n10 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire \c0.tx2.n10_cascade_ ;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire \c0.tx2.n12775 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.n18061 ;
    wire r_SM_Main_2;
    wire n11096;
    wire \c0.n18260_cascade_ ;
    wire \c0.n130 ;
    wire \c0.n3465 ;
    wire \c0.n4806 ;
    wire byte_transmit_counter_6;
    wire tx_transmit_N_1947_6;
    wire tx_transmit_N_1947_4;
    wire \c0.n4_cascade_ ;
    wire n5341_cascade_;
    wire tx_transmit_N_1947_7;
    wire byte_transmit_counter_7;
    wire \c0.tx_transmit_N_1947_5 ;
    wire n10973;
    wire n5341;
    wire \c0.byte_transmit_counter_5 ;
    wire \c0.n17998 ;
    wire \c0.tx.n17938 ;
    wire n10_adj_2536;
    wire n5440_cascade_;
    wire n18016;
    wire n18016_cascade_;
    wire \c0.n8_adj_2207 ;
    wire \c0.tx.n13802 ;
    wire \c0.tx.n13802_cascade_ ;
    wire \c0.tx.n6796_cascade_ ;
    wire r_Bit_Index_1;
    wire \c0.tx.n18167 ;
    wire r_Bit_Index_2;
    wire \c0.tx.n18711 ;
    wire r_Tx_Data_1;
    wire \c0.tx.n18040 ;
    wire \c0.n8_adj_2205 ;
    wire \c0.tx.r_SM_Main_2 ;
    wire \c0.tx.r_SM_Main_0 ;
    wire \c0.tx.r_SM_Main_1 ;
    wire \c0.tx.r_SM_Main_2_N_2031_1 ;
    wire n18012;
    wire r_Bit_Index_0;
    wire r_Tx_Data_5;
    wire \c0.tx.n18166 ;
    wire \c0.n5_adj_2241 ;
    wire \c0.n18753 ;
    wire \c0.n2 ;
    wire \c0.n18189 ;
    wire n18876_cascade_;
    wire n10_adj_2531;
    wire \c0.n5_adj_2196_cascade_ ;
    wire \c0.n18873 ;
    wire n5_cascade_;
    wire \c0.n8_adj_2209 ;
    wire n10_adj_2533;
    wire n10_adj_2528_cascade_;
    wire r_Tx_Data_2;
    wire data_out_3_5;
    wire data_out_1_6;
    wire \c0.data_out_0_6 ;
    wire \c0.n1_adj_2272 ;
    wire data_out_2_5;
    wire \c0.n18335 ;
    wire \c0.data_out_2_3 ;
    wire \c0.n19_cascade_ ;
    wire \c0.data_out_frame2_19_1 ;
    wire \c0.n20 ;
    wire \c0.n18266 ;
    wire \c0.n18360 ;
    wire \c0.n18256 ;
    wire \c0.n14_adj_2359_cascade_ ;
    wire \c0.data_out_frame2_20_0 ;
    wire \c0.n15_adj_2429 ;
    wire \c0.n17847 ;
    wire \c0.n10867_cascade_ ;
    wire \c0.n17739_cascade_ ;
    wire data_out_frame2_17_0;
    wire \c0.n18840 ;
    wire \c0.n18795 ;
    wire data_out_frame2_18_7;
    wire data_out_frame2_5_1;
    wire \c0.n18837 ;
    wire data_out_frame2_18_1;
    wire data_out_frame2_17_7;
    wire \c0.n17727 ;
    wire data_out_frame2_7_1;
    wire bfn_11_7_0_;
    wire \c0.n16634 ;
    wire \c0.n16635 ;
    wire \c0.n16636 ;
    wire \c0.n16637 ;
    wire \c0.n16638 ;
    wire \c0.n16639 ;
    wire \c0.n16640 ;
    wire \c0.n16641 ;
    wire bfn_11_8_0_;
    wire \c0.n16642 ;
    wire \c0.n16643 ;
    wire \c0.n16644 ;
    wire \c0.n16645 ;
    wire \c0.n16646 ;
    wire \c0.delay_counter_2 ;
    wire \c0.delay_counter_5 ;
    wire n26_adj_2466;
    wire \c0.n18019 ;
    wire n129;
    wire \c0.r_SM_Main_2_N_2034_0 ;
    wire n129_cascade_;
    wire \c0.tx_active ;
    wire \c0.n1707 ;
    wire \c0.delay_counter_11 ;
    wire \c0.delay_counter_12 ;
    wire \c0.delay_counter_4 ;
    wire \c0.delay_counter_7 ;
    wire \c0.n24 ;
    wire n12227;
    wire n574_cascade_;
    wire \c0.n98 ;
    wire \c0.n18230 ;
    wire n17978_cascade_;
    wire UART_TRANSMITTER_state_7_N_1223_1;
    wire n18202;
    wire n574;
    wire n4;
    wire n22_adj_2522;
    wire \c0.n18226 ;
    wire n21_adj_2524;
    wire n6_adj_2470;
    wire n18368;
    wire \c0.n18861_cascade_ ;
    wire \c0.n18377 ;
    wire n18864_cascade_;
    wire n10_adj_2529_cascade_;
    wire r_Tx_Data_3;
    wire n10_adj_2499;
    wire \c0.n10550_cascade_ ;
    wire \c0.n10524 ;
    wire \c0.n10550 ;
    wire \c0.n10746 ;
    wire \c0.n6_adj_2361 ;
    wire \c0.n10746_cascade_ ;
    wire n17758_cascade_;
    wire \c0.n10734 ;
    wire \c0.n8_adj_2232 ;
    wire n10_adj_2461;
    wire data_out_8_7;
    wire \c0.n17742_cascade_ ;
    wire \c0.n17742 ;
    wire \c0.n10558 ;
    wire \c0.data_out_9_5 ;
    wire \c0.n6_adj_2365_cascade_ ;
    wire \c0.n5_adj_2220 ;
    wire r_Tx_Data_4;
    wire \c0.n18265 ;
    wire n9667;
    wire byte_transmit_counter_4;
    wire r_Tx_Data_0;
    wire \c0.n1_cascade_ ;
    wire n22;
    wire \c0.n18849 ;
    wire n18852_cascade_;
    wire n10;
    wire \c0.n18264 ;
    wire \c0.n8 ;
    wire n10_adj_2527;
    wire \c0.n18322 ;
    wire data_out_0_1;
    wire n11017_cascade_;
    wire data_out_0_0;
    wire data_out_3_4;
    wire \control.PHASES_5_N_2152_1 ;
    wire \control.pwm_delay_9 ;
    wire \control.n18 ;
    wire \control.n17926 ;
    wire \control.PHASES_5__N_2160_cascade_ ;
    wire \control.n5 ;
    wire \control.n17950 ;
    wire \control.n9 ;
    wire \c0.n18639_cascade_ ;
    wire \c0.n10700_cascade_ ;
    wire \c0.n21 ;
    wire \c0.n17804 ;
    wire \c0.n17874 ;
    wire \c0.n17908 ;
    wire \c0.n18_adj_2423 ;
    wire \c0.n17908_cascade_ ;
    wire \c0.n28_adj_2425 ;
    wire \c0.n30_adj_2424_cascade_ ;
    wire \c0.n29_adj_2427 ;
    wire data_out_frame2_17_5;
    wire data_out_frame2_12_1;
    wire \c0.n10829_cascade_ ;
    wire \c0.FRAME_MATCHER_state_1 ;
    wire \c0.n14161 ;
    wire \c0.FRAME_MATCHER_state_2 ;
    wire \c0.n50 ;
    wire n11114_cascade_;
    wire data_out_frame2_18_0;
    wire data_out_frame2_6_7;
    wire \c0.delay_counter_10 ;
    wire \c0.delay_counter_0 ;
    wire \c0.delay_counter_13 ;
    wire \c0.delay_counter_6 ;
    wire \c0.n18810 ;
    wire \c0.tx_transmit_N_1947_0 ;
    wire \c0.tx_transmit_N_1947_1 ;
    wire \c0.tx_transmit_N_1947_2 ;
    wire \c0.n155 ;
    wire \c0.delay_counter_9 ;
    wire \c0.delay_counter_1 ;
    wire \c0.n22 ;
    wire n25_adj_2468;
    wire \c0.n18807 ;
    wire \c0.n5_adj_2436 ;
    wire r_Bit_Index_0_adj_2519;
    wire r_Bit_Index_1_adj_2518;
    wire tx_transmit_N_1947_3;
    wire \c0.n85 ;
    wire \c0.n14068 ;
    wire \c0.n18259 ;
    wire n18014;
    wire n4_adj_2472;
    wire n11545;
    wire r_Bit_Index_2_adj_2517;
    wire \c0.n17715 ;
    wire \c0.delay_counter_3 ;
    wire \c0.delay_counter_8 ;
    wire \c0.n18 ;
    wire data_in_3_1;
    wire data_in_2_1;
    wire data_in_3_3;
    wire rx_data_ready;
    wire data_in_2_3;
    wire \c0.n18365 ;
    wire data_out_frame2_18_5;
    wire n1;
    wire n24_adj_2523;
    wire n18_adj_2526;
    wire \c0.n17761_cascade_ ;
    wire n9_adj_2477;
    wire \c0.n17761 ;
    wire \c0.n18747 ;
    wire \c0.n17807_cascade_ ;
    wire data_out_9_2;
    wire \c0.n6_adj_2318_cascade_ ;
    wire \c0.data_out_9_0 ;
    wire \c0.data_out_9_6 ;
    wire \c0.n6_adj_2367 ;
    wire \c0.n17850 ;
    wire \c0.n10749 ;
    wire \c0.data_out_9__2__N_367_cascade_ ;
    wire \c0.n15_adj_2319_cascade_ ;
    wire \c0.n14_adj_2320 ;
    wire \c0.data_out_10_2 ;
    wire \c0.n17826 ;
    wire \c0.data_out_9_7 ;
    wire \c0.n17774 ;
    wire \c0.n17774_cascade_ ;
    wire \c0.data_out_10_3 ;
    wire \c0.data_out_10_5 ;
    wire \c0.n6_adj_2314 ;
    wire \c0.n17883 ;
    wire \c0.n10801_cascade_ ;
    wire \c0.data_out_10_0 ;
    wire \c0.n17768 ;
    wire \c0.n10_adj_2366_cascade_ ;
    wire \c0.data_out_10_1 ;
    wire \c0.data_out_6_1 ;
    wire \c0.n17819 ;
    wire \c0.n6_adj_2277 ;
    wire \c0.data_out_9_4 ;
    wire \c0.n8_adj_2211_cascade_ ;
    wire \c0.n18222_cascade_ ;
    wire \c0.n18693_cascade_ ;
    wire n18696;
    wire \c0.data_out_6_2 ;
    wire \c0.n5_adj_2347 ;
    wire byte_transmit_counter_1;
    wire \c0.n18191 ;
    wire \c0.n18867_cascade_ ;
    wire byte_transmit_counter_2;
    wire n10_adj_2505;
    wire n18870_cascade_;
    wire byte_transmit_counter_3;
    wire n10_adj_2530;
    wire \c0.n5_adj_2214 ;
    wire \c0.data_out_1_4 ;
    wire \c0.n18190 ;
    wire \c0.n2_adj_2348 ;
    wire \c0.n18334 ;
    wire \c0.data_out_7_4 ;
    wire data_out_3_2;
    wire \c0.data_out_1_2 ;
    wire \c0.n18223 ;
    wire data_out_2_2;
    wire PIN_24_c_3;
    wire \control.n6 ;
    wire \control.n17251 ;
    wire PIN_23_c_4;
    wire \control.n6_adj_2460 ;
    wire \control.n10490 ;
    wire hall3;
    wire hall2;
    wire hall1;
    wire \control.PHASES_5__N_2160 ;
    wire \control.PHASES_5_N_2130_5 ;
    wire \c0.n17748 ;
    wire data_out_frame2_15_1;
    wire \c0.n10829 ;
    wire \c0.n10890_cascade_ ;
    wire \c0.n17_adj_2449 ;
    wire \c0.n16_adj_2448_cascade_ ;
    wire \c0.n17911 ;
    wire \c0.n15_adj_2445 ;
    wire \c0.n14_adj_2444_cascade_ ;
    wire data_out_frame2_16_1;
    wire \c0.data_out_frame2_20_5 ;
    wire \c0.n16_adj_2358 ;
    wire \c0.n10720_cascade_ ;
    wire data_out_frame2_10_2;
    wire \c0.n10819 ;
    wire \c0.n17886 ;
    wire \c0.n20_adj_2442 ;
    wire \c0.n16_cascade_ ;
    wire \c0.n17795 ;
    wire \c0.data_out_frame2_19_5 ;
    wire \c0.n10839 ;
    wire \c0.n10890 ;
    wire data_out_frame2_10_5;
    wire \c0.n10816 ;
    wire \c0.n12_adj_2446_cascade_ ;
    wire data_out_frame2_6_4;
    wire \c0.n10864 ;
    wire \c0.n10_adj_2440 ;
    wire \c0.n6_adj_2357 ;
    wire \c0.n18879_cascade_ ;
    wire \c0.n10852 ;
    wire \c0.n10867 ;
    wire data_out_frame2_8_5;
    wire \c0.n14_adj_2447 ;
    wire \c0.data_out_frame2_19_4 ;
    wire data_out_frame2_15_3;
    wire \c0.n6_adj_2422_cascade_ ;
    wire data_out_frame2_18_4;
    wire \c0.n10870_cascade_ ;
    wire \c0.n27_adj_2428 ;
    wire \c0.n5_adj_2274 ;
    wire data_out_8_2;
    wire \c0.n11056 ;
    wire \c0.n18199_cascade_ ;
    wire \c0.n17832 ;
    wire \c0.n18242_cascade_ ;
    wire \c0.data_out_6_6 ;
    wire \c0.n5 ;
    wire \c0.n18247 ;
    wire \c0.n18238_cascade_ ;
    wire \c0.data_out_6_4 ;
    wire \c0.n6_adj_2276 ;
    wire \c0.data_out_6_7 ;
    wire \c0.data_out_6_5 ;
    wire data_out_8_4;
    wire \c0.n17745 ;
    wire \c0.n10542 ;
    wire \c0.n17745_cascade_ ;
    wire \c0.data_out_10_7 ;
    wire data_out_8_3;
    wire \c0.n8_adj_2219 ;
    wire data_out_0_3;
    wire \c0.n18376 ;
    wire data_out_10_6;
    wire \c0.data_out_7_2 ;
    wire \c0.data_out_9_1 ;
    wire \c0.n17730 ;
    wire \c0.n17835 ;
    wire \c0.n17844 ;
    wire \c0.n17730_cascade_ ;
    wire n17758;
    wire \c0.n14_adj_2363_cascade_ ;
    wire \c0.n13 ;
    wire \c0.data_out_9_3 ;
    wire \c0.n17816_cascade_ ;
    wire \c0.n17877 ;
    wire \c0.n12 ;
    wire \c0.n17786 ;
    wire \c0.n18184 ;
    wire \c0.data_out_7_1 ;
    wire \c0.n10537 ;
    wire data_out_6_0;
    wire \c0.n10680 ;
    wire \c0.n17816 ;
    wire \c0.n10680_cascade_ ;
    wire \c0.data_out_5_5 ;
    wire data_out_8_6;
    wire data_out_8_5;
    wire \c0.n17771 ;
    wire data_out_5_1;
    wire \c0.data_out_5_4 ;
    wire data_out_frame2_13_2;
    wire data_out_frame2_16_0;
    wire data_out_frame2_8_6;
    wire \c0.n18759_cascade_ ;
    wire data_out_frame2_6_0;
    wire \c0.n10920 ;
    wire \c0.n17783_cascade_ ;
    wire \c0.n10849 ;
    wire \c0.n17859 ;
    wire \c0.n15_cascade_ ;
    wire \c0.data_out_frame2_19_0 ;
    wire \c0.n10688 ;
    wire \c0.n10813_cascade_ ;
    wire \c0.n10577 ;
    wire \c0.n17783 ;
    wire \c0.n15_adj_2414_cascade_ ;
    wire \c0.data_out_frame2_20_1 ;
    wire \c0.n31 ;
    wire \c0.n32_cascade_ ;
    wire \c0.data_out_frame2_19_7 ;
    wire \c0.data_out_frame2_0_7 ;
    wire \c0.n17777 ;
    wire \c0.n6_adj_2430 ;
    wire \c0.n17777_cascade_ ;
    wire data_out_frame2_5_5;
    wire \c0.n10617_cascade_ ;
    wire \c0.n17765 ;
    wire \c0.data_out_frame2_0_4 ;
    wire \c0.n18681 ;
    wire bfn_14_5_0_;
    wire n16547;
    wire n16548;
    wire n16549;
    wire n16550;
    wire n16551;
    wire n16552;
    wire n16553;
    wire n16554;
    wire bfn_14_6_0_;
    wire n16555;
    wire n16556;
    wire n16557;
    wire n16558;
    wire n16559;
    wire n16560;
    wire n16561;
    wire n16562;
    wire bfn_14_7_0_;
    wire n16563;
    wire n16564;
    wire n16565;
    wire n16566;
    wire n16567;
    wire n16568;
    wire n16569;
    wire n16570;
    wire bfn_14_8_0_;
    wire n16571;
    wire n16572;
    wire n16573;
    wire n16574;
    wire n16575;
    wire n16576;
    wire n16577;
    wire rand_data_0;
    wire bfn_14_9_0_;
    wire rand_data_1;
    wire n16578;
    wire rand_data_2;
    wire rand_setpoint_2;
    wire n16579;
    wire rand_data_3;
    wire rand_setpoint_3;
    wire n16580;
    wire rand_data_4;
    wire rand_setpoint_4;
    wire n16581;
    wire rand_setpoint_5;
    wire n16582;
    wire rand_setpoint_6;
    wire n16583;
    wire rand_setpoint_7;
    wire n16584;
    wire n16585;
    wire rand_data_8;
    wire bfn_14_10_0_;
    wire rand_data_9;
    wire rand_setpoint_9;
    wire n16586;
    wire rand_data_10;
    wire rand_setpoint_10;
    wire n16587;
    wire n16588;
    wire rand_setpoint_12;
    wire n16589;
    wire rand_data_13;
    wire n16590;
    wire rand_data_14;
    wire n16591;
    wire rand_data_15;
    wire rand_setpoint_15;
    wire n16592;
    wire n16593;
    wire rand_data_16;
    wire rand_setpoint_16;
    wire bfn_14_11_0_;
    wire rand_data_17;
    wire rand_setpoint_17;
    wire n16594;
    wire rand_setpoint_18;
    wire n16595;
    wire rand_data_19;
    wire rand_setpoint_19;
    wire n16596;
    wire rand_data_20;
    wire rand_setpoint_20;
    wire n16597;
    wire rand_data_21;
    wire rand_setpoint_21;
    wire n16598;
    wire rand_data_22;
    wire rand_setpoint_22;
    wire n16599;
    wire rand_data_23;
    wire rand_setpoint_23;
    wire n16600;
    wire n16601;
    wire rand_data_24;
    wire bfn_14_12_0_;
    wire rand_data_25;
    wire rand_setpoint_25;
    wire n16602;
    wire rand_data_26;
    wire n16603;
    wire n16604;
    wire rand_setpoint_28;
    wire n16605;
    wire rand_data_29;
    wire rand_setpoint_29;
    wire n16606;
    wire rand_data_30;
    wire n16607;
    wire rand_data_31;
    wire n16608;
    wire rand_setpoint_13;
    wire \c0.n18234 ;
    wire rand_setpoint_1;
    wire \c0.data_out_8_1 ;
    wire \c0.data_out_7_5 ;
    wire \c0.data_out_7_7 ;
    wire \c0.n10533 ;
    wire rand_setpoint_26;
    wire \c0.data_out_5_2 ;
    wire rand_setpoint_30;
    wire rand_setpoint_27;
    wire \c0.data_out_5_3 ;
    wire \c0.n17718 ;
    wire \c0.n17829 ;
    wire \c0.data_out_10_4 ;
    wire n2837;
    wire data_out_3_0;
    wire \c0.n2_adj_2221 ;
    wire data_out_2_0;
    wire \c0.n5_adj_2433 ;
    wire data_out_frame2_14_7;
    wire \c0.n17899 ;
    wire \c0.n17899_cascade_ ;
    wire \c0.n34 ;
    wire \c0.n17736 ;
    wire \c0.n17736_cascade_ ;
    wire \c0.n18813 ;
    wire \c0.n18816 ;
    wire data_out_frame2_9_6;
    wire \c0.n10725 ;
    wire data_out_frame2_7_0;
    wire \c0.n10700 ;
    wire \c0.n16_adj_2412 ;
    wire \c0.n17_adj_2413_cascade_ ;
    wire \c0.data_out_frame2_0_1 ;
    wire \c0.n10782 ;
    wire data_out_frame2_14_1;
    wire \c0.n17862 ;
    wire \c0.n17862_cascade_ ;
    wire \c0.n17841 ;
    wire \c0.n12_adj_2410_cascade_ ;
    wire data_out_frame2_16_7;
    wire data_out_frame2_15_7;
    wire \c0.n17889 ;
    wire rand_data_18;
    wire data_out_frame2_6_2;
    wire \c0.n18645 ;
    wire \c0.n18_adj_2441 ;
    wire data_out_frame2_8_3;
    wire data_out_frame2_10_1;
    wire \c0.n17838 ;
    wire \c0.n17792 ;
    wire \c0.n33 ;
    wire data_out_frame2_6_6;
    wire data_out_frame2_10_3;
    wire \c0.n18663 ;
    wire data_out_frame2_5_0;
    wire \c0.n10911 ;
    wire data_out_frame2_11_6;
    wire rand_data_6;
    wire data_out_frame2_9_4;
    wire data_out_frame2_7_7;
    wire data_out_frame2_9_7;
    wire \c0.n10617 ;
    wire \c0.n14_adj_2362 ;
    wire data_out_frame2_12_2;
    wire data_out_frame2_10_4;
    wire \c0.n17880 ;
    wire \c0.n17789 ;
    wire data_out_frame2_5_6;
    wire \c0.n5_adj_2439 ;
    wire \c0.data_out_frame2_0_6 ;
    wire data_out_frame2_15_6;
    wire data_out_frame2_13_1;
    wire data_out_frame2_8_7;
    wire \c0.data_out_frame2_0_0 ;
    wire \c0.n10_adj_2431 ;
    wire data_out_frame2_5_2;
    wire \c0.n17865 ;
    wire rand_data_28;
    wire rand_data_11;
    wire data_out_frame2_13_7;
    wire \c0.n10_adj_2411 ;
    wire \c0.n18705 ;
    wire data_out_frame2_13_6;
    wire rand_data_27;
    wire rand_data_7;
    wire data_out_frame2_13_3;
    wire \c0.n18657 ;
    wire data_out_frame2_18_3;
    wire \c0.data_out_frame2_19_3 ;
    wire data_out_frame2_17_3;
    wire \c0.n18651_cascade_ ;
    wire data_out_frame2_16_3;
    wire \c0.data_out_frame2_20_3 ;
    wire \c0.n18654_cascade_ ;
    wire \c0.n18666 ;
    wire \c0.n18660 ;
    wire \c0.n18371 ;
    wire \c0.n18735_cascade_ ;
    wire \c0.n6_adj_2360 ;
    wire \c0.n22_adj_2259 ;
    wire \c0.n18738_cascade_ ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire data_out_frame2_18_6;
    wire \c0.n18708 ;
    wire \c0.n18762 ;
    wire \c0.n18308 ;
    wire \c0.n18777_cascade_ ;
    wire \c0.n6_adj_2218 ;
    wire \c0.n18699 ;
    wire data_out_frame2_17_6;
    wire data_out_frame2_16_6;
    wire \c0.n18702_cascade_ ;
    wire \c0.n18780 ;
    wire \c0.n22_adj_2240_cascade_ ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire \c0.n18783_cascade_ ;
    wire data_out_frame2_13_4;
    wire \c0.data_out_7__2__N_447 ;
    wire \c0.n18311 ;
    wire rand_setpoint_11;
    wire byte_transmit_counter_0;
    wire \c0.data_out_6_3 ;
    wire \c0.n5_adj_2217 ;
    wire \c0.n18201 ;
    wire \c0.data_out_7_3 ;
    wire rand_setpoint_24;
    wire \c0.data_out_6__1__N_537 ;
    wire rand_setpoint_31;
    wire \c0.data_out_7__3__N_441 ;
    wire \c0.n11277 ;
    wire \c0.data_out_1_1 ;
    wire n11017;
    wire \c0.n18250 ;
    wire rand_setpoint_8;
    wire \c0.data_out_7_0 ;
    wire \c0.n18648 ;
    wire \c0.n18642 ;
    wire \c0.n18221 ;
    wire \c0.n18765_cascade_ ;
    wire \c0.n6_adj_2227 ;
    wire \c0.n18768_cascade_ ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire data_out_frame2_18_2;
    wire \c0.data_out_frame2_19_2 ;
    wire data_out_frame2_17_2;
    wire \c0.n18633_cascade_ ;
    wire \c0.data_out_frame2_20_2 ;
    wire \c0.n18636_cascade_ ;
    wire \c0.n22_adj_2268 ;
    wire \c0.n17892 ;
    wire data_out_frame2_9_1;
    wire \c0.n10893 ;
    wire \c0.n20_adj_2438_cascade_ ;
    wire \c0.n17755 ;
    wire \c0.data_out_frame2_19_6 ;
    wire data_out_frame2_5_3;
    wire data_out_frame2_12_3;
    wire \c0.n10905 ;
    wire \c0.n10905_cascade_ ;
    wire \c0.n16_adj_2391 ;
    wire data_out_frame2_8_2;
    wire data_out_frame2_14_6;
    wire data_out_frame2_11_7;
    wire data_out_frame2_14_5;
    wire data_out_frame2_12_6;
    wire \c0.n10929 ;
    wire \c0.n10929_cascade_ ;
    wire \c0.n17823 ;
    wire \c0.n17853 ;
    wire \c0.n17823_cascade_ ;
    wire \c0.n17895 ;
    wire \c0.n17_adj_2401_cascade_ ;
    wire \c0.n17914 ;
    wire \c0.data_out_frame2_20_6 ;
    wire \c0.n10703 ;
    wire data_out_frame2_14_4;
    wire \c0.n10825 ;
    wire \c0.data_out_frame2_0_5 ;
    wire data_out_frame2_8_1;
    wire data_out_frame2_12_7;
    wire rand_data_5;
    wire data_out_frame2_12_5;
    wire data_out_frame2_6_3;
    wire \c0.n5_adj_2381 ;
    wire data_out_frame2_6_1;
    wire \c0.n30_adj_2434 ;
    wire data_out_frame2_7_3;
    wire \c0.data_out_frame2_0_3 ;
    wire data_out_frame2_14_3;
    wire data_out_frame2_15_4;
    wire data_out_frame2_7_4;
    wire \c0.n10710 ;
    wire \c0.n10710_cascade_ ;
    wire \c0.n18_adj_2402 ;
    wire \c0.n20_adj_2404 ;
    wire data_out_frame2_6_5;
    wire data_out_frame2_7_5;
    wire \c0.n5_adj_2386 ;
    wire data_out_frame2_13_5;
    wire data_out_frame2_10_7;
    wire \c0.n10877 ;
    wire \c0.n10593_cascade_ ;
    wire \c0.n14 ;
    wire data_out_frame2_7_6;
    wire data_out_frame2_5_7;
    wire data_out_frame2_9_5;
    wire data_out_frame2_9_3;
    wire \c0.n17810 ;
    wire data_out_frame2_11_2;
    wire data_out_frame2_11_3;
    wire data_out_frame2_11_1;
    wire \c0.n17798 ;
    wire \c0.n17751 ;
    wire \c0.n17868 ;
    wire \c0.n17798_cascade_ ;
    wire \c0.n17902 ;
    wire \c0.n18_adj_2393 ;
    wire data_out_frame2_16_5;
    wire \c0.n24_adj_2394_cascade_ ;
    wire data_out_frame2_15_5;
    wire \c0.n17920 ;
    wire \c0.n22_adj_2395 ;
    wire \c0.n26_adj_2396_cascade_ ;
    wire \c0.n17917 ;
    wire \c0.data_out_frame2_20_7 ;
    wire \c0.n10778 ;
    wire \c0.n17871 ;
    wire \c0.n14_adj_2406_cascade_ ;
    wire \c0.n10583 ;
    wire data_out_frame2_11_5;
    wire data_out_frame2_12_4;
    wire \c0.n17780 ;
    wire \c0.n15_adj_2407 ;
    wire data_out_frame2_5_4;
    wire \c0.n17856 ;
    wire data_out_frame2_16_2;
    wire data_out_frame2_9_2;
    wire \c0.n10887 ;
    wire \c0.n16_adj_2399 ;
    wire data_out_frame2_10_0;
    wire data_out_frame2_11_0;
    wire data_out_frame2_9_0;
    wire \c0.n18891_cascade_ ;
    wire data_out_frame2_8_0;
    wire data_out_frame2_14_0;
    wire data_out_frame2_15_0;
    wire \c0.byte_transmit_counter2_0 ;
    wire data_out_frame2_13_0;
    wire \c0.n18897_cascade_ ;
    wire data_out_frame2_12_0;
    wire \c0.n18060 ;
    wire \c0.n18057_cascade_ ;
    wire \c0.n18374 ;
    wire \c0.n18723_cascade_ ;
    wire \c0.n6_adj_2275 ;
    wire \c0.n22_adj_2373 ;
    wire \c0.n18726_cascade_ ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire \c0.n18160 ;
    wire \c0.n18161 ;
    wire \c0.n18067 ;
    wire \c0.n18771_cascade_ ;
    wire \c0.n18068 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.n18774_cascade_ ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.tx2.n9639 ;
    wire \c0.n18669 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire data_out_frame2_16_4;
    wire \c0.data_out_frame2_20_4 ;
    wire \c0.n7263 ;
    wire \c0.n18672_cascade_ ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n22_adj_2243 ;
    wire rand_setpoint_14;
    wire \c0.n11016 ;
    wire n2732;
    wire \c0.data_out_7_6 ;
    wire UART_TRANSMITTER_state_2;
    wire UART_TRANSMITTER_state_0;
    wire UART_TRANSMITTER_state_1;
    wire data_out_10__7__N_110;
    wire rand_setpoint_0;
    wire data_out_10__7__N_110_cascade_;
    wire data_out_8_0;
    wire data_out_frame2_8_4;
    wire \c0.n10788 ;
    wire data_out_frame2_10_6;
    wire \c0.n18_adj_2437 ;
    wire data_out_frame2_7_2;
    wire data_out_frame2_15_2;
    wire \c0.data_out_frame2_0_2 ;
    wire data_out_frame2_14_2;
    wire \c0.n6_adj_2409_cascade_ ;
    wire data_out_frame2_11_4;
    wire \c0.n17905 ;
    wire rand_data_12;
    wire n11114;
    wire data_out_frame2_17_4;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__51094),
            .DIN(N__51093),
            .DOUT(N__51092),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__51094),
            .PADOUT(N__51093),
            .PADIN(N__51092),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22809),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_1_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_1_pad_iopad (
            .OE(N__51085),
            .DIN(N__51084),
            .DOUT(N__51083),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_1_pad_preio (
            .PADOEN(N__51085),
            .PADOUT(N__51084),
            .PADIN(N__51083),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24903),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_22_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_22_pad_iopad (
            .OE(N__51076),
            .DIN(N__51075),
            .DOUT(N__51074),
            .PACKAGEPIN(PIN_22));
    defparam PIN_22_pad_preio.PIN_TYPE=6'b010101;
    defparam PIN_22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_22_pad_preio (
            .PADOEN(N__51076),
            .PADOUT(N__51075),
            .PADIN(N__51074),
            .CLOCKENABLE(N__32793),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35292),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__49893),
            .OUTPUTENABLE());
    defparam PIN_23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_23_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_23_pad_iopad (
            .OE(N__51067),
            .DIN(N__51066),
            .DOUT(N__51065),
            .PACKAGEPIN(PIN_23));
    defparam PIN_23_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_23_pad_preio (
            .PADOEN(N__51067),
            .PADOUT(N__51066),
            .PADIN(N__51065),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35742),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_24_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_24_pad_iopad (
            .OE(N__51058),
            .DIN(N__51057),
            .DOUT(N__51056),
            .PACKAGEPIN(PIN_24));
    defparam PIN_24_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_24_pad_preio (
            .PADOEN(N__51058),
            .PADOUT(N__51057),
            .PADIN(N__51056),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35778),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__51049),
            .DIN(N__51048),
            .DOUT(N__51047),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__51049),
            .PADOUT(N__51048),
            .PADIN(N__51047),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__18558),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_3_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_3_pad_iopad (
            .OE(N__51040),
            .DIN(N__51039),
            .DOUT(N__51038),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_3_pad_preio (
            .PADOEN(N__51040),
            .PADOUT(N__51039),
            .PADIN(N__51038),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22797),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__51031),
            .DIN(N__51030),
            .DOUT(N__51029),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__51031),
            .PADOUT(N__51030),
            .PADIN(N__51029),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__51022),
            .DIN(N__51021),
            .DOUT(N__51020),
            .PACKAGEPIN(PIN_4));
    defparam hall1_input_preio.PIN_TYPE=6'b000001;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__51022),
            .PADOUT(N__51021),
            .PADIN(N__51020),
            .CLOCKENABLE(),
            .DIN0(hall1),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__51013),
            .DIN(N__51012),
            .DOUT(N__51011),
            .PACKAGEPIN(PIN_5));
    defparam hall2_input_preio.PIN_TYPE=6'b000001;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__51013),
            .PADOUT(N__51012),
            .PADIN(N__51011),
            .CLOCKENABLE(),
            .DIN0(hall2),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__51004),
            .DIN(N__51003),
            .DOUT(N__51002),
            .PACKAGEPIN(PIN_6));
    defparam hall3_input_preio.PIN_TYPE=6'b000001;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__51004),
            .PADOUT(N__51003),
            .PADIN(N__51002),
            .CLOCKENABLE(),
            .DIN0(hall3),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__50995),
            .DIN(N__50994),
            .DOUT(N__50993),
            .PACKAGEPIN(PIN_12));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__50995),
            .PADOUT(N__50994),
            .PADIN(N__50993),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__49822),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__50986),
            .DIN(N__50985),
            .DOUT(N__50984),
            .PACKAGEPIN(PIN_11));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__50986),
            .PADOUT(N__50985),
            .PADIN(N__50984),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22769),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__22734));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__50977),
            .DIN(N__50976),
            .DOUT(N__50975),
            .PACKAGEPIN(PIN_10));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__50977),
            .PADOUT(N__50976),
            .PADIN(N__50975),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29367),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__29121));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__50968),
            .DIN(N__50967),
            .DOUT(N__50966),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__50968),
            .PADOUT(N__50967),
            .PADIN(N__50966),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__12716 (
            .O(N__50949),
            .I(N__50946));
    LocalMux I__12715 (
            .O(N__50946),
            .I(N__50942));
    CascadeMux I__12714 (
            .O(N__50945),
            .I(N__50939));
    Span4Mux_v I__12713 (
            .O(N__50942),
            .I(N__50936));
    InMux I__12712 (
            .O(N__50939),
            .I(N__50933));
    Odrv4 I__12711 (
            .O(N__50936),
            .I(rand_setpoint_0));
    LocalMux I__12710 (
            .O(N__50933),
            .I(rand_setpoint_0));
    CascadeMux I__12709 (
            .O(N__50928),
            .I(data_out_10__7__N_110_cascade_));
    InMux I__12708 (
            .O(N__50925),
            .I(N__50918));
    InMux I__12707 (
            .O(N__50924),
            .I(N__50918));
    CascadeMux I__12706 (
            .O(N__50923),
            .I(N__50915));
    LocalMux I__12705 (
            .O(N__50918),
            .I(N__50911));
    InMux I__12704 (
            .O(N__50915),
            .I(N__50905));
    InMux I__12703 (
            .O(N__50914),
            .I(N__50905));
    Span4Mux_h I__12702 (
            .O(N__50911),
            .I(N__50902));
    InMux I__12701 (
            .O(N__50910),
            .I(N__50899));
    LocalMux I__12700 (
            .O(N__50905),
            .I(N__50896));
    Span4Mux_h I__12699 (
            .O(N__50902),
            .I(N__50893));
    LocalMux I__12698 (
            .O(N__50899),
            .I(data_out_8_0));
    Odrv12 I__12697 (
            .O(N__50896),
            .I(data_out_8_0));
    Odrv4 I__12696 (
            .O(N__50893),
            .I(data_out_8_0));
    InMux I__12695 (
            .O(N__50886),
            .I(N__50882));
    InMux I__12694 (
            .O(N__50885),
            .I(N__50878));
    LocalMux I__12693 (
            .O(N__50882),
            .I(N__50875));
    InMux I__12692 (
            .O(N__50881),
            .I(N__50872));
    LocalMux I__12691 (
            .O(N__50878),
            .I(N__50865));
    Span4Mux_v I__12690 (
            .O(N__50875),
            .I(N__50860));
    LocalMux I__12689 (
            .O(N__50872),
            .I(N__50860));
    InMux I__12688 (
            .O(N__50871),
            .I(N__50857));
    InMux I__12687 (
            .O(N__50870),
            .I(N__50854));
    InMux I__12686 (
            .O(N__50869),
            .I(N__50851));
    InMux I__12685 (
            .O(N__50868),
            .I(N__50848));
    Span4Mux_v I__12684 (
            .O(N__50865),
            .I(N__50839));
    Span4Mux_h I__12683 (
            .O(N__50860),
            .I(N__50839));
    LocalMux I__12682 (
            .O(N__50857),
            .I(N__50839));
    LocalMux I__12681 (
            .O(N__50854),
            .I(N__50839));
    LocalMux I__12680 (
            .O(N__50851),
            .I(data_out_frame2_8_4));
    LocalMux I__12679 (
            .O(N__50848),
            .I(data_out_frame2_8_4));
    Odrv4 I__12678 (
            .O(N__50839),
            .I(data_out_frame2_8_4));
    CascadeMux I__12677 (
            .O(N__50832),
            .I(N__50829));
    InMux I__12676 (
            .O(N__50829),
            .I(N__50826));
    LocalMux I__12675 (
            .O(N__50826),
            .I(\c0.n10788 ));
    InMux I__12674 (
            .O(N__50823),
            .I(N__50816));
    InMux I__12673 (
            .O(N__50822),
            .I(N__50813));
    InMux I__12672 (
            .O(N__50821),
            .I(N__50810));
    InMux I__12671 (
            .O(N__50820),
            .I(N__50807));
    InMux I__12670 (
            .O(N__50819),
            .I(N__50804));
    LocalMux I__12669 (
            .O(N__50816),
            .I(N__50801));
    LocalMux I__12668 (
            .O(N__50813),
            .I(N__50798));
    LocalMux I__12667 (
            .O(N__50810),
            .I(N__50793));
    LocalMux I__12666 (
            .O(N__50807),
            .I(N__50793));
    LocalMux I__12665 (
            .O(N__50804),
            .I(N__50790));
    Span4Mux_s0_v I__12664 (
            .O(N__50801),
            .I(N__50786));
    Span4Mux_h I__12663 (
            .O(N__50798),
            .I(N__50779));
    Span4Mux_v I__12662 (
            .O(N__50793),
            .I(N__50779));
    Span4Mux_s1_v I__12661 (
            .O(N__50790),
            .I(N__50779));
    InMux I__12660 (
            .O(N__50789),
            .I(N__50776));
    Span4Mux_v I__12659 (
            .O(N__50786),
            .I(N__50773));
    Span4Mux_h I__12658 (
            .O(N__50779),
            .I(N__50770));
    LocalMux I__12657 (
            .O(N__50776),
            .I(data_out_frame2_10_6));
    Odrv4 I__12656 (
            .O(N__50773),
            .I(data_out_frame2_10_6));
    Odrv4 I__12655 (
            .O(N__50770),
            .I(data_out_frame2_10_6));
    InMux I__12654 (
            .O(N__50763),
            .I(N__50760));
    LocalMux I__12653 (
            .O(N__50760),
            .I(\c0.n18_adj_2437 ));
    InMux I__12652 (
            .O(N__50757),
            .I(N__50753));
    InMux I__12651 (
            .O(N__50756),
            .I(N__50750));
    LocalMux I__12650 (
            .O(N__50753),
            .I(N__50747));
    LocalMux I__12649 (
            .O(N__50750),
            .I(N__50744));
    Span4Mux_s2_v I__12648 (
            .O(N__50747),
            .I(N__50739));
    Span4Mux_h I__12647 (
            .O(N__50744),
            .I(N__50736));
    CascadeMux I__12646 (
            .O(N__50743),
            .I(N__50733));
    InMux I__12645 (
            .O(N__50742),
            .I(N__50730));
    Span4Mux_h I__12644 (
            .O(N__50739),
            .I(N__50727));
    Span4Mux_h I__12643 (
            .O(N__50736),
            .I(N__50724));
    InMux I__12642 (
            .O(N__50733),
            .I(N__50721));
    LocalMux I__12641 (
            .O(N__50730),
            .I(data_out_frame2_7_2));
    Odrv4 I__12640 (
            .O(N__50727),
            .I(data_out_frame2_7_2));
    Odrv4 I__12639 (
            .O(N__50724),
            .I(data_out_frame2_7_2));
    LocalMux I__12638 (
            .O(N__50721),
            .I(data_out_frame2_7_2));
    InMux I__12637 (
            .O(N__50712),
            .I(N__50707));
    InMux I__12636 (
            .O(N__50711),
            .I(N__50704));
    InMux I__12635 (
            .O(N__50710),
            .I(N__50699));
    LocalMux I__12634 (
            .O(N__50707),
            .I(N__50696));
    LocalMux I__12633 (
            .O(N__50704),
            .I(N__50693));
    InMux I__12632 (
            .O(N__50703),
            .I(N__50690));
    InMux I__12631 (
            .O(N__50702),
            .I(N__50687));
    LocalMux I__12630 (
            .O(N__50699),
            .I(data_out_frame2_15_2));
    Odrv12 I__12629 (
            .O(N__50696),
            .I(data_out_frame2_15_2));
    Odrv4 I__12628 (
            .O(N__50693),
            .I(data_out_frame2_15_2));
    LocalMux I__12627 (
            .O(N__50690),
            .I(data_out_frame2_15_2));
    LocalMux I__12626 (
            .O(N__50687),
            .I(data_out_frame2_15_2));
    InMux I__12625 (
            .O(N__50676),
            .I(N__50673));
    LocalMux I__12624 (
            .O(N__50673),
            .I(N__50668));
    InMux I__12623 (
            .O(N__50672),
            .I(N__50665));
    InMux I__12622 (
            .O(N__50671),
            .I(N__50661));
    Span4Mux_h I__12621 (
            .O(N__50668),
            .I(N__50656));
    LocalMux I__12620 (
            .O(N__50665),
            .I(N__50656));
    CascadeMux I__12619 (
            .O(N__50664),
            .I(N__50652));
    LocalMux I__12618 (
            .O(N__50661),
            .I(N__50649));
    Span4Mux_s3_v I__12617 (
            .O(N__50656),
            .I(N__50646));
    InMux I__12616 (
            .O(N__50655),
            .I(N__50643));
    InMux I__12615 (
            .O(N__50652),
            .I(N__50640));
    Span4Mux_h I__12614 (
            .O(N__50649),
            .I(N__50637));
    Span4Mux_h I__12613 (
            .O(N__50646),
            .I(N__50634));
    LocalMux I__12612 (
            .O(N__50643),
            .I(\c0.data_out_frame2_0_2 ));
    LocalMux I__12611 (
            .O(N__50640),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv4 I__12610 (
            .O(N__50637),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv4 I__12609 (
            .O(N__50634),
            .I(\c0.data_out_frame2_0_2 ));
    InMux I__12608 (
            .O(N__50625),
            .I(N__50622));
    LocalMux I__12607 (
            .O(N__50622),
            .I(N__50617));
    CascadeMux I__12606 (
            .O(N__50621),
            .I(N__50614));
    InMux I__12605 (
            .O(N__50620),
            .I(N__50610));
    Span4Mux_h I__12604 (
            .O(N__50617),
            .I(N__50607));
    InMux I__12603 (
            .O(N__50614),
            .I(N__50604));
    InMux I__12602 (
            .O(N__50613),
            .I(N__50601));
    LocalMux I__12601 (
            .O(N__50610),
            .I(N__50594));
    Span4Mux_h I__12600 (
            .O(N__50607),
            .I(N__50594));
    LocalMux I__12599 (
            .O(N__50604),
            .I(N__50594));
    LocalMux I__12598 (
            .O(N__50601),
            .I(data_out_frame2_14_2));
    Odrv4 I__12597 (
            .O(N__50594),
            .I(data_out_frame2_14_2));
    CascadeMux I__12596 (
            .O(N__50589),
            .I(\c0.n6_adj_2409_cascade_ ));
    InMux I__12595 (
            .O(N__50586),
            .I(N__50582));
    InMux I__12594 (
            .O(N__50585),
            .I(N__50578));
    LocalMux I__12593 (
            .O(N__50582),
            .I(N__50575));
    CascadeMux I__12592 (
            .O(N__50581),
            .I(N__50572));
    LocalMux I__12591 (
            .O(N__50578),
            .I(N__50568));
    Span4Mux_h I__12590 (
            .O(N__50575),
            .I(N__50565));
    InMux I__12589 (
            .O(N__50572),
            .I(N__50560));
    InMux I__12588 (
            .O(N__50571),
            .I(N__50560));
    Odrv4 I__12587 (
            .O(N__50568),
            .I(data_out_frame2_11_4));
    Odrv4 I__12586 (
            .O(N__50565),
            .I(data_out_frame2_11_4));
    LocalMux I__12585 (
            .O(N__50560),
            .I(data_out_frame2_11_4));
    InMux I__12584 (
            .O(N__50553),
            .I(N__50549));
    CascadeMux I__12583 (
            .O(N__50552),
            .I(N__50546));
    LocalMux I__12582 (
            .O(N__50549),
            .I(N__50543));
    InMux I__12581 (
            .O(N__50546),
            .I(N__50540));
    Span4Mux_s3_v I__12580 (
            .O(N__50543),
            .I(N__50537));
    LocalMux I__12579 (
            .O(N__50540),
            .I(N__50534));
    Odrv4 I__12578 (
            .O(N__50537),
            .I(\c0.n17905 ));
    Odrv4 I__12577 (
            .O(N__50534),
            .I(\c0.n17905 ));
    InMux I__12576 (
            .O(N__50529),
            .I(N__50526));
    LocalMux I__12575 (
            .O(N__50526),
            .I(N__50520));
    InMux I__12574 (
            .O(N__50525),
            .I(N__50517));
    InMux I__12573 (
            .O(N__50524),
            .I(N__50514));
    InMux I__12572 (
            .O(N__50523),
            .I(N__50511));
    Span4Mux_h I__12571 (
            .O(N__50520),
            .I(N__50506));
    LocalMux I__12570 (
            .O(N__50517),
            .I(N__50506));
    LocalMux I__12569 (
            .O(N__50514),
            .I(N__50501));
    LocalMux I__12568 (
            .O(N__50511),
            .I(N__50498));
    Span4Mux_h I__12567 (
            .O(N__50506),
            .I(N__50495));
    InMux I__12566 (
            .O(N__50505),
            .I(N__50492));
    InMux I__12565 (
            .O(N__50504),
            .I(N__50489));
    Span4Mux_v I__12564 (
            .O(N__50501),
            .I(N__50484));
    Span4Mux_v I__12563 (
            .O(N__50498),
            .I(N__50484));
    Odrv4 I__12562 (
            .O(N__50495),
            .I(rand_data_12));
    LocalMux I__12561 (
            .O(N__50492),
            .I(rand_data_12));
    LocalMux I__12560 (
            .O(N__50489),
            .I(rand_data_12));
    Odrv4 I__12559 (
            .O(N__50484),
            .I(rand_data_12));
    CEMux I__12558 (
            .O(N__50475),
            .I(N__50470));
    CEMux I__12557 (
            .O(N__50474),
            .I(N__50459));
    InMux I__12556 (
            .O(N__50473),
            .I(N__50456));
    LocalMux I__12555 (
            .O(N__50470),
            .I(N__50441));
    CEMux I__12554 (
            .O(N__50469),
            .I(N__50438));
    CEMux I__12553 (
            .O(N__50468),
            .I(N__50420));
    CEMux I__12552 (
            .O(N__50467),
            .I(N__50416));
    CEMux I__12551 (
            .O(N__50466),
            .I(N__50413));
    InMux I__12550 (
            .O(N__50465),
            .I(N__50406));
    InMux I__12549 (
            .O(N__50464),
            .I(N__50406));
    InMux I__12548 (
            .O(N__50463),
            .I(N__50406));
    CEMux I__12547 (
            .O(N__50462),
            .I(N__50395));
    LocalMux I__12546 (
            .O(N__50459),
            .I(N__50392));
    LocalMux I__12545 (
            .O(N__50456),
            .I(N__50389));
    InMux I__12544 (
            .O(N__50455),
            .I(N__50380));
    InMux I__12543 (
            .O(N__50454),
            .I(N__50380));
    InMux I__12542 (
            .O(N__50453),
            .I(N__50380));
    InMux I__12541 (
            .O(N__50452),
            .I(N__50380));
    InMux I__12540 (
            .O(N__50451),
            .I(N__50377));
    InMux I__12539 (
            .O(N__50450),
            .I(N__50374));
    InMux I__12538 (
            .O(N__50449),
            .I(N__50371));
    InMux I__12537 (
            .O(N__50448),
            .I(N__50364));
    InMux I__12536 (
            .O(N__50447),
            .I(N__50364));
    InMux I__12535 (
            .O(N__50446),
            .I(N__50364));
    InMux I__12534 (
            .O(N__50445),
            .I(N__50361));
    CEMux I__12533 (
            .O(N__50444),
            .I(N__50351));
    Span4Mux_s2_v I__12532 (
            .O(N__50441),
            .I(N__50345));
    LocalMux I__12531 (
            .O(N__50438),
            .I(N__50345));
    CEMux I__12530 (
            .O(N__50437),
            .I(N__50342));
    InMux I__12529 (
            .O(N__50436),
            .I(N__50339));
    InMux I__12528 (
            .O(N__50435),
            .I(N__50336));
    InMux I__12527 (
            .O(N__50434),
            .I(N__50327));
    InMux I__12526 (
            .O(N__50433),
            .I(N__50327));
    InMux I__12525 (
            .O(N__50432),
            .I(N__50327));
    InMux I__12524 (
            .O(N__50431),
            .I(N__50327));
    InMux I__12523 (
            .O(N__50430),
            .I(N__50324));
    InMux I__12522 (
            .O(N__50429),
            .I(N__50317));
    InMux I__12521 (
            .O(N__50428),
            .I(N__50317));
    InMux I__12520 (
            .O(N__50427),
            .I(N__50317));
    CEMux I__12519 (
            .O(N__50426),
            .I(N__50310));
    InMux I__12518 (
            .O(N__50425),
            .I(N__50303));
    InMux I__12517 (
            .O(N__50424),
            .I(N__50303));
    InMux I__12516 (
            .O(N__50423),
            .I(N__50303));
    LocalMux I__12515 (
            .O(N__50420),
            .I(N__50294));
    CEMux I__12514 (
            .O(N__50419),
            .I(N__50291));
    LocalMux I__12513 (
            .O(N__50416),
            .I(N__50288));
    LocalMux I__12512 (
            .O(N__50413),
            .I(N__50285));
    LocalMux I__12511 (
            .O(N__50406),
            .I(N__50282));
    InMux I__12510 (
            .O(N__50405),
            .I(N__50277));
    InMux I__12509 (
            .O(N__50404),
            .I(N__50277));
    InMux I__12508 (
            .O(N__50403),
            .I(N__50264));
    InMux I__12507 (
            .O(N__50402),
            .I(N__50264));
    InMux I__12506 (
            .O(N__50401),
            .I(N__50264));
    InMux I__12505 (
            .O(N__50400),
            .I(N__50264));
    InMux I__12504 (
            .O(N__50399),
            .I(N__50264));
    InMux I__12503 (
            .O(N__50398),
            .I(N__50264));
    LocalMux I__12502 (
            .O(N__50395),
            .I(N__50237));
    Span4Mux_s3_v I__12501 (
            .O(N__50392),
            .I(N__50234));
    Span4Mux_s3_v I__12500 (
            .O(N__50389),
            .I(N__50229));
    LocalMux I__12499 (
            .O(N__50380),
            .I(N__50229));
    LocalMux I__12498 (
            .O(N__50377),
            .I(N__50226));
    LocalMux I__12497 (
            .O(N__50374),
            .I(N__50219));
    LocalMux I__12496 (
            .O(N__50371),
            .I(N__50219));
    LocalMux I__12495 (
            .O(N__50364),
            .I(N__50219));
    LocalMux I__12494 (
            .O(N__50361),
            .I(N__50216));
    InMux I__12493 (
            .O(N__50360),
            .I(N__50201));
    InMux I__12492 (
            .O(N__50359),
            .I(N__50201));
    InMux I__12491 (
            .O(N__50358),
            .I(N__50201));
    InMux I__12490 (
            .O(N__50357),
            .I(N__50201));
    InMux I__12489 (
            .O(N__50356),
            .I(N__50201));
    InMux I__12488 (
            .O(N__50355),
            .I(N__50201));
    InMux I__12487 (
            .O(N__50354),
            .I(N__50201));
    LocalMux I__12486 (
            .O(N__50351),
            .I(N__50198));
    CEMux I__12485 (
            .O(N__50350),
            .I(N__50195));
    Span4Mux_v I__12484 (
            .O(N__50345),
            .I(N__50188));
    LocalMux I__12483 (
            .O(N__50342),
            .I(N__50188));
    LocalMux I__12482 (
            .O(N__50339),
            .I(N__50188));
    LocalMux I__12481 (
            .O(N__50336),
            .I(N__50179));
    LocalMux I__12480 (
            .O(N__50327),
            .I(N__50179));
    LocalMux I__12479 (
            .O(N__50324),
            .I(N__50179));
    LocalMux I__12478 (
            .O(N__50317),
            .I(N__50179));
    InMux I__12477 (
            .O(N__50316),
            .I(N__50170));
    InMux I__12476 (
            .O(N__50315),
            .I(N__50170));
    InMux I__12475 (
            .O(N__50314),
            .I(N__50170));
    InMux I__12474 (
            .O(N__50313),
            .I(N__50170));
    LocalMux I__12473 (
            .O(N__50310),
            .I(N__50165));
    LocalMux I__12472 (
            .O(N__50303),
            .I(N__50165));
    InMux I__12471 (
            .O(N__50302),
            .I(N__50152));
    InMux I__12470 (
            .O(N__50301),
            .I(N__50152));
    InMux I__12469 (
            .O(N__50300),
            .I(N__50152));
    InMux I__12468 (
            .O(N__50299),
            .I(N__50152));
    InMux I__12467 (
            .O(N__50298),
            .I(N__50152));
    InMux I__12466 (
            .O(N__50297),
            .I(N__50152));
    Span4Mux_v I__12465 (
            .O(N__50294),
            .I(N__50115));
    LocalMux I__12464 (
            .O(N__50291),
            .I(N__50112));
    Span4Mux_s3_v I__12463 (
            .O(N__50288),
            .I(N__50109));
    Span4Mux_h I__12462 (
            .O(N__50285),
            .I(N__50100));
    Span4Mux_v I__12461 (
            .O(N__50282),
            .I(N__50100));
    LocalMux I__12460 (
            .O(N__50277),
            .I(N__50100));
    LocalMux I__12459 (
            .O(N__50264),
            .I(N__50100));
    InMux I__12458 (
            .O(N__50263),
            .I(N__50091));
    InMux I__12457 (
            .O(N__50262),
            .I(N__50091));
    InMux I__12456 (
            .O(N__50261),
            .I(N__50091));
    InMux I__12455 (
            .O(N__50260),
            .I(N__50091));
    InMux I__12454 (
            .O(N__50259),
            .I(N__50076));
    InMux I__12453 (
            .O(N__50258),
            .I(N__50076));
    InMux I__12452 (
            .O(N__50257),
            .I(N__50076));
    InMux I__12451 (
            .O(N__50256),
            .I(N__50076));
    InMux I__12450 (
            .O(N__50255),
            .I(N__50076));
    InMux I__12449 (
            .O(N__50254),
            .I(N__50076));
    InMux I__12448 (
            .O(N__50253),
            .I(N__50076));
    InMux I__12447 (
            .O(N__50252),
            .I(N__50059));
    InMux I__12446 (
            .O(N__50251),
            .I(N__50059));
    InMux I__12445 (
            .O(N__50250),
            .I(N__50059));
    InMux I__12444 (
            .O(N__50249),
            .I(N__50059));
    InMux I__12443 (
            .O(N__50248),
            .I(N__50059));
    InMux I__12442 (
            .O(N__50247),
            .I(N__50059));
    InMux I__12441 (
            .O(N__50246),
            .I(N__50059));
    InMux I__12440 (
            .O(N__50245),
            .I(N__50059));
    InMux I__12439 (
            .O(N__50244),
            .I(N__50048));
    InMux I__12438 (
            .O(N__50243),
            .I(N__50048));
    InMux I__12437 (
            .O(N__50242),
            .I(N__50048));
    InMux I__12436 (
            .O(N__50241),
            .I(N__50048));
    InMux I__12435 (
            .O(N__50240),
            .I(N__50048));
    Span4Mux_s3_v I__12434 (
            .O(N__50237),
            .I(N__50033));
    Span4Mux_h I__12433 (
            .O(N__50234),
            .I(N__50033));
    Span4Mux_v I__12432 (
            .O(N__50229),
            .I(N__50033));
    Span4Mux_s3_v I__12431 (
            .O(N__50226),
            .I(N__50033));
    Span4Mux_h I__12430 (
            .O(N__50219),
            .I(N__50033));
    Span4Mux_h I__12429 (
            .O(N__50216),
            .I(N__50033));
    LocalMux I__12428 (
            .O(N__50201),
            .I(N__50033));
    Span4Mux_s2_v I__12427 (
            .O(N__50198),
            .I(N__50018));
    LocalMux I__12426 (
            .O(N__50195),
            .I(N__50018));
    Span4Mux_h I__12425 (
            .O(N__50188),
            .I(N__50018));
    Span4Mux_v I__12424 (
            .O(N__50179),
            .I(N__50018));
    LocalMux I__12423 (
            .O(N__50170),
            .I(N__50018));
    Span4Mux_s2_v I__12422 (
            .O(N__50165),
            .I(N__50018));
    LocalMux I__12421 (
            .O(N__50152),
            .I(N__50018));
    InMux I__12420 (
            .O(N__50151),
            .I(N__50001));
    InMux I__12419 (
            .O(N__50150),
            .I(N__50001));
    InMux I__12418 (
            .O(N__50149),
            .I(N__50001));
    InMux I__12417 (
            .O(N__50148),
            .I(N__50001));
    InMux I__12416 (
            .O(N__50147),
            .I(N__50001));
    InMux I__12415 (
            .O(N__50146),
            .I(N__50001));
    InMux I__12414 (
            .O(N__50145),
            .I(N__50001));
    InMux I__12413 (
            .O(N__50144),
            .I(N__50001));
    InMux I__12412 (
            .O(N__50143),
            .I(N__49988));
    InMux I__12411 (
            .O(N__50142),
            .I(N__49988));
    InMux I__12410 (
            .O(N__50141),
            .I(N__49988));
    InMux I__12409 (
            .O(N__50140),
            .I(N__49988));
    InMux I__12408 (
            .O(N__50139),
            .I(N__49988));
    InMux I__12407 (
            .O(N__50138),
            .I(N__49988));
    InMux I__12406 (
            .O(N__50137),
            .I(N__49973));
    InMux I__12405 (
            .O(N__50136),
            .I(N__49973));
    InMux I__12404 (
            .O(N__50135),
            .I(N__49973));
    InMux I__12403 (
            .O(N__50134),
            .I(N__49973));
    InMux I__12402 (
            .O(N__50133),
            .I(N__49973));
    InMux I__12401 (
            .O(N__50132),
            .I(N__49973));
    InMux I__12400 (
            .O(N__50131),
            .I(N__49973));
    InMux I__12399 (
            .O(N__50130),
            .I(N__49958));
    InMux I__12398 (
            .O(N__50129),
            .I(N__49958));
    InMux I__12397 (
            .O(N__50128),
            .I(N__49958));
    InMux I__12396 (
            .O(N__50127),
            .I(N__49958));
    InMux I__12395 (
            .O(N__50126),
            .I(N__49958));
    InMux I__12394 (
            .O(N__50125),
            .I(N__49958));
    InMux I__12393 (
            .O(N__50124),
            .I(N__49958));
    InMux I__12392 (
            .O(N__50123),
            .I(N__49945));
    InMux I__12391 (
            .O(N__50122),
            .I(N__49945));
    InMux I__12390 (
            .O(N__50121),
            .I(N__49945));
    InMux I__12389 (
            .O(N__50120),
            .I(N__49945));
    InMux I__12388 (
            .O(N__50119),
            .I(N__49945));
    InMux I__12387 (
            .O(N__50118),
            .I(N__49945));
    Odrv4 I__12386 (
            .O(N__50115),
            .I(n11114));
    Odrv4 I__12385 (
            .O(N__50112),
            .I(n11114));
    Odrv4 I__12384 (
            .O(N__50109),
            .I(n11114));
    Odrv4 I__12383 (
            .O(N__50100),
            .I(n11114));
    LocalMux I__12382 (
            .O(N__50091),
            .I(n11114));
    LocalMux I__12381 (
            .O(N__50076),
            .I(n11114));
    LocalMux I__12380 (
            .O(N__50059),
            .I(n11114));
    LocalMux I__12379 (
            .O(N__50048),
            .I(n11114));
    Odrv4 I__12378 (
            .O(N__50033),
            .I(n11114));
    Odrv4 I__12377 (
            .O(N__50018),
            .I(n11114));
    LocalMux I__12376 (
            .O(N__50001),
            .I(n11114));
    LocalMux I__12375 (
            .O(N__49988),
            .I(n11114));
    LocalMux I__12374 (
            .O(N__49973),
            .I(n11114));
    LocalMux I__12373 (
            .O(N__49958),
            .I(n11114));
    LocalMux I__12372 (
            .O(N__49945),
            .I(n11114));
    CascadeMux I__12371 (
            .O(N__49914),
            .I(N__49911));
    InMux I__12370 (
            .O(N__49911),
            .I(N__49908));
    LocalMux I__12369 (
            .O(N__49908),
            .I(N__49904));
    InMux I__12368 (
            .O(N__49907),
            .I(N__49901));
    Span4Mux_v I__12367 (
            .O(N__49904),
            .I(N__49898));
    LocalMux I__12366 (
            .O(N__49901),
            .I(data_out_frame2_17_4));
    Odrv4 I__12365 (
            .O(N__49898),
            .I(data_out_frame2_17_4));
    ClkMux I__12364 (
            .O(N__49893),
            .I(N__49206));
    ClkMux I__12363 (
            .O(N__49892),
            .I(N__49206));
    ClkMux I__12362 (
            .O(N__49891),
            .I(N__49206));
    ClkMux I__12361 (
            .O(N__49890),
            .I(N__49206));
    ClkMux I__12360 (
            .O(N__49889),
            .I(N__49206));
    ClkMux I__12359 (
            .O(N__49888),
            .I(N__49206));
    ClkMux I__12358 (
            .O(N__49887),
            .I(N__49206));
    ClkMux I__12357 (
            .O(N__49886),
            .I(N__49206));
    ClkMux I__12356 (
            .O(N__49885),
            .I(N__49206));
    ClkMux I__12355 (
            .O(N__49884),
            .I(N__49206));
    ClkMux I__12354 (
            .O(N__49883),
            .I(N__49206));
    ClkMux I__12353 (
            .O(N__49882),
            .I(N__49206));
    ClkMux I__12352 (
            .O(N__49881),
            .I(N__49206));
    ClkMux I__12351 (
            .O(N__49880),
            .I(N__49206));
    ClkMux I__12350 (
            .O(N__49879),
            .I(N__49206));
    ClkMux I__12349 (
            .O(N__49878),
            .I(N__49206));
    ClkMux I__12348 (
            .O(N__49877),
            .I(N__49206));
    ClkMux I__12347 (
            .O(N__49876),
            .I(N__49206));
    ClkMux I__12346 (
            .O(N__49875),
            .I(N__49206));
    ClkMux I__12345 (
            .O(N__49874),
            .I(N__49206));
    ClkMux I__12344 (
            .O(N__49873),
            .I(N__49206));
    ClkMux I__12343 (
            .O(N__49872),
            .I(N__49206));
    ClkMux I__12342 (
            .O(N__49871),
            .I(N__49206));
    ClkMux I__12341 (
            .O(N__49870),
            .I(N__49206));
    ClkMux I__12340 (
            .O(N__49869),
            .I(N__49206));
    ClkMux I__12339 (
            .O(N__49868),
            .I(N__49206));
    ClkMux I__12338 (
            .O(N__49867),
            .I(N__49206));
    ClkMux I__12337 (
            .O(N__49866),
            .I(N__49206));
    ClkMux I__12336 (
            .O(N__49865),
            .I(N__49206));
    ClkMux I__12335 (
            .O(N__49864),
            .I(N__49206));
    ClkMux I__12334 (
            .O(N__49863),
            .I(N__49206));
    ClkMux I__12333 (
            .O(N__49862),
            .I(N__49206));
    ClkMux I__12332 (
            .O(N__49861),
            .I(N__49206));
    ClkMux I__12331 (
            .O(N__49860),
            .I(N__49206));
    ClkMux I__12330 (
            .O(N__49859),
            .I(N__49206));
    ClkMux I__12329 (
            .O(N__49858),
            .I(N__49206));
    ClkMux I__12328 (
            .O(N__49857),
            .I(N__49206));
    ClkMux I__12327 (
            .O(N__49856),
            .I(N__49206));
    ClkMux I__12326 (
            .O(N__49855),
            .I(N__49206));
    ClkMux I__12325 (
            .O(N__49854),
            .I(N__49206));
    ClkMux I__12324 (
            .O(N__49853),
            .I(N__49206));
    ClkMux I__12323 (
            .O(N__49852),
            .I(N__49206));
    ClkMux I__12322 (
            .O(N__49851),
            .I(N__49206));
    ClkMux I__12321 (
            .O(N__49850),
            .I(N__49206));
    ClkMux I__12320 (
            .O(N__49849),
            .I(N__49206));
    ClkMux I__12319 (
            .O(N__49848),
            .I(N__49206));
    ClkMux I__12318 (
            .O(N__49847),
            .I(N__49206));
    ClkMux I__12317 (
            .O(N__49846),
            .I(N__49206));
    ClkMux I__12316 (
            .O(N__49845),
            .I(N__49206));
    ClkMux I__12315 (
            .O(N__49844),
            .I(N__49206));
    ClkMux I__12314 (
            .O(N__49843),
            .I(N__49206));
    ClkMux I__12313 (
            .O(N__49842),
            .I(N__49206));
    ClkMux I__12312 (
            .O(N__49841),
            .I(N__49206));
    ClkMux I__12311 (
            .O(N__49840),
            .I(N__49206));
    ClkMux I__12310 (
            .O(N__49839),
            .I(N__49206));
    ClkMux I__12309 (
            .O(N__49838),
            .I(N__49206));
    ClkMux I__12308 (
            .O(N__49837),
            .I(N__49206));
    ClkMux I__12307 (
            .O(N__49836),
            .I(N__49206));
    ClkMux I__12306 (
            .O(N__49835),
            .I(N__49206));
    ClkMux I__12305 (
            .O(N__49834),
            .I(N__49206));
    ClkMux I__12304 (
            .O(N__49833),
            .I(N__49206));
    ClkMux I__12303 (
            .O(N__49832),
            .I(N__49206));
    ClkMux I__12302 (
            .O(N__49831),
            .I(N__49206));
    ClkMux I__12301 (
            .O(N__49830),
            .I(N__49206));
    ClkMux I__12300 (
            .O(N__49829),
            .I(N__49206));
    ClkMux I__12299 (
            .O(N__49828),
            .I(N__49206));
    ClkMux I__12298 (
            .O(N__49827),
            .I(N__49206));
    ClkMux I__12297 (
            .O(N__49826),
            .I(N__49206));
    ClkMux I__12296 (
            .O(N__49825),
            .I(N__49206));
    ClkMux I__12295 (
            .O(N__49824),
            .I(N__49206));
    ClkMux I__12294 (
            .O(N__49823),
            .I(N__49206));
    ClkMux I__12293 (
            .O(N__49822),
            .I(N__49206));
    ClkMux I__12292 (
            .O(N__49821),
            .I(N__49206));
    ClkMux I__12291 (
            .O(N__49820),
            .I(N__49206));
    ClkMux I__12290 (
            .O(N__49819),
            .I(N__49206));
    ClkMux I__12289 (
            .O(N__49818),
            .I(N__49206));
    ClkMux I__12288 (
            .O(N__49817),
            .I(N__49206));
    ClkMux I__12287 (
            .O(N__49816),
            .I(N__49206));
    ClkMux I__12286 (
            .O(N__49815),
            .I(N__49206));
    ClkMux I__12285 (
            .O(N__49814),
            .I(N__49206));
    ClkMux I__12284 (
            .O(N__49813),
            .I(N__49206));
    ClkMux I__12283 (
            .O(N__49812),
            .I(N__49206));
    ClkMux I__12282 (
            .O(N__49811),
            .I(N__49206));
    ClkMux I__12281 (
            .O(N__49810),
            .I(N__49206));
    ClkMux I__12280 (
            .O(N__49809),
            .I(N__49206));
    ClkMux I__12279 (
            .O(N__49808),
            .I(N__49206));
    ClkMux I__12278 (
            .O(N__49807),
            .I(N__49206));
    ClkMux I__12277 (
            .O(N__49806),
            .I(N__49206));
    ClkMux I__12276 (
            .O(N__49805),
            .I(N__49206));
    ClkMux I__12275 (
            .O(N__49804),
            .I(N__49206));
    ClkMux I__12274 (
            .O(N__49803),
            .I(N__49206));
    ClkMux I__12273 (
            .O(N__49802),
            .I(N__49206));
    ClkMux I__12272 (
            .O(N__49801),
            .I(N__49206));
    ClkMux I__12271 (
            .O(N__49800),
            .I(N__49206));
    ClkMux I__12270 (
            .O(N__49799),
            .I(N__49206));
    ClkMux I__12269 (
            .O(N__49798),
            .I(N__49206));
    ClkMux I__12268 (
            .O(N__49797),
            .I(N__49206));
    ClkMux I__12267 (
            .O(N__49796),
            .I(N__49206));
    ClkMux I__12266 (
            .O(N__49795),
            .I(N__49206));
    ClkMux I__12265 (
            .O(N__49794),
            .I(N__49206));
    ClkMux I__12264 (
            .O(N__49793),
            .I(N__49206));
    ClkMux I__12263 (
            .O(N__49792),
            .I(N__49206));
    ClkMux I__12262 (
            .O(N__49791),
            .I(N__49206));
    ClkMux I__12261 (
            .O(N__49790),
            .I(N__49206));
    ClkMux I__12260 (
            .O(N__49789),
            .I(N__49206));
    ClkMux I__12259 (
            .O(N__49788),
            .I(N__49206));
    ClkMux I__12258 (
            .O(N__49787),
            .I(N__49206));
    ClkMux I__12257 (
            .O(N__49786),
            .I(N__49206));
    ClkMux I__12256 (
            .O(N__49785),
            .I(N__49206));
    ClkMux I__12255 (
            .O(N__49784),
            .I(N__49206));
    ClkMux I__12254 (
            .O(N__49783),
            .I(N__49206));
    ClkMux I__12253 (
            .O(N__49782),
            .I(N__49206));
    ClkMux I__12252 (
            .O(N__49781),
            .I(N__49206));
    ClkMux I__12251 (
            .O(N__49780),
            .I(N__49206));
    ClkMux I__12250 (
            .O(N__49779),
            .I(N__49206));
    ClkMux I__12249 (
            .O(N__49778),
            .I(N__49206));
    ClkMux I__12248 (
            .O(N__49777),
            .I(N__49206));
    ClkMux I__12247 (
            .O(N__49776),
            .I(N__49206));
    ClkMux I__12246 (
            .O(N__49775),
            .I(N__49206));
    ClkMux I__12245 (
            .O(N__49774),
            .I(N__49206));
    ClkMux I__12244 (
            .O(N__49773),
            .I(N__49206));
    ClkMux I__12243 (
            .O(N__49772),
            .I(N__49206));
    ClkMux I__12242 (
            .O(N__49771),
            .I(N__49206));
    ClkMux I__12241 (
            .O(N__49770),
            .I(N__49206));
    ClkMux I__12240 (
            .O(N__49769),
            .I(N__49206));
    ClkMux I__12239 (
            .O(N__49768),
            .I(N__49206));
    ClkMux I__12238 (
            .O(N__49767),
            .I(N__49206));
    ClkMux I__12237 (
            .O(N__49766),
            .I(N__49206));
    ClkMux I__12236 (
            .O(N__49765),
            .I(N__49206));
    ClkMux I__12235 (
            .O(N__49764),
            .I(N__49206));
    ClkMux I__12234 (
            .O(N__49763),
            .I(N__49206));
    ClkMux I__12233 (
            .O(N__49762),
            .I(N__49206));
    ClkMux I__12232 (
            .O(N__49761),
            .I(N__49206));
    ClkMux I__12231 (
            .O(N__49760),
            .I(N__49206));
    ClkMux I__12230 (
            .O(N__49759),
            .I(N__49206));
    ClkMux I__12229 (
            .O(N__49758),
            .I(N__49206));
    ClkMux I__12228 (
            .O(N__49757),
            .I(N__49206));
    ClkMux I__12227 (
            .O(N__49756),
            .I(N__49206));
    ClkMux I__12226 (
            .O(N__49755),
            .I(N__49206));
    ClkMux I__12225 (
            .O(N__49754),
            .I(N__49206));
    ClkMux I__12224 (
            .O(N__49753),
            .I(N__49206));
    ClkMux I__12223 (
            .O(N__49752),
            .I(N__49206));
    ClkMux I__12222 (
            .O(N__49751),
            .I(N__49206));
    ClkMux I__12221 (
            .O(N__49750),
            .I(N__49206));
    ClkMux I__12220 (
            .O(N__49749),
            .I(N__49206));
    ClkMux I__12219 (
            .O(N__49748),
            .I(N__49206));
    ClkMux I__12218 (
            .O(N__49747),
            .I(N__49206));
    ClkMux I__12217 (
            .O(N__49746),
            .I(N__49206));
    ClkMux I__12216 (
            .O(N__49745),
            .I(N__49206));
    ClkMux I__12215 (
            .O(N__49744),
            .I(N__49206));
    ClkMux I__12214 (
            .O(N__49743),
            .I(N__49206));
    ClkMux I__12213 (
            .O(N__49742),
            .I(N__49206));
    ClkMux I__12212 (
            .O(N__49741),
            .I(N__49206));
    ClkMux I__12211 (
            .O(N__49740),
            .I(N__49206));
    ClkMux I__12210 (
            .O(N__49739),
            .I(N__49206));
    ClkMux I__12209 (
            .O(N__49738),
            .I(N__49206));
    ClkMux I__12208 (
            .O(N__49737),
            .I(N__49206));
    ClkMux I__12207 (
            .O(N__49736),
            .I(N__49206));
    ClkMux I__12206 (
            .O(N__49735),
            .I(N__49206));
    ClkMux I__12205 (
            .O(N__49734),
            .I(N__49206));
    ClkMux I__12204 (
            .O(N__49733),
            .I(N__49206));
    ClkMux I__12203 (
            .O(N__49732),
            .I(N__49206));
    ClkMux I__12202 (
            .O(N__49731),
            .I(N__49206));
    ClkMux I__12201 (
            .O(N__49730),
            .I(N__49206));
    ClkMux I__12200 (
            .O(N__49729),
            .I(N__49206));
    ClkMux I__12199 (
            .O(N__49728),
            .I(N__49206));
    ClkMux I__12198 (
            .O(N__49727),
            .I(N__49206));
    ClkMux I__12197 (
            .O(N__49726),
            .I(N__49206));
    ClkMux I__12196 (
            .O(N__49725),
            .I(N__49206));
    ClkMux I__12195 (
            .O(N__49724),
            .I(N__49206));
    ClkMux I__12194 (
            .O(N__49723),
            .I(N__49206));
    ClkMux I__12193 (
            .O(N__49722),
            .I(N__49206));
    ClkMux I__12192 (
            .O(N__49721),
            .I(N__49206));
    ClkMux I__12191 (
            .O(N__49720),
            .I(N__49206));
    ClkMux I__12190 (
            .O(N__49719),
            .I(N__49206));
    ClkMux I__12189 (
            .O(N__49718),
            .I(N__49206));
    ClkMux I__12188 (
            .O(N__49717),
            .I(N__49206));
    ClkMux I__12187 (
            .O(N__49716),
            .I(N__49206));
    ClkMux I__12186 (
            .O(N__49715),
            .I(N__49206));
    ClkMux I__12185 (
            .O(N__49714),
            .I(N__49206));
    ClkMux I__12184 (
            .O(N__49713),
            .I(N__49206));
    ClkMux I__12183 (
            .O(N__49712),
            .I(N__49206));
    ClkMux I__12182 (
            .O(N__49711),
            .I(N__49206));
    ClkMux I__12181 (
            .O(N__49710),
            .I(N__49206));
    ClkMux I__12180 (
            .O(N__49709),
            .I(N__49206));
    ClkMux I__12179 (
            .O(N__49708),
            .I(N__49206));
    ClkMux I__12178 (
            .O(N__49707),
            .I(N__49206));
    ClkMux I__12177 (
            .O(N__49706),
            .I(N__49206));
    ClkMux I__12176 (
            .O(N__49705),
            .I(N__49206));
    ClkMux I__12175 (
            .O(N__49704),
            .I(N__49206));
    ClkMux I__12174 (
            .O(N__49703),
            .I(N__49206));
    ClkMux I__12173 (
            .O(N__49702),
            .I(N__49206));
    ClkMux I__12172 (
            .O(N__49701),
            .I(N__49206));
    ClkMux I__12171 (
            .O(N__49700),
            .I(N__49206));
    ClkMux I__12170 (
            .O(N__49699),
            .I(N__49206));
    ClkMux I__12169 (
            .O(N__49698),
            .I(N__49206));
    ClkMux I__12168 (
            .O(N__49697),
            .I(N__49206));
    ClkMux I__12167 (
            .O(N__49696),
            .I(N__49206));
    ClkMux I__12166 (
            .O(N__49695),
            .I(N__49206));
    ClkMux I__12165 (
            .O(N__49694),
            .I(N__49206));
    ClkMux I__12164 (
            .O(N__49693),
            .I(N__49206));
    ClkMux I__12163 (
            .O(N__49692),
            .I(N__49206));
    ClkMux I__12162 (
            .O(N__49691),
            .I(N__49206));
    ClkMux I__12161 (
            .O(N__49690),
            .I(N__49206));
    ClkMux I__12160 (
            .O(N__49689),
            .I(N__49206));
    ClkMux I__12159 (
            .O(N__49688),
            .I(N__49206));
    ClkMux I__12158 (
            .O(N__49687),
            .I(N__49206));
    ClkMux I__12157 (
            .O(N__49686),
            .I(N__49206));
    ClkMux I__12156 (
            .O(N__49685),
            .I(N__49206));
    ClkMux I__12155 (
            .O(N__49684),
            .I(N__49206));
    ClkMux I__12154 (
            .O(N__49683),
            .I(N__49206));
    ClkMux I__12153 (
            .O(N__49682),
            .I(N__49206));
    ClkMux I__12152 (
            .O(N__49681),
            .I(N__49206));
    ClkMux I__12151 (
            .O(N__49680),
            .I(N__49206));
    ClkMux I__12150 (
            .O(N__49679),
            .I(N__49206));
    ClkMux I__12149 (
            .O(N__49678),
            .I(N__49206));
    ClkMux I__12148 (
            .O(N__49677),
            .I(N__49206));
    ClkMux I__12147 (
            .O(N__49676),
            .I(N__49206));
    ClkMux I__12146 (
            .O(N__49675),
            .I(N__49206));
    ClkMux I__12145 (
            .O(N__49674),
            .I(N__49206));
    ClkMux I__12144 (
            .O(N__49673),
            .I(N__49206));
    ClkMux I__12143 (
            .O(N__49672),
            .I(N__49206));
    ClkMux I__12142 (
            .O(N__49671),
            .I(N__49206));
    ClkMux I__12141 (
            .O(N__49670),
            .I(N__49206));
    ClkMux I__12140 (
            .O(N__49669),
            .I(N__49206));
    ClkMux I__12139 (
            .O(N__49668),
            .I(N__49206));
    ClkMux I__12138 (
            .O(N__49667),
            .I(N__49206));
    ClkMux I__12137 (
            .O(N__49666),
            .I(N__49206));
    ClkMux I__12136 (
            .O(N__49665),
            .I(N__49206));
    GlobalMux I__12135 (
            .O(N__49206),
            .I(N__49203));
    gio2CtrlBuf I__12134 (
            .O(N__49203),
            .I(CLK_c));
    InMux I__12133 (
            .O(N__49200),
            .I(N__49197));
    LocalMux I__12132 (
            .O(N__49197),
            .I(N__49194));
    Span4Mux_v I__12131 (
            .O(N__49194),
            .I(N__49191));
    Span4Mux_s2_v I__12130 (
            .O(N__49191),
            .I(N__49188));
    Span4Mux_h I__12129 (
            .O(N__49188),
            .I(N__49185));
    Odrv4 I__12128 (
            .O(N__49185),
            .I(\c0.n22_adj_2373 ));
    CascadeMux I__12127 (
            .O(N__49182),
            .I(\c0.n18726_cascade_ ));
    InMux I__12126 (
            .O(N__49179),
            .I(N__49176));
    LocalMux I__12125 (
            .O(N__49176),
            .I(N__49173));
    Odrv12 I__12124 (
            .O(N__49173),
            .I(\c0.tx2.r_Tx_Data_0 ));
    InMux I__12123 (
            .O(N__49170),
            .I(N__49167));
    LocalMux I__12122 (
            .O(N__49167),
            .I(N__49164));
    Span4Mux_h I__12121 (
            .O(N__49164),
            .I(N__49161));
    Odrv4 I__12120 (
            .O(N__49161),
            .I(\c0.n18160 ));
    CascadeMux I__12119 (
            .O(N__49158),
            .I(N__49155));
    InMux I__12118 (
            .O(N__49155),
            .I(N__49152));
    LocalMux I__12117 (
            .O(N__49152),
            .I(\c0.n18161 ));
    InMux I__12116 (
            .O(N__49149),
            .I(N__49146));
    LocalMux I__12115 (
            .O(N__49146),
            .I(N__49143));
    Span4Mux_v I__12114 (
            .O(N__49143),
            .I(N__49140));
    Span4Mux_h I__12113 (
            .O(N__49140),
            .I(N__49137));
    Span4Mux_v I__12112 (
            .O(N__49137),
            .I(N__49134));
    Odrv4 I__12111 (
            .O(N__49134),
            .I(\c0.n18067 ));
    CascadeMux I__12110 (
            .O(N__49131),
            .I(\c0.n18771_cascade_ ));
    InMux I__12109 (
            .O(N__49128),
            .I(N__49125));
    LocalMux I__12108 (
            .O(N__49125),
            .I(N__49122));
    Span4Mux_h I__12107 (
            .O(N__49122),
            .I(N__49119));
    Odrv4 I__12106 (
            .O(N__49119),
            .I(\c0.n18068 ));
    InMux I__12105 (
            .O(N__49116),
            .I(N__49100));
    InMux I__12104 (
            .O(N__49115),
            .I(N__49100));
    InMux I__12103 (
            .O(N__49114),
            .I(N__49100));
    InMux I__12102 (
            .O(N__49113),
            .I(N__49087));
    InMux I__12101 (
            .O(N__49112),
            .I(N__49087));
    InMux I__12100 (
            .O(N__49111),
            .I(N__49087));
    InMux I__12099 (
            .O(N__49110),
            .I(N__49080));
    InMux I__12098 (
            .O(N__49109),
            .I(N__49080));
    InMux I__12097 (
            .O(N__49108),
            .I(N__49080));
    InMux I__12096 (
            .O(N__49107),
            .I(N__49077));
    LocalMux I__12095 (
            .O(N__49100),
            .I(N__49071));
    InMux I__12094 (
            .O(N__49099),
            .I(N__49064));
    InMux I__12093 (
            .O(N__49098),
            .I(N__49064));
    InMux I__12092 (
            .O(N__49097),
            .I(N__49064));
    InMux I__12091 (
            .O(N__49096),
            .I(N__49057));
    InMux I__12090 (
            .O(N__49095),
            .I(N__49057));
    InMux I__12089 (
            .O(N__49094),
            .I(N__49057));
    LocalMux I__12088 (
            .O(N__49087),
            .I(N__49054));
    LocalMux I__12087 (
            .O(N__49080),
            .I(N__49051));
    LocalMux I__12086 (
            .O(N__49077),
            .I(N__49042));
    InMux I__12085 (
            .O(N__49076),
            .I(N__49035));
    InMux I__12084 (
            .O(N__49075),
            .I(N__49035));
    InMux I__12083 (
            .O(N__49074),
            .I(N__49035));
    Span4Mux_h I__12082 (
            .O(N__49071),
            .I(N__49028));
    LocalMux I__12081 (
            .O(N__49064),
            .I(N__49028));
    LocalMux I__12080 (
            .O(N__49057),
            .I(N__49028));
    Span4Mux_v I__12079 (
            .O(N__49054),
            .I(N__49022));
    Span4Mux_s2_v I__12078 (
            .O(N__49051),
            .I(N__49022));
    InMux I__12077 (
            .O(N__49050),
            .I(N__49015));
    InMux I__12076 (
            .O(N__49049),
            .I(N__49015));
    InMux I__12075 (
            .O(N__49048),
            .I(N__49015));
    InMux I__12074 (
            .O(N__49047),
            .I(N__49008));
    InMux I__12073 (
            .O(N__49046),
            .I(N__49008));
    InMux I__12072 (
            .O(N__49045),
            .I(N__49008));
    Span4Mux_v I__12071 (
            .O(N__49042),
            .I(N__49005));
    LocalMux I__12070 (
            .O(N__49035),
            .I(N__49002));
    Span4Mux_v I__12069 (
            .O(N__49028),
            .I(N__48999));
    InMux I__12068 (
            .O(N__49027),
            .I(N__48995));
    Span4Mux_h I__12067 (
            .O(N__49022),
            .I(N__48992));
    LocalMux I__12066 (
            .O(N__49015),
            .I(N__48987));
    LocalMux I__12065 (
            .O(N__49008),
            .I(N__48987));
    Span4Mux_h I__12064 (
            .O(N__49005),
            .I(N__48979));
    Span4Mux_s3_v I__12063 (
            .O(N__49002),
            .I(N__48979));
    Span4Mux_h I__12062 (
            .O(N__48999),
            .I(N__48979));
    InMux I__12061 (
            .O(N__48998),
            .I(N__48976));
    LocalMux I__12060 (
            .O(N__48995),
            .I(N__48969));
    Span4Mux_h I__12059 (
            .O(N__48992),
            .I(N__48969));
    Span4Mux_s2_v I__12058 (
            .O(N__48987),
            .I(N__48969));
    InMux I__12057 (
            .O(N__48986),
            .I(N__48966));
    Span4Mux_h I__12056 (
            .O(N__48979),
            .I(N__48961));
    LocalMux I__12055 (
            .O(N__48976),
            .I(N__48961));
    Odrv4 I__12054 (
            .O(N__48969),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__12053 (
            .O(N__48966),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__12052 (
            .O(N__48961),
            .I(\c0.byte_transmit_counter2_3 ));
    CascadeMux I__12051 (
            .O(N__48954),
            .I(\c0.n18774_cascade_ ));
    InMux I__12050 (
            .O(N__48951),
            .I(N__48944));
    InMux I__12049 (
            .O(N__48950),
            .I(N__48941));
    InMux I__12048 (
            .O(N__48949),
            .I(N__48938));
    InMux I__12047 (
            .O(N__48948),
            .I(N__48935));
    InMux I__12046 (
            .O(N__48947),
            .I(N__48932));
    LocalMux I__12045 (
            .O(N__48944),
            .I(N__48929));
    LocalMux I__12044 (
            .O(N__48941),
            .I(N__48918));
    LocalMux I__12043 (
            .O(N__48938),
            .I(N__48918));
    LocalMux I__12042 (
            .O(N__48935),
            .I(N__48913));
    LocalMux I__12041 (
            .O(N__48932),
            .I(N__48913));
    Span4Mux_s1_v I__12040 (
            .O(N__48929),
            .I(N__48910));
    InMux I__12039 (
            .O(N__48928),
            .I(N__48907));
    InMux I__12038 (
            .O(N__48927),
            .I(N__48904));
    InMux I__12037 (
            .O(N__48926),
            .I(N__48901));
    InMux I__12036 (
            .O(N__48925),
            .I(N__48898));
    InMux I__12035 (
            .O(N__48924),
            .I(N__48895));
    InMux I__12034 (
            .O(N__48923),
            .I(N__48892));
    Span4Mux_v I__12033 (
            .O(N__48918),
            .I(N__48888));
    Span4Mux_v I__12032 (
            .O(N__48913),
            .I(N__48883));
    Span4Mux_v I__12031 (
            .O(N__48910),
            .I(N__48883));
    LocalMux I__12030 (
            .O(N__48907),
            .I(N__48880));
    LocalMux I__12029 (
            .O(N__48904),
            .I(N__48875));
    LocalMux I__12028 (
            .O(N__48901),
            .I(N__48875));
    LocalMux I__12027 (
            .O(N__48898),
            .I(N__48872));
    LocalMux I__12026 (
            .O(N__48895),
            .I(N__48867));
    LocalMux I__12025 (
            .O(N__48892),
            .I(N__48867));
    InMux I__12024 (
            .O(N__48891),
            .I(N__48864));
    Sp12to4 I__12023 (
            .O(N__48888),
            .I(N__48857));
    Sp12to4 I__12022 (
            .O(N__48883),
            .I(N__48857));
    Span12Mux_s5_h I__12021 (
            .O(N__48880),
            .I(N__48857));
    Span4Mux_s2_v I__12020 (
            .O(N__48875),
            .I(N__48852));
    Span4Mux_h I__12019 (
            .O(N__48872),
            .I(N__48852));
    Span4Mux_h I__12018 (
            .O(N__48867),
            .I(N__48849));
    LocalMux I__12017 (
            .O(N__48864),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv12 I__12016 (
            .O(N__48857),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__12015 (
            .O(N__48852),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__12014 (
            .O(N__48849),
            .I(\c0.byte_transmit_counter2_4 ));
    InMux I__12013 (
            .O(N__48840),
            .I(N__48837));
    LocalMux I__12012 (
            .O(N__48837),
            .I(N__48834));
    Span12Mux_s6_h I__12011 (
            .O(N__48834),
            .I(N__48831));
    Odrv12 I__12010 (
            .O(N__48831),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CEMux I__12009 (
            .O(N__48828),
            .I(N__48825));
    LocalMux I__12008 (
            .O(N__48825),
            .I(N__48820));
    CEMux I__12007 (
            .O(N__48824),
            .I(N__48817));
    CEMux I__12006 (
            .O(N__48823),
            .I(N__48813));
    Span4Mux_v I__12005 (
            .O(N__48820),
            .I(N__48806));
    LocalMux I__12004 (
            .O(N__48817),
            .I(N__48806));
    CEMux I__12003 (
            .O(N__48816),
            .I(N__48803));
    LocalMux I__12002 (
            .O(N__48813),
            .I(N__48800));
    CEMux I__12001 (
            .O(N__48812),
            .I(N__48797));
    CEMux I__12000 (
            .O(N__48811),
            .I(N__48793));
    Span4Mux_v I__11999 (
            .O(N__48806),
            .I(N__48790));
    LocalMux I__11998 (
            .O(N__48803),
            .I(N__48787));
    Span4Mux_v I__11997 (
            .O(N__48800),
            .I(N__48783));
    LocalMux I__11996 (
            .O(N__48797),
            .I(N__48780));
    CEMux I__11995 (
            .O(N__48796),
            .I(N__48777));
    LocalMux I__11994 (
            .O(N__48793),
            .I(N__48774));
    Span4Mux_h I__11993 (
            .O(N__48790),
            .I(N__48771));
    Span4Mux_v I__11992 (
            .O(N__48787),
            .I(N__48768));
    CEMux I__11991 (
            .O(N__48786),
            .I(N__48765));
    Span4Mux_h I__11990 (
            .O(N__48783),
            .I(N__48762));
    Span4Mux_h I__11989 (
            .O(N__48780),
            .I(N__48757));
    LocalMux I__11988 (
            .O(N__48777),
            .I(N__48757));
    Span4Mux_h I__11987 (
            .O(N__48774),
            .I(N__48754));
    Span4Mux_h I__11986 (
            .O(N__48771),
            .I(N__48751));
    Span4Mux_h I__11985 (
            .O(N__48768),
            .I(N__48748));
    LocalMux I__11984 (
            .O(N__48765),
            .I(N__48745));
    Span4Mux_h I__11983 (
            .O(N__48762),
            .I(N__48742));
    Span4Mux_h I__11982 (
            .O(N__48757),
            .I(N__48737));
    Span4Mux_h I__11981 (
            .O(N__48754),
            .I(N__48737));
    Span4Mux_v I__11980 (
            .O(N__48751),
            .I(N__48734));
    Span4Mux_h I__11979 (
            .O(N__48748),
            .I(N__48731));
    Span4Mux_h I__11978 (
            .O(N__48745),
            .I(N__48726));
    Span4Mux_v I__11977 (
            .O(N__48742),
            .I(N__48726));
    Odrv4 I__11976 (
            .O(N__48737),
            .I(\c0.tx2.n9639 ));
    Odrv4 I__11975 (
            .O(N__48734),
            .I(\c0.tx2.n9639 ));
    Odrv4 I__11974 (
            .O(N__48731),
            .I(\c0.tx2.n9639 ));
    Odrv4 I__11973 (
            .O(N__48726),
            .I(\c0.tx2.n9639 ));
    InMux I__11972 (
            .O(N__48717),
            .I(N__48714));
    LocalMux I__11971 (
            .O(N__48714),
            .I(N__48711));
    Span4Mux_v I__11970 (
            .O(N__48711),
            .I(N__48708));
    Odrv4 I__11969 (
            .O(N__48708),
            .I(\c0.n18669 ));
    InMux I__11968 (
            .O(N__48705),
            .I(N__48697));
    CascadeMux I__11967 (
            .O(N__48704),
            .I(N__48675));
    CascadeMux I__11966 (
            .O(N__48703),
            .I(N__48672));
    CascadeMux I__11965 (
            .O(N__48702),
            .I(N__48669));
    CascadeMux I__11964 (
            .O(N__48701),
            .I(N__48666));
    CascadeMux I__11963 (
            .O(N__48700),
            .I(N__48663));
    LocalMux I__11962 (
            .O(N__48697),
            .I(N__48660));
    InMux I__11961 (
            .O(N__48696),
            .I(N__48653));
    InMux I__11960 (
            .O(N__48695),
            .I(N__48653));
    InMux I__11959 (
            .O(N__48694),
            .I(N__48653));
    CascadeMux I__11958 (
            .O(N__48693),
            .I(N__48650));
    InMux I__11957 (
            .O(N__48692),
            .I(N__48645));
    CascadeMux I__11956 (
            .O(N__48691),
            .I(N__48642));
    InMux I__11955 (
            .O(N__48690),
            .I(N__48639));
    CascadeMux I__11954 (
            .O(N__48689),
            .I(N__48632));
    CascadeMux I__11953 (
            .O(N__48688),
            .I(N__48628));
    CascadeMux I__11952 (
            .O(N__48687),
            .I(N__48625));
    InMux I__11951 (
            .O(N__48686),
            .I(N__48613));
    InMux I__11950 (
            .O(N__48685),
            .I(N__48613));
    CascadeMux I__11949 (
            .O(N__48684),
            .I(N__48610));
    CascadeMux I__11948 (
            .O(N__48683),
            .I(N__48599));
    CascadeMux I__11947 (
            .O(N__48682),
            .I(N__48596));
    CascadeMux I__11946 (
            .O(N__48681),
            .I(N__48592));
    InMux I__11945 (
            .O(N__48680),
            .I(N__48586));
    InMux I__11944 (
            .O(N__48679),
            .I(N__48586));
    InMux I__11943 (
            .O(N__48678),
            .I(N__48579));
    InMux I__11942 (
            .O(N__48675),
            .I(N__48579));
    InMux I__11941 (
            .O(N__48672),
            .I(N__48579));
    InMux I__11940 (
            .O(N__48669),
            .I(N__48574));
    InMux I__11939 (
            .O(N__48666),
            .I(N__48574));
    InMux I__11938 (
            .O(N__48663),
            .I(N__48571));
    Span4Mux_v I__11937 (
            .O(N__48660),
            .I(N__48565));
    LocalMux I__11936 (
            .O(N__48653),
            .I(N__48565));
    InMux I__11935 (
            .O(N__48650),
            .I(N__48562));
    CascadeMux I__11934 (
            .O(N__48649),
            .I(N__48559));
    CascadeMux I__11933 (
            .O(N__48648),
            .I(N__48553));
    LocalMux I__11932 (
            .O(N__48645),
            .I(N__48550));
    InMux I__11931 (
            .O(N__48642),
            .I(N__48547));
    LocalMux I__11930 (
            .O(N__48639),
            .I(N__48544));
    InMux I__11929 (
            .O(N__48638),
            .I(N__48539));
    InMux I__11928 (
            .O(N__48637),
            .I(N__48539));
    InMux I__11927 (
            .O(N__48636),
            .I(N__48532));
    InMux I__11926 (
            .O(N__48635),
            .I(N__48532));
    InMux I__11925 (
            .O(N__48632),
            .I(N__48532));
    InMux I__11924 (
            .O(N__48631),
            .I(N__48525));
    InMux I__11923 (
            .O(N__48628),
            .I(N__48525));
    InMux I__11922 (
            .O(N__48625),
            .I(N__48525));
    InMux I__11921 (
            .O(N__48624),
            .I(N__48521));
    InMux I__11920 (
            .O(N__48623),
            .I(N__48518));
    InMux I__11919 (
            .O(N__48622),
            .I(N__48515));
    InMux I__11918 (
            .O(N__48621),
            .I(N__48510));
    InMux I__11917 (
            .O(N__48620),
            .I(N__48510));
    InMux I__11916 (
            .O(N__48619),
            .I(N__48505));
    InMux I__11915 (
            .O(N__48618),
            .I(N__48505));
    LocalMux I__11914 (
            .O(N__48613),
            .I(N__48502));
    InMux I__11913 (
            .O(N__48610),
            .I(N__48497));
    InMux I__11912 (
            .O(N__48609),
            .I(N__48497));
    InMux I__11911 (
            .O(N__48608),
            .I(N__48492));
    InMux I__11910 (
            .O(N__48607),
            .I(N__48492));
    CascadeMux I__11909 (
            .O(N__48606),
            .I(N__48484));
    InMux I__11908 (
            .O(N__48605),
            .I(N__48475));
    InMux I__11907 (
            .O(N__48604),
            .I(N__48475));
    InMux I__11906 (
            .O(N__48603),
            .I(N__48470));
    InMux I__11905 (
            .O(N__48602),
            .I(N__48470));
    InMux I__11904 (
            .O(N__48599),
            .I(N__48459));
    InMux I__11903 (
            .O(N__48596),
            .I(N__48459));
    InMux I__11902 (
            .O(N__48595),
            .I(N__48459));
    InMux I__11901 (
            .O(N__48592),
            .I(N__48459));
    InMux I__11900 (
            .O(N__48591),
            .I(N__48459));
    LocalMux I__11899 (
            .O(N__48586),
            .I(N__48454));
    LocalMux I__11898 (
            .O(N__48579),
            .I(N__48454));
    LocalMux I__11897 (
            .O(N__48574),
            .I(N__48449));
    LocalMux I__11896 (
            .O(N__48571),
            .I(N__48449));
    CascadeMux I__11895 (
            .O(N__48570),
            .I(N__48446));
    Span4Mux_v I__11894 (
            .O(N__48565),
            .I(N__48441));
    LocalMux I__11893 (
            .O(N__48562),
            .I(N__48441));
    InMux I__11892 (
            .O(N__48559),
            .I(N__48438));
    InMux I__11891 (
            .O(N__48558),
            .I(N__48429));
    InMux I__11890 (
            .O(N__48557),
            .I(N__48429));
    InMux I__11889 (
            .O(N__48556),
            .I(N__48429));
    InMux I__11888 (
            .O(N__48553),
            .I(N__48429));
    Span4Mux_v I__11887 (
            .O(N__48550),
            .I(N__48424));
    LocalMux I__11886 (
            .O(N__48547),
            .I(N__48424));
    Span4Mux_v I__11885 (
            .O(N__48544),
            .I(N__48415));
    LocalMux I__11884 (
            .O(N__48539),
            .I(N__48415));
    LocalMux I__11883 (
            .O(N__48532),
            .I(N__48415));
    LocalMux I__11882 (
            .O(N__48525),
            .I(N__48415));
    InMux I__11881 (
            .O(N__48524),
            .I(N__48412));
    LocalMux I__11880 (
            .O(N__48521),
            .I(N__48407));
    LocalMux I__11879 (
            .O(N__48518),
            .I(N__48407));
    LocalMux I__11878 (
            .O(N__48515),
            .I(N__48404));
    LocalMux I__11877 (
            .O(N__48510),
            .I(N__48399));
    LocalMux I__11876 (
            .O(N__48505),
            .I(N__48390));
    Span4Mux_s3_v I__11875 (
            .O(N__48502),
            .I(N__48390));
    LocalMux I__11874 (
            .O(N__48497),
            .I(N__48390));
    LocalMux I__11873 (
            .O(N__48492),
            .I(N__48390));
    CascadeMux I__11872 (
            .O(N__48491),
            .I(N__48386));
    CascadeMux I__11871 (
            .O(N__48490),
            .I(N__48383));
    InMux I__11870 (
            .O(N__48489),
            .I(N__48378));
    InMux I__11869 (
            .O(N__48488),
            .I(N__48378));
    InMux I__11868 (
            .O(N__48487),
            .I(N__48373));
    InMux I__11867 (
            .O(N__48484),
            .I(N__48373));
    InMux I__11866 (
            .O(N__48483),
            .I(N__48367));
    InMux I__11865 (
            .O(N__48482),
            .I(N__48367));
    InMux I__11864 (
            .O(N__48481),
            .I(N__48362));
    InMux I__11863 (
            .O(N__48480),
            .I(N__48362));
    LocalMux I__11862 (
            .O(N__48475),
            .I(N__48355));
    LocalMux I__11861 (
            .O(N__48470),
            .I(N__48355));
    LocalMux I__11860 (
            .O(N__48459),
            .I(N__48355));
    Span4Mux_h I__11859 (
            .O(N__48454),
            .I(N__48352));
    Span4Mux_h I__11858 (
            .O(N__48449),
            .I(N__48349));
    InMux I__11857 (
            .O(N__48446),
            .I(N__48346));
    Span4Mux_h I__11856 (
            .O(N__48441),
            .I(N__48343));
    LocalMux I__11855 (
            .O(N__48438),
            .I(N__48332));
    LocalMux I__11854 (
            .O(N__48429),
            .I(N__48332));
    Span4Mux_h I__11853 (
            .O(N__48424),
            .I(N__48332));
    Span4Mux_v I__11852 (
            .O(N__48415),
            .I(N__48332));
    LocalMux I__11851 (
            .O(N__48412),
            .I(N__48332));
    Span4Mux_s3_v I__11850 (
            .O(N__48407),
            .I(N__48329));
    Span4Mux_s3_v I__11849 (
            .O(N__48404),
            .I(N__48326));
    InMux I__11848 (
            .O(N__48403),
            .I(N__48321));
    InMux I__11847 (
            .O(N__48402),
            .I(N__48321));
    Span4Mux_v I__11846 (
            .O(N__48399),
            .I(N__48316));
    Span4Mux_v I__11845 (
            .O(N__48390),
            .I(N__48316));
    InMux I__11844 (
            .O(N__48389),
            .I(N__48311));
    InMux I__11843 (
            .O(N__48386),
            .I(N__48311));
    InMux I__11842 (
            .O(N__48383),
            .I(N__48308));
    LocalMux I__11841 (
            .O(N__48378),
            .I(N__48303));
    LocalMux I__11840 (
            .O(N__48373),
            .I(N__48303));
    InMux I__11839 (
            .O(N__48372),
            .I(N__48300));
    LocalMux I__11838 (
            .O(N__48367),
            .I(N__48295));
    LocalMux I__11837 (
            .O(N__48362),
            .I(N__48295));
    Span4Mux_h I__11836 (
            .O(N__48355),
            .I(N__48292));
    Span4Mux_v I__11835 (
            .O(N__48352),
            .I(N__48287));
    Span4Mux_v I__11834 (
            .O(N__48349),
            .I(N__48287));
    LocalMux I__11833 (
            .O(N__48346),
            .I(N__48283));
    Span4Mux_h I__11832 (
            .O(N__48343),
            .I(N__48278));
    Span4Mux_h I__11831 (
            .O(N__48332),
            .I(N__48278));
    Span4Mux_v I__11830 (
            .O(N__48329),
            .I(N__48273));
    Span4Mux_v I__11829 (
            .O(N__48326),
            .I(N__48273));
    LocalMux I__11828 (
            .O(N__48321),
            .I(N__48266));
    Sp12to4 I__11827 (
            .O(N__48316),
            .I(N__48266));
    LocalMux I__11826 (
            .O(N__48311),
            .I(N__48266));
    LocalMux I__11825 (
            .O(N__48308),
            .I(N__48259));
    Sp12to4 I__11824 (
            .O(N__48303),
            .I(N__48259));
    LocalMux I__11823 (
            .O(N__48300),
            .I(N__48259));
    Span4Mux_v I__11822 (
            .O(N__48295),
            .I(N__48252));
    Span4Mux_v I__11821 (
            .O(N__48292),
            .I(N__48252));
    Span4Mux_h I__11820 (
            .O(N__48287),
            .I(N__48252));
    InMux I__11819 (
            .O(N__48286),
            .I(N__48249));
    Span4Mux_h I__11818 (
            .O(N__48283),
            .I(N__48246));
    Span4Mux_h I__11817 (
            .O(N__48278),
            .I(N__48243));
    Sp12to4 I__11816 (
            .O(N__48273),
            .I(N__48236));
    Span12Mux_h I__11815 (
            .O(N__48266),
            .I(N__48236));
    Span12Mux_s7_v I__11814 (
            .O(N__48259),
            .I(N__48236));
    Span4Mux_h I__11813 (
            .O(N__48252),
            .I(N__48233));
    LocalMux I__11812 (
            .O(N__48249),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11811 (
            .O(N__48246),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11810 (
            .O(N__48243),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__11809 (
            .O(N__48236),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__11808 (
            .O(N__48233),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__11807 (
            .O(N__48222),
            .I(N__48216));
    InMux I__11806 (
            .O(N__48221),
            .I(N__48213));
    InMux I__11805 (
            .O(N__48220),
            .I(N__48210));
    InMux I__11804 (
            .O(N__48219),
            .I(N__48207));
    LocalMux I__11803 (
            .O(N__48216),
            .I(N__48204));
    LocalMux I__11802 (
            .O(N__48213),
            .I(N__48201));
    LocalMux I__11801 (
            .O(N__48210),
            .I(N__48198));
    LocalMux I__11800 (
            .O(N__48207),
            .I(N__48193));
    Span4Mux_v I__11799 (
            .O(N__48204),
            .I(N__48193));
    Span4Mux_h I__11798 (
            .O(N__48201),
            .I(N__48190));
    Span4Mux_s1_v I__11797 (
            .O(N__48198),
            .I(N__48187));
    Odrv4 I__11796 (
            .O(N__48193),
            .I(data_out_frame2_16_4));
    Odrv4 I__11795 (
            .O(N__48190),
            .I(data_out_frame2_16_4));
    Odrv4 I__11794 (
            .O(N__48187),
            .I(data_out_frame2_16_4));
    InMux I__11793 (
            .O(N__48180),
            .I(N__48177));
    LocalMux I__11792 (
            .O(N__48177),
            .I(N__48174));
    Odrv12 I__11791 (
            .O(N__48174),
            .I(\c0.data_out_frame2_20_4 ));
    InMux I__11790 (
            .O(N__48171),
            .I(N__48165));
    InMux I__11789 (
            .O(N__48170),
            .I(N__48162));
    InMux I__11788 (
            .O(N__48169),
            .I(N__48158));
    InMux I__11787 (
            .O(N__48168),
            .I(N__48154));
    LocalMux I__11786 (
            .O(N__48165),
            .I(N__48149));
    LocalMux I__11785 (
            .O(N__48162),
            .I(N__48149));
    InMux I__11784 (
            .O(N__48161),
            .I(N__48146));
    LocalMux I__11783 (
            .O(N__48158),
            .I(N__48143));
    InMux I__11782 (
            .O(N__48157),
            .I(N__48140));
    LocalMux I__11781 (
            .O(N__48154),
            .I(N__48135));
    Span4Mux_h I__11780 (
            .O(N__48149),
            .I(N__48130));
    LocalMux I__11779 (
            .O(N__48146),
            .I(N__48130));
    Span4Mux_s2_v I__11778 (
            .O(N__48143),
            .I(N__48127));
    LocalMux I__11777 (
            .O(N__48140),
            .I(N__48124));
    InMux I__11776 (
            .O(N__48139),
            .I(N__48121));
    InMux I__11775 (
            .O(N__48138),
            .I(N__48118));
    Span4Mux_s3_v I__11774 (
            .O(N__48135),
            .I(N__48115));
    Sp12to4 I__11773 (
            .O(N__48130),
            .I(N__48112));
    Span4Mux_v I__11772 (
            .O(N__48127),
            .I(N__48105));
    Span4Mux_v I__11771 (
            .O(N__48124),
            .I(N__48105));
    LocalMux I__11770 (
            .O(N__48121),
            .I(N__48105));
    LocalMux I__11769 (
            .O(N__48118),
            .I(N__48102));
    Span4Mux_h I__11768 (
            .O(N__48115),
            .I(N__48099));
    Span12Mux_s7_v I__11767 (
            .O(N__48112),
            .I(N__48096));
    Span4Mux_h I__11766 (
            .O(N__48105),
            .I(N__48093));
    Odrv4 I__11765 (
            .O(N__48102),
            .I(\c0.n7263 ));
    Odrv4 I__11764 (
            .O(N__48099),
            .I(\c0.n7263 ));
    Odrv12 I__11763 (
            .O(N__48096),
            .I(\c0.n7263 ));
    Odrv4 I__11762 (
            .O(N__48093),
            .I(\c0.n7263 ));
    CascadeMux I__11761 (
            .O(N__48084),
            .I(\c0.n18672_cascade_ ));
    InMux I__11760 (
            .O(N__48081),
            .I(N__48072));
    InMux I__11759 (
            .O(N__48080),
            .I(N__48065));
    InMux I__11758 (
            .O(N__48079),
            .I(N__48065));
    InMux I__11757 (
            .O(N__48078),
            .I(N__48062));
    InMux I__11756 (
            .O(N__48077),
            .I(N__48057));
    InMux I__11755 (
            .O(N__48076),
            .I(N__48057));
    InMux I__11754 (
            .O(N__48075),
            .I(N__48054));
    LocalMux I__11753 (
            .O(N__48072),
            .I(N__48051));
    InMux I__11752 (
            .O(N__48071),
            .I(N__48046));
    InMux I__11751 (
            .O(N__48070),
            .I(N__48046));
    LocalMux I__11750 (
            .O(N__48065),
            .I(N__48043));
    LocalMux I__11749 (
            .O(N__48062),
            .I(N__48036));
    LocalMux I__11748 (
            .O(N__48057),
            .I(N__48036));
    LocalMux I__11747 (
            .O(N__48054),
            .I(N__48036));
    Span4Mux_v I__11746 (
            .O(N__48051),
            .I(N__48026));
    LocalMux I__11745 (
            .O(N__48046),
            .I(N__48023));
    Span4Mux_v I__11744 (
            .O(N__48043),
            .I(N__48018));
    Span4Mux_v I__11743 (
            .O(N__48036),
            .I(N__48018));
    InMux I__11742 (
            .O(N__48035),
            .I(N__48012));
    InMux I__11741 (
            .O(N__48034),
            .I(N__48012));
    CascadeMux I__11740 (
            .O(N__48033),
            .I(N__48009));
    InMux I__11739 (
            .O(N__48032),
            .I(N__48004));
    InMux I__11738 (
            .O(N__48031),
            .I(N__48004));
    InMux I__11737 (
            .O(N__48030),
            .I(N__47999));
    InMux I__11736 (
            .O(N__48029),
            .I(N__47999));
    Span4Mux_v I__11735 (
            .O(N__48026),
            .I(N__47994));
    Span4Mux_s1_v I__11734 (
            .O(N__48023),
            .I(N__47994));
    Span4Mux_h I__11733 (
            .O(N__48018),
            .I(N__47991));
    InMux I__11732 (
            .O(N__48017),
            .I(N__47988));
    LocalMux I__11731 (
            .O(N__48012),
            .I(N__47985));
    InMux I__11730 (
            .O(N__48009),
            .I(N__47982));
    LocalMux I__11729 (
            .O(N__48004),
            .I(N__47978));
    LocalMux I__11728 (
            .O(N__47999),
            .I(N__47972));
    Span4Mux_h I__11727 (
            .O(N__47994),
            .I(N__47972));
    Span4Mux_h I__11726 (
            .O(N__47991),
            .I(N__47969));
    LocalMux I__11725 (
            .O(N__47988),
            .I(N__47966));
    Span4Mux_s2_v I__11724 (
            .O(N__47985),
            .I(N__47961));
    LocalMux I__11723 (
            .O(N__47982),
            .I(N__47961));
    InMux I__11722 (
            .O(N__47981),
            .I(N__47957));
    Span4Mux_s1_v I__11721 (
            .O(N__47978),
            .I(N__47954));
    InMux I__11720 (
            .O(N__47977),
            .I(N__47951));
    Span4Mux_h I__11719 (
            .O(N__47972),
            .I(N__47944));
    Span4Mux_v I__11718 (
            .O(N__47969),
            .I(N__47944));
    Span4Mux_v I__11717 (
            .O(N__47966),
            .I(N__47944));
    Span4Mux_h I__11716 (
            .O(N__47961),
            .I(N__47941));
    InMux I__11715 (
            .O(N__47960),
            .I(N__47938));
    LocalMux I__11714 (
            .O(N__47957),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__11713 (
            .O(N__47954),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__11712 (
            .O(N__47951),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__11711 (
            .O(N__47944),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__11710 (
            .O(N__47941),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__11709 (
            .O(N__47938),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__11708 (
            .O(N__47925),
            .I(N__47922));
    LocalMux I__11707 (
            .O(N__47922),
            .I(\c0.n22_adj_2243 ));
    InMux I__11706 (
            .O(N__47919),
            .I(N__47916));
    LocalMux I__11705 (
            .O(N__47916),
            .I(N__47912));
    CascadeMux I__11704 (
            .O(N__47915),
            .I(N__47909));
    Span4Mux_h I__11703 (
            .O(N__47912),
            .I(N__47906));
    InMux I__11702 (
            .O(N__47909),
            .I(N__47903));
    Odrv4 I__11701 (
            .O(N__47906),
            .I(rand_setpoint_14));
    LocalMux I__11700 (
            .O(N__47903),
            .I(rand_setpoint_14));
    CEMux I__11699 (
            .O(N__47898),
            .I(N__47895));
    LocalMux I__11698 (
            .O(N__47895),
            .I(N__47890));
    InMux I__11697 (
            .O(N__47894),
            .I(N__47887));
    CEMux I__11696 (
            .O(N__47893),
            .I(N__47880));
    Span4Mux_v I__11695 (
            .O(N__47890),
            .I(N__47875));
    LocalMux I__11694 (
            .O(N__47887),
            .I(N__47875));
    InMux I__11693 (
            .O(N__47886),
            .I(N__47872));
    CEMux I__11692 (
            .O(N__47885),
            .I(N__47868));
    CEMux I__11691 (
            .O(N__47884),
            .I(N__47865));
    InMux I__11690 (
            .O(N__47883),
            .I(N__47862));
    LocalMux I__11689 (
            .O(N__47880),
            .I(N__47859));
    Span4Mux_h I__11688 (
            .O(N__47875),
            .I(N__47854));
    LocalMux I__11687 (
            .O(N__47872),
            .I(N__47854));
    InMux I__11686 (
            .O(N__47871),
            .I(N__47851));
    LocalMux I__11685 (
            .O(N__47868),
            .I(N__47848));
    LocalMux I__11684 (
            .O(N__47865),
            .I(N__47845));
    LocalMux I__11683 (
            .O(N__47862),
            .I(N__47842));
    Span4Mux_h I__11682 (
            .O(N__47859),
            .I(N__47839));
    Span4Mux_v I__11681 (
            .O(N__47854),
            .I(N__47834));
    LocalMux I__11680 (
            .O(N__47851),
            .I(N__47834));
    Span4Mux_v I__11679 (
            .O(N__47848),
            .I(N__47831));
    Span4Mux_h I__11678 (
            .O(N__47845),
            .I(N__47826));
    Span4Mux_v I__11677 (
            .O(N__47842),
            .I(N__47826));
    Span4Mux_h I__11676 (
            .O(N__47839),
            .I(N__47821));
    Span4Mux_h I__11675 (
            .O(N__47834),
            .I(N__47821));
    Odrv4 I__11674 (
            .O(N__47831),
            .I(\c0.n11016 ));
    Odrv4 I__11673 (
            .O(N__47826),
            .I(\c0.n11016 ));
    Odrv4 I__11672 (
            .O(N__47821),
            .I(\c0.n11016 ));
    CascadeMux I__11671 (
            .O(N__47814),
            .I(N__47811));
    InMux I__11670 (
            .O(N__47811),
            .I(N__47806));
    CascadeMux I__11669 (
            .O(N__47810),
            .I(N__47803));
    CascadeMux I__11668 (
            .O(N__47809),
            .I(N__47800));
    LocalMux I__11667 (
            .O(N__47806),
            .I(N__47795));
    InMux I__11666 (
            .O(N__47803),
            .I(N__47792));
    InMux I__11665 (
            .O(N__47800),
            .I(N__47788));
    CascadeMux I__11664 (
            .O(N__47799),
            .I(N__47785));
    CascadeMux I__11663 (
            .O(N__47798),
            .I(N__47782));
    Span4Mux_v I__11662 (
            .O(N__47795),
            .I(N__47777));
    LocalMux I__11661 (
            .O(N__47792),
            .I(N__47777));
    CascadeMux I__11660 (
            .O(N__47791),
            .I(N__47774));
    LocalMux I__11659 (
            .O(N__47788),
            .I(N__47771));
    InMux I__11658 (
            .O(N__47785),
            .I(N__47768));
    InMux I__11657 (
            .O(N__47782),
            .I(N__47765));
    Span4Mux_h I__11656 (
            .O(N__47777),
            .I(N__47762));
    InMux I__11655 (
            .O(N__47774),
            .I(N__47759));
    Span4Mux_h I__11654 (
            .O(N__47771),
            .I(N__47754));
    LocalMux I__11653 (
            .O(N__47768),
            .I(N__47754));
    LocalMux I__11652 (
            .O(N__47765),
            .I(N__47751));
    Span4Mux_v I__11651 (
            .O(N__47762),
            .I(N__47746));
    LocalMux I__11650 (
            .O(N__47759),
            .I(N__47746));
    Span4Mux_v I__11649 (
            .O(N__47754),
            .I(N__47741));
    Span4Mux_h I__11648 (
            .O(N__47751),
            .I(N__47741));
    Odrv4 I__11647 (
            .O(N__47746),
            .I(n2732));
    Odrv4 I__11646 (
            .O(N__47741),
            .I(n2732));
    InMux I__11645 (
            .O(N__47736),
            .I(N__47730));
    InMux I__11644 (
            .O(N__47735),
            .I(N__47727));
    InMux I__11643 (
            .O(N__47734),
            .I(N__47724));
    InMux I__11642 (
            .O(N__47733),
            .I(N__47720));
    LocalMux I__11641 (
            .O(N__47730),
            .I(N__47715));
    LocalMux I__11640 (
            .O(N__47727),
            .I(N__47715));
    LocalMux I__11639 (
            .O(N__47724),
            .I(N__47712));
    InMux I__11638 (
            .O(N__47723),
            .I(N__47709));
    LocalMux I__11637 (
            .O(N__47720),
            .I(N__47706));
    Span4Mux_v I__11636 (
            .O(N__47715),
            .I(N__47703));
    Span4Mux_h I__11635 (
            .O(N__47712),
            .I(N__47700));
    LocalMux I__11634 (
            .O(N__47709),
            .I(\c0.data_out_7_6 ));
    Odrv12 I__11633 (
            .O(N__47706),
            .I(\c0.data_out_7_6 ));
    Odrv4 I__11632 (
            .O(N__47703),
            .I(\c0.data_out_7_6 ));
    Odrv4 I__11631 (
            .O(N__47700),
            .I(\c0.data_out_7_6 ));
    CascadeMux I__11630 (
            .O(N__47691),
            .I(N__47682));
    InMux I__11629 (
            .O(N__47690),
            .I(N__47673));
    InMux I__11628 (
            .O(N__47689),
            .I(N__47665));
    InMux I__11627 (
            .O(N__47688),
            .I(N__47662));
    InMux I__11626 (
            .O(N__47687),
            .I(N__47655));
    InMux I__11625 (
            .O(N__47686),
            .I(N__47655));
    InMux I__11624 (
            .O(N__47685),
            .I(N__47652));
    InMux I__11623 (
            .O(N__47682),
            .I(N__47647));
    InMux I__11622 (
            .O(N__47681),
            .I(N__47647));
    InMux I__11621 (
            .O(N__47680),
            .I(N__47641));
    InMux I__11620 (
            .O(N__47679),
            .I(N__47641));
    InMux I__11619 (
            .O(N__47678),
            .I(N__47638));
    InMux I__11618 (
            .O(N__47677),
            .I(N__47635));
    InMux I__11617 (
            .O(N__47676),
            .I(N__47629));
    LocalMux I__11616 (
            .O(N__47673),
            .I(N__47626));
    CascadeMux I__11615 (
            .O(N__47672),
            .I(N__47622));
    InMux I__11614 (
            .O(N__47671),
            .I(N__47619));
    CascadeMux I__11613 (
            .O(N__47670),
            .I(N__47616));
    CascadeMux I__11612 (
            .O(N__47669),
            .I(N__47611));
    InMux I__11611 (
            .O(N__47668),
            .I(N__47607));
    LocalMux I__11610 (
            .O(N__47665),
            .I(N__47604));
    LocalMux I__11609 (
            .O(N__47662),
            .I(N__47599));
    InMux I__11608 (
            .O(N__47661),
            .I(N__47596));
    InMux I__11607 (
            .O(N__47660),
            .I(N__47593));
    LocalMux I__11606 (
            .O(N__47655),
            .I(N__47590));
    LocalMux I__11605 (
            .O(N__47652),
            .I(N__47587));
    LocalMux I__11604 (
            .O(N__47647),
            .I(N__47584));
    InMux I__11603 (
            .O(N__47646),
            .I(N__47581));
    LocalMux I__11602 (
            .O(N__47641),
            .I(N__47578));
    LocalMux I__11601 (
            .O(N__47638),
            .I(N__47573));
    LocalMux I__11600 (
            .O(N__47635),
            .I(N__47573));
    InMux I__11599 (
            .O(N__47634),
            .I(N__47570));
    InMux I__11598 (
            .O(N__47633),
            .I(N__47567));
    InMux I__11597 (
            .O(N__47632),
            .I(N__47564));
    LocalMux I__11596 (
            .O(N__47629),
            .I(N__47561));
    Span4Mux_h I__11595 (
            .O(N__47626),
            .I(N__47558));
    InMux I__11594 (
            .O(N__47625),
            .I(N__47555));
    InMux I__11593 (
            .O(N__47622),
            .I(N__47551));
    LocalMux I__11592 (
            .O(N__47619),
            .I(N__47546));
    InMux I__11591 (
            .O(N__47616),
            .I(N__47543));
    CascadeMux I__11590 (
            .O(N__47615),
            .I(N__47540));
    CascadeMux I__11589 (
            .O(N__47614),
            .I(N__47537));
    InMux I__11588 (
            .O(N__47611),
            .I(N__47533));
    InMux I__11587 (
            .O(N__47610),
            .I(N__47530));
    LocalMux I__11586 (
            .O(N__47607),
            .I(N__47527));
    Span4Mux_v I__11585 (
            .O(N__47604),
            .I(N__47524));
    InMux I__11584 (
            .O(N__47603),
            .I(N__47519));
    InMux I__11583 (
            .O(N__47602),
            .I(N__47519));
    Span4Mux_v I__11582 (
            .O(N__47599),
            .I(N__47512));
    LocalMux I__11581 (
            .O(N__47596),
            .I(N__47512));
    LocalMux I__11580 (
            .O(N__47593),
            .I(N__47512));
    Span4Mux_v I__11579 (
            .O(N__47590),
            .I(N__47509));
    Span4Mux_v I__11578 (
            .O(N__47587),
            .I(N__47506));
    Span4Mux_v I__11577 (
            .O(N__47584),
            .I(N__47495));
    LocalMux I__11576 (
            .O(N__47581),
            .I(N__47495));
    Span4Mux_v I__11575 (
            .O(N__47578),
            .I(N__47495));
    Span4Mux_v I__11574 (
            .O(N__47573),
            .I(N__47495));
    LocalMux I__11573 (
            .O(N__47570),
            .I(N__47495));
    LocalMux I__11572 (
            .O(N__47567),
            .I(N__47492));
    LocalMux I__11571 (
            .O(N__47564),
            .I(N__47483));
    Span12Mux_h I__11570 (
            .O(N__47561),
            .I(N__47483));
    Sp12to4 I__11569 (
            .O(N__47558),
            .I(N__47483));
    LocalMux I__11568 (
            .O(N__47555),
            .I(N__47483));
    InMux I__11567 (
            .O(N__47554),
            .I(N__47480));
    LocalMux I__11566 (
            .O(N__47551),
            .I(N__47477));
    InMux I__11565 (
            .O(N__47550),
            .I(N__47474));
    InMux I__11564 (
            .O(N__47549),
            .I(N__47471));
    Span4Mux_h I__11563 (
            .O(N__47546),
            .I(N__47466));
    LocalMux I__11562 (
            .O(N__47543),
            .I(N__47466));
    InMux I__11561 (
            .O(N__47540),
            .I(N__47463));
    InMux I__11560 (
            .O(N__47537),
            .I(N__47458));
    InMux I__11559 (
            .O(N__47536),
            .I(N__47458));
    LocalMux I__11558 (
            .O(N__47533),
            .I(N__47439));
    LocalMux I__11557 (
            .O(N__47530),
            .I(N__47439));
    Span4Mux_v I__11556 (
            .O(N__47527),
            .I(N__47439));
    Span4Mux_h I__11555 (
            .O(N__47524),
            .I(N__47439));
    LocalMux I__11554 (
            .O(N__47519),
            .I(N__47439));
    Span4Mux_v I__11553 (
            .O(N__47512),
            .I(N__47439));
    Span4Mux_h I__11552 (
            .O(N__47509),
            .I(N__47439));
    Span4Mux_h I__11551 (
            .O(N__47506),
            .I(N__47439));
    Span4Mux_v I__11550 (
            .O(N__47495),
            .I(N__47439));
    Span12Mux_v I__11549 (
            .O(N__47492),
            .I(N__47436));
    Span12Mux_v I__11548 (
            .O(N__47483),
            .I(N__47433));
    LocalMux I__11547 (
            .O(N__47480),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11546 (
            .O(N__47477),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11545 (
            .O(N__47474),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11544 (
            .O(N__47471),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11543 (
            .O(N__47466),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11542 (
            .O(N__47463),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11541 (
            .O(N__47458),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11540 (
            .O(N__47439),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__11539 (
            .O(N__47436),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__11538 (
            .O(N__47433),
            .I(UART_TRANSMITTER_state_2));
    InMux I__11537 (
            .O(N__47412),
            .I(N__47395));
    InMux I__11536 (
            .O(N__47411),
            .I(N__47391));
    InMux I__11535 (
            .O(N__47410),
            .I(N__47388));
    InMux I__11534 (
            .O(N__47409),
            .I(N__47381));
    InMux I__11533 (
            .O(N__47408),
            .I(N__47381));
    InMux I__11532 (
            .O(N__47407),
            .I(N__47381));
    InMux I__11531 (
            .O(N__47406),
            .I(N__47375));
    InMux I__11530 (
            .O(N__47405),
            .I(N__47375));
    InMux I__11529 (
            .O(N__47404),
            .I(N__47372));
    InMux I__11528 (
            .O(N__47403),
            .I(N__47369));
    InMux I__11527 (
            .O(N__47402),
            .I(N__47366));
    InMux I__11526 (
            .O(N__47401),
            .I(N__47362));
    InMux I__11525 (
            .O(N__47400),
            .I(N__47359));
    InMux I__11524 (
            .O(N__47399),
            .I(N__47350));
    InMux I__11523 (
            .O(N__47398),
            .I(N__47347));
    LocalMux I__11522 (
            .O(N__47395),
            .I(N__47342));
    InMux I__11521 (
            .O(N__47394),
            .I(N__47339));
    LocalMux I__11520 (
            .O(N__47391),
            .I(N__47332));
    LocalMux I__11519 (
            .O(N__47388),
            .I(N__47332));
    LocalMux I__11518 (
            .O(N__47381),
            .I(N__47332));
    InMux I__11517 (
            .O(N__47380),
            .I(N__47329));
    LocalMux I__11516 (
            .O(N__47375),
            .I(N__47324));
    LocalMux I__11515 (
            .O(N__47372),
            .I(N__47324));
    LocalMux I__11514 (
            .O(N__47369),
            .I(N__47321));
    LocalMux I__11513 (
            .O(N__47366),
            .I(N__47317));
    InMux I__11512 (
            .O(N__47365),
            .I(N__47314));
    LocalMux I__11511 (
            .O(N__47362),
            .I(N__47308));
    LocalMux I__11510 (
            .O(N__47359),
            .I(N__47308));
    InMux I__11509 (
            .O(N__47358),
            .I(N__47299));
    InMux I__11508 (
            .O(N__47357),
            .I(N__47299));
    InMux I__11507 (
            .O(N__47356),
            .I(N__47299));
    InMux I__11506 (
            .O(N__47355),
            .I(N__47299));
    InMux I__11505 (
            .O(N__47354),
            .I(N__47294));
    InMux I__11504 (
            .O(N__47353),
            .I(N__47294));
    LocalMux I__11503 (
            .O(N__47350),
            .I(N__47288));
    LocalMux I__11502 (
            .O(N__47347),
            .I(N__47285));
    InMux I__11501 (
            .O(N__47346),
            .I(N__47282));
    InMux I__11500 (
            .O(N__47345),
            .I(N__47279));
    Span4Mux_v I__11499 (
            .O(N__47342),
            .I(N__47276));
    LocalMux I__11498 (
            .O(N__47339),
            .I(N__47273));
    Span4Mux_v I__11497 (
            .O(N__47332),
            .I(N__47264));
    LocalMux I__11496 (
            .O(N__47329),
            .I(N__47264));
    Span4Mux_v I__11495 (
            .O(N__47324),
            .I(N__47264));
    Span4Mux_h I__11494 (
            .O(N__47321),
            .I(N__47264));
    InMux I__11493 (
            .O(N__47320),
            .I(N__47261));
    Span4Mux_v I__11492 (
            .O(N__47317),
            .I(N__47249));
    LocalMux I__11491 (
            .O(N__47314),
            .I(N__47249));
    InMux I__11490 (
            .O(N__47313),
            .I(N__47246));
    Span4Mux_v I__11489 (
            .O(N__47308),
            .I(N__47243));
    LocalMux I__11488 (
            .O(N__47299),
            .I(N__47238));
    LocalMux I__11487 (
            .O(N__47294),
            .I(N__47238));
    InMux I__11486 (
            .O(N__47293),
            .I(N__47229));
    InMux I__11485 (
            .O(N__47292),
            .I(N__47229));
    InMux I__11484 (
            .O(N__47291),
            .I(N__47229));
    Span4Mux_h I__11483 (
            .O(N__47288),
            .I(N__47225));
    Span4Mux_h I__11482 (
            .O(N__47285),
            .I(N__47210));
    LocalMux I__11481 (
            .O(N__47282),
            .I(N__47210));
    LocalMux I__11480 (
            .O(N__47279),
            .I(N__47210));
    Span4Mux_h I__11479 (
            .O(N__47276),
            .I(N__47210));
    Span4Mux_h I__11478 (
            .O(N__47273),
            .I(N__47210));
    Span4Mux_h I__11477 (
            .O(N__47264),
            .I(N__47210));
    LocalMux I__11476 (
            .O(N__47261),
            .I(N__47210));
    InMux I__11475 (
            .O(N__47260),
            .I(N__47205));
    InMux I__11474 (
            .O(N__47259),
            .I(N__47205));
    InMux I__11473 (
            .O(N__47258),
            .I(N__47202));
    InMux I__11472 (
            .O(N__47257),
            .I(N__47197));
    InMux I__11471 (
            .O(N__47256),
            .I(N__47197));
    InMux I__11470 (
            .O(N__47255),
            .I(N__47192));
    InMux I__11469 (
            .O(N__47254),
            .I(N__47192));
    Span4Mux_v I__11468 (
            .O(N__47249),
            .I(N__47183));
    LocalMux I__11467 (
            .O(N__47246),
            .I(N__47183));
    Span4Mux_v I__11466 (
            .O(N__47243),
            .I(N__47183));
    Span4Mux_v I__11465 (
            .O(N__47238),
            .I(N__47183));
    InMux I__11464 (
            .O(N__47237),
            .I(N__47178));
    InMux I__11463 (
            .O(N__47236),
            .I(N__47178));
    LocalMux I__11462 (
            .O(N__47229),
            .I(N__47175));
    InMux I__11461 (
            .O(N__47228),
            .I(N__47172));
    Span4Mux_h I__11460 (
            .O(N__47225),
            .I(N__47167));
    Span4Mux_v I__11459 (
            .O(N__47210),
            .I(N__47167));
    LocalMux I__11458 (
            .O(N__47205),
            .I(N__47162));
    LocalMux I__11457 (
            .O(N__47202),
            .I(N__47162));
    LocalMux I__11456 (
            .O(N__47197),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11455 (
            .O(N__47192),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11454 (
            .O(N__47183),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11453 (
            .O(N__47178),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__11452 (
            .O(N__47175),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11451 (
            .O(N__47172),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11450 (
            .O(N__47167),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11449 (
            .O(N__47162),
            .I(UART_TRANSMITTER_state_0));
    InMux I__11448 (
            .O(N__47145),
            .I(N__47134));
    InMux I__11447 (
            .O(N__47144),
            .I(N__47131));
    InMux I__11446 (
            .O(N__47143),
            .I(N__47124));
    InMux I__11445 (
            .O(N__47142),
            .I(N__47112));
    InMux I__11444 (
            .O(N__47141),
            .I(N__47108));
    InMux I__11443 (
            .O(N__47140),
            .I(N__47105));
    InMux I__11442 (
            .O(N__47139),
            .I(N__47102));
    InMux I__11441 (
            .O(N__47138),
            .I(N__47097));
    InMux I__11440 (
            .O(N__47137),
            .I(N__47097));
    LocalMux I__11439 (
            .O(N__47134),
            .I(N__47092));
    LocalMux I__11438 (
            .O(N__47131),
            .I(N__47092));
    InMux I__11437 (
            .O(N__47130),
            .I(N__47089));
    InMux I__11436 (
            .O(N__47129),
            .I(N__47086));
    CascadeMux I__11435 (
            .O(N__47128),
            .I(N__47082));
    InMux I__11434 (
            .O(N__47127),
            .I(N__47077));
    LocalMux I__11433 (
            .O(N__47124),
            .I(N__47074));
    InMux I__11432 (
            .O(N__47123),
            .I(N__47067));
    InMux I__11431 (
            .O(N__47122),
            .I(N__47060));
    InMux I__11430 (
            .O(N__47121),
            .I(N__47055));
    InMux I__11429 (
            .O(N__47120),
            .I(N__47050));
    InMux I__11428 (
            .O(N__47119),
            .I(N__47050));
    InMux I__11427 (
            .O(N__47118),
            .I(N__47047));
    InMux I__11426 (
            .O(N__47117),
            .I(N__47040));
    InMux I__11425 (
            .O(N__47116),
            .I(N__47040));
    InMux I__11424 (
            .O(N__47115),
            .I(N__47040));
    LocalMux I__11423 (
            .O(N__47112),
            .I(N__47037));
    InMux I__11422 (
            .O(N__47111),
            .I(N__47034));
    LocalMux I__11421 (
            .O(N__47108),
            .I(N__47027));
    LocalMux I__11420 (
            .O(N__47105),
            .I(N__47027));
    LocalMux I__11419 (
            .O(N__47102),
            .I(N__47027));
    LocalMux I__11418 (
            .O(N__47097),
            .I(N__47024));
    Span4Mux_v I__11417 (
            .O(N__47092),
            .I(N__47019));
    LocalMux I__11416 (
            .O(N__47089),
            .I(N__47019));
    LocalMux I__11415 (
            .O(N__47086),
            .I(N__47016));
    InMux I__11414 (
            .O(N__47085),
            .I(N__47011));
    InMux I__11413 (
            .O(N__47082),
            .I(N__47011));
    InMux I__11412 (
            .O(N__47081),
            .I(N__47006));
    InMux I__11411 (
            .O(N__47080),
            .I(N__47006));
    LocalMux I__11410 (
            .O(N__47077),
            .I(N__47003));
    Span4Mux_h I__11409 (
            .O(N__47074),
            .I(N__47000));
    InMux I__11408 (
            .O(N__47073),
            .I(N__46995));
    InMux I__11407 (
            .O(N__47072),
            .I(N__46995));
    InMux I__11406 (
            .O(N__47071),
            .I(N__46990));
    InMux I__11405 (
            .O(N__47070),
            .I(N__46990));
    LocalMux I__11404 (
            .O(N__47067),
            .I(N__46987));
    InMux I__11403 (
            .O(N__47066),
            .I(N__46978));
    InMux I__11402 (
            .O(N__47065),
            .I(N__46978));
    InMux I__11401 (
            .O(N__47064),
            .I(N__46978));
    InMux I__11400 (
            .O(N__47063),
            .I(N__46978));
    LocalMux I__11399 (
            .O(N__47060),
            .I(N__46975));
    InMux I__11398 (
            .O(N__47059),
            .I(N__46963));
    InMux I__11397 (
            .O(N__47058),
            .I(N__46963));
    LocalMux I__11396 (
            .O(N__47055),
            .I(N__46945));
    LocalMux I__11395 (
            .O(N__47050),
            .I(N__46945));
    LocalMux I__11394 (
            .O(N__47047),
            .I(N__46945));
    LocalMux I__11393 (
            .O(N__47040),
            .I(N__46945));
    Span4Mux_h I__11392 (
            .O(N__47037),
            .I(N__46945));
    LocalMux I__11391 (
            .O(N__47034),
            .I(N__46945));
    Span4Mux_v I__11390 (
            .O(N__47027),
            .I(N__46940));
    Span4Mux_v I__11389 (
            .O(N__47024),
            .I(N__46940));
    Span4Mux_v I__11388 (
            .O(N__47019),
            .I(N__46933));
    Span4Mux_h I__11387 (
            .O(N__47016),
            .I(N__46933));
    LocalMux I__11386 (
            .O(N__47011),
            .I(N__46933));
    LocalMux I__11385 (
            .O(N__47006),
            .I(N__46922));
    Span4Mux_h I__11384 (
            .O(N__47003),
            .I(N__46922));
    Span4Mux_h I__11383 (
            .O(N__47000),
            .I(N__46922));
    LocalMux I__11382 (
            .O(N__46995),
            .I(N__46922));
    LocalMux I__11381 (
            .O(N__46990),
            .I(N__46922));
    Span12Mux_h I__11380 (
            .O(N__46987),
            .I(N__46919));
    LocalMux I__11379 (
            .O(N__46978),
            .I(N__46914));
    Span12Mux_v I__11378 (
            .O(N__46975),
            .I(N__46914));
    InMux I__11377 (
            .O(N__46974),
            .I(N__46899));
    InMux I__11376 (
            .O(N__46973),
            .I(N__46899));
    InMux I__11375 (
            .O(N__46972),
            .I(N__46899));
    InMux I__11374 (
            .O(N__46971),
            .I(N__46899));
    InMux I__11373 (
            .O(N__46970),
            .I(N__46899));
    InMux I__11372 (
            .O(N__46969),
            .I(N__46899));
    InMux I__11371 (
            .O(N__46968),
            .I(N__46899));
    LocalMux I__11370 (
            .O(N__46963),
            .I(N__46896));
    InMux I__11369 (
            .O(N__46962),
            .I(N__46891));
    InMux I__11368 (
            .O(N__46961),
            .I(N__46891));
    InMux I__11367 (
            .O(N__46960),
            .I(N__46884));
    InMux I__11366 (
            .O(N__46959),
            .I(N__46884));
    InMux I__11365 (
            .O(N__46958),
            .I(N__46884));
    Span4Mux_v I__11364 (
            .O(N__46945),
            .I(N__46879));
    Span4Mux_h I__11363 (
            .O(N__46940),
            .I(N__46879));
    Span4Mux_h I__11362 (
            .O(N__46933),
            .I(N__46874));
    Span4Mux_v I__11361 (
            .O(N__46922),
            .I(N__46874));
    Odrv12 I__11360 (
            .O(N__46919),
            .I(UART_TRANSMITTER_state_1));
    Odrv12 I__11359 (
            .O(N__46914),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11358 (
            .O(N__46899),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11357 (
            .O(N__46896),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11356 (
            .O(N__46891),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11355 (
            .O(N__46884),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11354 (
            .O(N__46879),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11353 (
            .O(N__46874),
            .I(UART_TRANSMITTER_state_1));
    CEMux I__11352 (
            .O(N__46857),
            .I(N__46848));
    CEMux I__11351 (
            .O(N__46856),
            .I(N__46840));
    InMux I__11350 (
            .O(N__46855),
            .I(N__46837));
    CEMux I__11349 (
            .O(N__46854),
            .I(N__46834));
    InMux I__11348 (
            .O(N__46853),
            .I(N__46831));
    InMux I__11347 (
            .O(N__46852),
            .I(N__46828));
    InMux I__11346 (
            .O(N__46851),
            .I(N__46825));
    LocalMux I__11345 (
            .O(N__46848),
            .I(N__46822));
    InMux I__11344 (
            .O(N__46847),
            .I(N__46818));
    InMux I__11343 (
            .O(N__46846),
            .I(N__46815));
    CEMux I__11342 (
            .O(N__46845),
            .I(N__46811));
    CEMux I__11341 (
            .O(N__46844),
            .I(N__46808));
    CEMux I__11340 (
            .O(N__46843),
            .I(N__46805));
    LocalMux I__11339 (
            .O(N__46840),
            .I(N__46802));
    LocalMux I__11338 (
            .O(N__46837),
            .I(N__46799));
    LocalMux I__11337 (
            .O(N__46834),
            .I(N__46792));
    LocalMux I__11336 (
            .O(N__46831),
            .I(N__46792));
    LocalMux I__11335 (
            .O(N__46828),
            .I(N__46792));
    LocalMux I__11334 (
            .O(N__46825),
            .I(N__46789));
    Span4Mux_v I__11333 (
            .O(N__46822),
            .I(N__46786));
    CEMux I__11332 (
            .O(N__46821),
            .I(N__46783));
    LocalMux I__11331 (
            .O(N__46818),
            .I(N__46778));
    LocalMux I__11330 (
            .O(N__46815),
            .I(N__46778));
    InMux I__11329 (
            .O(N__46814),
            .I(N__46775));
    LocalMux I__11328 (
            .O(N__46811),
            .I(N__46772));
    LocalMux I__11327 (
            .O(N__46808),
            .I(N__46769));
    LocalMux I__11326 (
            .O(N__46805),
            .I(N__46762));
    Span4Mux_v I__11325 (
            .O(N__46802),
            .I(N__46762));
    Span4Mux_h I__11324 (
            .O(N__46799),
            .I(N__46762));
    Span4Mux_v I__11323 (
            .O(N__46792),
            .I(N__46757));
    Span4Mux_v I__11322 (
            .O(N__46789),
            .I(N__46757));
    Span4Mux_h I__11321 (
            .O(N__46786),
            .I(N__46752));
    LocalMux I__11320 (
            .O(N__46783),
            .I(N__46752));
    Span4Mux_h I__11319 (
            .O(N__46778),
            .I(N__46747));
    LocalMux I__11318 (
            .O(N__46775),
            .I(N__46747));
    Span12Mux_h I__11317 (
            .O(N__46772),
            .I(N__46744));
    Span4Mux_h I__11316 (
            .O(N__46769),
            .I(N__46741));
    Span4Mux_h I__11315 (
            .O(N__46762),
            .I(N__46738));
    Span4Mux_h I__11314 (
            .O(N__46757),
            .I(N__46735));
    Span4Mux_h I__11313 (
            .O(N__46752),
            .I(N__46730));
    Span4Mux_h I__11312 (
            .O(N__46747),
            .I(N__46730));
    Odrv12 I__11311 (
            .O(N__46744),
            .I(data_out_10__7__N_110));
    Odrv4 I__11310 (
            .O(N__46741),
            .I(data_out_10__7__N_110));
    Odrv4 I__11309 (
            .O(N__46738),
            .I(data_out_10__7__N_110));
    Odrv4 I__11308 (
            .O(N__46735),
            .I(data_out_10__7__N_110));
    Odrv4 I__11307 (
            .O(N__46730),
            .I(data_out_10__7__N_110));
    CascadeMux I__11306 (
            .O(N__46719),
            .I(N__46716));
    InMux I__11305 (
            .O(N__46716),
            .I(N__46712));
    InMux I__11304 (
            .O(N__46715),
            .I(N__46709));
    LocalMux I__11303 (
            .O(N__46712),
            .I(N__46704));
    LocalMux I__11302 (
            .O(N__46709),
            .I(N__46701));
    CascadeMux I__11301 (
            .O(N__46708),
            .I(N__46698));
    InMux I__11300 (
            .O(N__46707),
            .I(N__46694));
    Span4Mux_h I__11299 (
            .O(N__46704),
            .I(N__46691));
    Span4Mux_v I__11298 (
            .O(N__46701),
            .I(N__46688));
    InMux I__11297 (
            .O(N__46698),
            .I(N__46685));
    InMux I__11296 (
            .O(N__46697),
            .I(N__46682));
    LocalMux I__11295 (
            .O(N__46694),
            .I(N__46679));
    Span4Mux_v I__11294 (
            .O(N__46691),
            .I(N__46676));
    Span4Mux_h I__11293 (
            .O(N__46688),
            .I(N__46671));
    LocalMux I__11292 (
            .O(N__46685),
            .I(N__46671));
    LocalMux I__11291 (
            .O(N__46682),
            .I(data_out_frame2_5_4));
    Odrv12 I__11290 (
            .O(N__46679),
            .I(data_out_frame2_5_4));
    Odrv4 I__11289 (
            .O(N__46676),
            .I(data_out_frame2_5_4));
    Odrv4 I__11288 (
            .O(N__46671),
            .I(data_out_frame2_5_4));
    InMux I__11287 (
            .O(N__46662),
            .I(N__46659));
    LocalMux I__11286 (
            .O(N__46659),
            .I(\c0.n17856 ));
    InMux I__11285 (
            .O(N__46656),
            .I(N__46649));
    InMux I__11284 (
            .O(N__46655),
            .I(N__46649));
    InMux I__11283 (
            .O(N__46654),
            .I(N__46646));
    LocalMux I__11282 (
            .O(N__46649),
            .I(N__46642));
    LocalMux I__11281 (
            .O(N__46646),
            .I(N__46639));
    CascadeMux I__11280 (
            .O(N__46645),
            .I(N__46634));
    Span4Mux_v I__11279 (
            .O(N__46642),
            .I(N__46629));
    Span4Mux_s3_v I__11278 (
            .O(N__46639),
            .I(N__46629));
    InMux I__11277 (
            .O(N__46638),
            .I(N__46626));
    InMux I__11276 (
            .O(N__46637),
            .I(N__46623));
    InMux I__11275 (
            .O(N__46634),
            .I(N__46620));
    Span4Mux_h I__11274 (
            .O(N__46629),
            .I(N__46615));
    LocalMux I__11273 (
            .O(N__46626),
            .I(N__46615));
    LocalMux I__11272 (
            .O(N__46623),
            .I(data_out_frame2_16_2));
    LocalMux I__11271 (
            .O(N__46620),
            .I(data_out_frame2_16_2));
    Odrv4 I__11270 (
            .O(N__46615),
            .I(data_out_frame2_16_2));
    CascadeMux I__11269 (
            .O(N__46608),
            .I(N__46605));
    InMux I__11268 (
            .O(N__46605),
            .I(N__46599));
    InMux I__11267 (
            .O(N__46604),
            .I(N__46599));
    LocalMux I__11266 (
            .O(N__46599),
            .I(N__46596));
    Span4Mux_h I__11265 (
            .O(N__46596),
            .I(N__46591));
    CascadeMux I__11264 (
            .O(N__46595),
            .I(N__46586));
    InMux I__11263 (
            .O(N__46594),
            .I(N__46583));
    Sp12to4 I__11262 (
            .O(N__46591),
            .I(N__46580));
    InMux I__11261 (
            .O(N__46590),
            .I(N__46575));
    InMux I__11260 (
            .O(N__46589),
            .I(N__46575));
    InMux I__11259 (
            .O(N__46586),
            .I(N__46572));
    LocalMux I__11258 (
            .O(N__46583),
            .I(data_out_frame2_9_2));
    Odrv12 I__11257 (
            .O(N__46580),
            .I(data_out_frame2_9_2));
    LocalMux I__11256 (
            .O(N__46575),
            .I(data_out_frame2_9_2));
    LocalMux I__11255 (
            .O(N__46572),
            .I(data_out_frame2_9_2));
    InMux I__11254 (
            .O(N__46563),
            .I(N__46559));
    InMux I__11253 (
            .O(N__46562),
            .I(N__46556));
    LocalMux I__11252 (
            .O(N__46559),
            .I(N__46553));
    LocalMux I__11251 (
            .O(N__46556),
            .I(N__46550));
    Odrv12 I__11250 (
            .O(N__46553),
            .I(\c0.n10887 ));
    Odrv4 I__11249 (
            .O(N__46550),
            .I(\c0.n10887 ));
    InMux I__11248 (
            .O(N__46545),
            .I(N__46542));
    LocalMux I__11247 (
            .O(N__46542),
            .I(N__46539));
    Odrv12 I__11246 (
            .O(N__46539),
            .I(\c0.n16_adj_2399 ));
    InMux I__11245 (
            .O(N__46536),
            .I(N__46530));
    InMux I__11244 (
            .O(N__46535),
            .I(N__46527));
    InMux I__11243 (
            .O(N__46534),
            .I(N__46524));
    InMux I__11242 (
            .O(N__46533),
            .I(N__46521));
    LocalMux I__11241 (
            .O(N__46530),
            .I(N__46517));
    LocalMux I__11240 (
            .O(N__46527),
            .I(N__46512));
    LocalMux I__11239 (
            .O(N__46524),
            .I(N__46512));
    LocalMux I__11238 (
            .O(N__46521),
            .I(N__46509));
    InMux I__11237 (
            .O(N__46520),
            .I(N__46506));
    Span4Mux_v I__11236 (
            .O(N__46517),
            .I(N__46503));
    Span4Mux_s3_v I__11235 (
            .O(N__46512),
            .I(N__46500));
    Span4Mux_h I__11234 (
            .O(N__46509),
            .I(N__46497));
    LocalMux I__11233 (
            .O(N__46506),
            .I(data_out_frame2_10_0));
    Odrv4 I__11232 (
            .O(N__46503),
            .I(data_out_frame2_10_0));
    Odrv4 I__11231 (
            .O(N__46500),
            .I(data_out_frame2_10_0));
    Odrv4 I__11230 (
            .O(N__46497),
            .I(data_out_frame2_10_0));
    CascadeMux I__11229 (
            .O(N__46488),
            .I(N__46482));
    InMux I__11228 (
            .O(N__46487),
            .I(N__46479));
    InMux I__11227 (
            .O(N__46486),
            .I(N__46476));
    InMux I__11226 (
            .O(N__46485),
            .I(N__46471));
    InMux I__11225 (
            .O(N__46482),
            .I(N__46468));
    LocalMux I__11224 (
            .O(N__46479),
            .I(N__46464));
    LocalMux I__11223 (
            .O(N__46476),
            .I(N__46461));
    InMux I__11222 (
            .O(N__46475),
            .I(N__46458));
    CascadeMux I__11221 (
            .O(N__46474),
            .I(N__46455));
    LocalMux I__11220 (
            .O(N__46471),
            .I(N__46452));
    LocalMux I__11219 (
            .O(N__46468),
            .I(N__46449));
    InMux I__11218 (
            .O(N__46467),
            .I(N__46446));
    Span4Mux_v I__11217 (
            .O(N__46464),
            .I(N__46443));
    Span4Mux_v I__11216 (
            .O(N__46461),
            .I(N__46440));
    LocalMux I__11215 (
            .O(N__46458),
            .I(N__46437));
    InMux I__11214 (
            .O(N__46455),
            .I(N__46434));
    Span4Mux_h I__11213 (
            .O(N__46452),
            .I(N__46429));
    Span4Mux_h I__11212 (
            .O(N__46449),
            .I(N__46429));
    LocalMux I__11211 (
            .O(N__46446),
            .I(data_out_frame2_11_0));
    Odrv4 I__11210 (
            .O(N__46443),
            .I(data_out_frame2_11_0));
    Odrv4 I__11209 (
            .O(N__46440),
            .I(data_out_frame2_11_0));
    Odrv4 I__11208 (
            .O(N__46437),
            .I(data_out_frame2_11_0));
    LocalMux I__11207 (
            .O(N__46434),
            .I(data_out_frame2_11_0));
    Odrv4 I__11206 (
            .O(N__46429),
            .I(data_out_frame2_11_0));
    InMux I__11205 (
            .O(N__46416),
            .I(N__46412));
    InMux I__11204 (
            .O(N__46415),
            .I(N__46407));
    LocalMux I__11203 (
            .O(N__46412),
            .I(N__46404));
    InMux I__11202 (
            .O(N__46411),
            .I(N__46401));
    InMux I__11201 (
            .O(N__46410),
            .I(N__46398));
    LocalMux I__11200 (
            .O(N__46407),
            .I(N__46394));
    Span4Mux_h I__11199 (
            .O(N__46404),
            .I(N__46389));
    LocalMux I__11198 (
            .O(N__46401),
            .I(N__46389));
    LocalMux I__11197 (
            .O(N__46398),
            .I(N__46386));
    InMux I__11196 (
            .O(N__46397),
            .I(N__46383));
    Span4Mux_s1_v I__11195 (
            .O(N__46394),
            .I(N__46379));
    Span4Mux_v I__11194 (
            .O(N__46389),
            .I(N__46372));
    Span4Mux_v I__11193 (
            .O(N__46386),
            .I(N__46372));
    LocalMux I__11192 (
            .O(N__46383),
            .I(N__46372));
    InMux I__11191 (
            .O(N__46382),
            .I(N__46369));
    Span4Mux_v I__11190 (
            .O(N__46379),
            .I(N__46366));
    Span4Mux_h I__11189 (
            .O(N__46372),
            .I(N__46363));
    LocalMux I__11188 (
            .O(N__46369),
            .I(data_out_frame2_9_0));
    Odrv4 I__11187 (
            .O(N__46366),
            .I(data_out_frame2_9_0));
    Odrv4 I__11186 (
            .O(N__46363),
            .I(data_out_frame2_9_0));
    CascadeMux I__11185 (
            .O(N__46356),
            .I(\c0.n18891_cascade_ ));
    InMux I__11184 (
            .O(N__46353),
            .I(N__46349));
    InMux I__11183 (
            .O(N__46352),
            .I(N__46346));
    LocalMux I__11182 (
            .O(N__46349),
            .I(N__46342));
    LocalMux I__11181 (
            .O(N__46346),
            .I(N__46338));
    InMux I__11180 (
            .O(N__46345),
            .I(N__46335));
    Span4Mux_h I__11179 (
            .O(N__46342),
            .I(N__46332));
    InMux I__11178 (
            .O(N__46341),
            .I(N__46328));
    Span4Mux_h I__11177 (
            .O(N__46338),
            .I(N__46325));
    LocalMux I__11176 (
            .O(N__46335),
            .I(N__46320));
    Span4Mux_v I__11175 (
            .O(N__46332),
            .I(N__46320));
    InMux I__11174 (
            .O(N__46331),
            .I(N__46317));
    LocalMux I__11173 (
            .O(N__46328),
            .I(data_out_frame2_8_0));
    Odrv4 I__11172 (
            .O(N__46325),
            .I(data_out_frame2_8_0));
    Odrv4 I__11171 (
            .O(N__46320),
            .I(data_out_frame2_8_0));
    LocalMux I__11170 (
            .O(N__46317),
            .I(data_out_frame2_8_0));
    InMux I__11169 (
            .O(N__46308),
            .I(N__46305));
    LocalMux I__11168 (
            .O(N__46305),
            .I(N__46300));
    InMux I__11167 (
            .O(N__46304),
            .I(N__46297));
    InMux I__11166 (
            .O(N__46303),
            .I(N__46294));
    Span4Mux_s2_v I__11165 (
            .O(N__46300),
            .I(N__46291));
    LocalMux I__11164 (
            .O(N__46297),
            .I(N__46288));
    LocalMux I__11163 (
            .O(N__46294),
            .I(N__46284));
    Span4Mux_v I__11162 (
            .O(N__46291),
            .I(N__46279));
    Span4Mux_h I__11161 (
            .O(N__46288),
            .I(N__46279));
    InMux I__11160 (
            .O(N__46287),
            .I(N__46276));
    Span12Mux_s9_v I__11159 (
            .O(N__46284),
            .I(N__46273));
    Span4Mux_h I__11158 (
            .O(N__46279),
            .I(N__46270));
    LocalMux I__11157 (
            .O(N__46276),
            .I(data_out_frame2_14_0));
    Odrv12 I__11156 (
            .O(N__46273),
            .I(data_out_frame2_14_0));
    Odrv4 I__11155 (
            .O(N__46270),
            .I(data_out_frame2_14_0));
    CascadeMux I__11154 (
            .O(N__46263),
            .I(N__46258));
    InMux I__11153 (
            .O(N__46262),
            .I(N__46255));
    InMux I__11152 (
            .O(N__46261),
            .I(N__46252));
    InMux I__11151 (
            .O(N__46258),
            .I(N__46249));
    LocalMux I__11150 (
            .O(N__46255),
            .I(N__46246));
    LocalMux I__11149 (
            .O(N__46252),
            .I(N__46243));
    LocalMux I__11148 (
            .O(N__46249),
            .I(N__46240));
    IoSpan4Mux I__11147 (
            .O(N__46246),
            .I(N__46235));
    Span4Mux_v I__11146 (
            .O(N__46243),
            .I(N__46235));
    Span4Mux_h I__11145 (
            .O(N__46240),
            .I(N__46230));
    Span4Mux_s0_v I__11144 (
            .O(N__46235),
            .I(N__46227));
    InMux I__11143 (
            .O(N__46234),
            .I(N__46222));
    InMux I__11142 (
            .O(N__46233),
            .I(N__46222));
    Span4Mux_v I__11141 (
            .O(N__46230),
            .I(N__46219));
    Odrv4 I__11140 (
            .O(N__46227),
            .I(data_out_frame2_15_0));
    LocalMux I__11139 (
            .O(N__46222),
            .I(data_out_frame2_15_0));
    Odrv4 I__11138 (
            .O(N__46219),
            .I(data_out_frame2_15_0));
    CascadeMux I__11137 (
            .O(N__46212),
            .I(N__46207));
    CascadeMux I__11136 (
            .O(N__46211),
            .I(N__46202));
    CascadeMux I__11135 (
            .O(N__46210),
            .I(N__46198));
    InMux I__11134 (
            .O(N__46207),
            .I(N__46181));
    InMux I__11133 (
            .O(N__46206),
            .I(N__46170));
    InMux I__11132 (
            .O(N__46205),
            .I(N__46170));
    InMux I__11131 (
            .O(N__46202),
            .I(N__46170));
    InMux I__11130 (
            .O(N__46201),
            .I(N__46170));
    InMux I__11129 (
            .O(N__46198),
            .I(N__46170));
    InMux I__11128 (
            .O(N__46197),
            .I(N__46167));
    InMux I__11127 (
            .O(N__46196),
            .I(N__46152));
    InMux I__11126 (
            .O(N__46195),
            .I(N__46152));
    InMux I__11125 (
            .O(N__46194),
            .I(N__46145));
    InMux I__11124 (
            .O(N__46193),
            .I(N__46145));
    InMux I__11123 (
            .O(N__46192),
            .I(N__46140));
    InMux I__11122 (
            .O(N__46191),
            .I(N__46140));
    InMux I__11121 (
            .O(N__46190),
            .I(N__46136));
    InMux I__11120 (
            .O(N__46189),
            .I(N__46127));
    InMux I__11119 (
            .O(N__46188),
            .I(N__46127));
    InMux I__11118 (
            .O(N__46187),
            .I(N__46127));
    InMux I__11117 (
            .O(N__46186),
            .I(N__46127));
    InMux I__11116 (
            .O(N__46185),
            .I(N__46124));
    InMux I__11115 (
            .O(N__46184),
            .I(N__46113));
    LocalMux I__11114 (
            .O(N__46181),
            .I(N__46106));
    LocalMux I__11113 (
            .O(N__46170),
            .I(N__46106));
    LocalMux I__11112 (
            .O(N__46167),
            .I(N__46106));
    InMux I__11111 (
            .O(N__46166),
            .I(N__46101));
    InMux I__11110 (
            .O(N__46165),
            .I(N__46101));
    InMux I__11109 (
            .O(N__46164),
            .I(N__46096));
    InMux I__11108 (
            .O(N__46163),
            .I(N__46096));
    InMux I__11107 (
            .O(N__46162),
            .I(N__46093));
    InMux I__11106 (
            .O(N__46161),
            .I(N__46085));
    InMux I__11105 (
            .O(N__46160),
            .I(N__46082));
    InMux I__11104 (
            .O(N__46159),
            .I(N__46077));
    InMux I__11103 (
            .O(N__46158),
            .I(N__46072));
    InMux I__11102 (
            .O(N__46157),
            .I(N__46072));
    LocalMux I__11101 (
            .O(N__46152),
            .I(N__46069));
    InMux I__11100 (
            .O(N__46151),
            .I(N__46066));
    InMux I__11099 (
            .O(N__46150),
            .I(N__46061));
    LocalMux I__11098 (
            .O(N__46145),
            .I(N__46056));
    LocalMux I__11097 (
            .O(N__46140),
            .I(N__46056));
    InMux I__11096 (
            .O(N__46139),
            .I(N__46053));
    LocalMux I__11095 (
            .O(N__46136),
            .I(N__46046));
    LocalMux I__11094 (
            .O(N__46127),
            .I(N__46046));
    LocalMux I__11093 (
            .O(N__46124),
            .I(N__46046));
    InMux I__11092 (
            .O(N__46123),
            .I(N__46039));
    InMux I__11091 (
            .O(N__46122),
            .I(N__46039));
    InMux I__11090 (
            .O(N__46121),
            .I(N__46039));
    InMux I__11089 (
            .O(N__46120),
            .I(N__46034));
    InMux I__11088 (
            .O(N__46119),
            .I(N__46034));
    InMux I__11087 (
            .O(N__46118),
            .I(N__46027));
    InMux I__11086 (
            .O(N__46117),
            .I(N__46027));
    InMux I__11085 (
            .O(N__46116),
            .I(N__46027));
    LocalMux I__11084 (
            .O(N__46113),
            .I(N__46018));
    Span4Mux_h I__11083 (
            .O(N__46106),
            .I(N__46018));
    LocalMux I__11082 (
            .O(N__46101),
            .I(N__46018));
    LocalMux I__11081 (
            .O(N__46096),
            .I(N__46018));
    LocalMux I__11080 (
            .O(N__46093),
            .I(N__46014));
    InMux I__11079 (
            .O(N__46092),
            .I(N__46007));
    InMux I__11078 (
            .O(N__46091),
            .I(N__46007));
    InMux I__11077 (
            .O(N__46090),
            .I(N__46007));
    InMux I__11076 (
            .O(N__46089),
            .I(N__46002));
    InMux I__11075 (
            .O(N__46088),
            .I(N__46002));
    LocalMux I__11074 (
            .O(N__46085),
            .I(N__45999));
    LocalMux I__11073 (
            .O(N__46082),
            .I(N__45996));
    InMux I__11072 (
            .O(N__46081),
            .I(N__45993));
    InMux I__11071 (
            .O(N__46080),
            .I(N__45990));
    LocalMux I__11070 (
            .O(N__46077),
            .I(N__45987));
    LocalMux I__11069 (
            .O(N__46072),
            .I(N__45982));
    Span4Mux_v I__11068 (
            .O(N__46069),
            .I(N__45982));
    LocalMux I__11067 (
            .O(N__46066),
            .I(N__45979));
    InMux I__11066 (
            .O(N__46065),
            .I(N__45976));
    InMux I__11065 (
            .O(N__46064),
            .I(N__45973));
    LocalMux I__11064 (
            .O(N__46061),
            .I(N__45968));
    Span4Mux_v I__11063 (
            .O(N__46056),
            .I(N__45968));
    LocalMux I__11062 (
            .O(N__46053),
            .I(N__45963));
    Span4Mux_v I__11061 (
            .O(N__46046),
            .I(N__45963));
    LocalMux I__11060 (
            .O(N__46039),
            .I(N__45956));
    LocalMux I__11059 (
            .O(N__46034),
            .I(N__45956));
    LocalMux I__11058 (
            .O(N__46027),
            .I(N__45956));
    Span4Mux_h I__11057 (
            .O(N__46018),
            .I(N__45953));
    InMux I__11056 (
            .O(N__46017),
            .I(N__45949));
    Span4Mux_s1_v I__11055 (
            .O(N__46014),
            .I(N__45944));
    LocalMux I__11054 (
            .O(N__46007),
            .I(N__45944));
    LocalMux I__11053 (
            .O(N__46002),
            .I(N__45939));
    Span4Mux_v I__11052 (
            .O(N__45999),
            .I(N__45939));
    Span4Mux_v I__11051 (
            .O(N__45996),
            .I(N__45936));
    LocalMux I__11050 (
            .O(N__45993),
            .I(N__45933));
    LocalMux I__11049 (
            .O(N__45990),
            .I(N__45926));
    Span4Mux_v I__11048 (
            .O(N__45987),
            .I(N__45926));
    Span4Mux_v I__11047 (
            .O(N__45982),
            .I(N__45926));
    Span4Mux_h I__11046 (
            .O(N__45979),
            .I(N__45921));
    LocalMux I__11045 (
            .O(N__45976),
            .I(N__45921));
    LocalMux I__11044 (
            .O(N__45973),
            .I(N__45916));
    Span4Mux_v I__11043 (
            .O(N__45968),
            .I(N__45916));
    Span4Mux_v I__11042 (
            .O(N__45963),
            .I(N__45913));
    Span4Mux_v I__11041 (
            .O(N__45956),
            .I(N__45908));
    Span4Mux_v I__11040 (
            .O(N__45953),
            .I(N__45908));
    InMux I__11039 (
            .O(N__45952),
            .I(N__45905));
    LocalMux I__11038 (
            .O(N__45949),
            .I(N__45902));
    Span4Mux_v I__11037 (
            .O(N__45944),
            .I(N__45899));
    Span4Mux_h I__11036 (
            .O(N__45939),
            .I(N__45896));
    Span4Mux_v I__11035 (
            .O(N__45936),
            .I(N__45889));
    Span4Mux_v I__11034 (
            .O(N__45933),
            .I(N__45889));
    Span4Mux_h I__11033 (
            .O(N__45926),
            .I(N__45889));
    Span4Mux_h I__11032 (
            .O(N__45921),
            .I(N__45886));
    Span4Mux_h I__11031 (
            .O(N__45916),
            .I(N__45881));
    Span4Mux_h I__11030 (
            .O(N__45913),
            .I(N__45881));
    Span4Mux_h I__11029 (
            .O(N__45908),
            .I(N__45878));
    LocalMux I__11028 (
            .O(N__45905),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__11027 (
            .O(N__45902),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11026 (
            .O(N__45899),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11025 (
            .O(N__45896),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11024 (
            .O(N__45889),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11023 (
            .O(N__45886),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11022 (
            .O(N__45881),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__11021 (
            .O(N__45878),
            .I(\c0.byte_transmit_counter2_0 ));
    CascadeMux I__11020 (
            .O(N__45861),
            .I(N__45858));
    InMux I__11019 (
            .O(N__45858),
            .I(N__45853));
    InMux I__11018 (
            .O(N__45857),
            .I(N__45850));
    InMux I__11017 (
            .O(N__45856),
            .I(N__45846));
    LocalMux I__11016 (
            .O(N__45853),
            .I(N__45843));
    LocalMux I__11015 (
            .O(N__45850),
            .I(N__45840));
    InMux I__11014 (
            .O(N__45849),
            .I(N__45837));
    LocalMux I__11013 (
            .O(N__45846),
            .I(N__45834));
    Span4Mux_h I__11012 (
            .O(N__45843),
            .I(N__45831));
    Span4Mux_v I__11011 (
            .O(N__45840),
            .I(N__45828));
    LocalMux I__11010 (
            .O(N__45837),
            .I(data_out_frame2_13_0));
    Odrv4 I__11009 (
            .O(N__45834),
            .I(data_out_frame2_13_0));
    Odrv4 I__11008 (
            .O(N__45831),
            .I(data_out_frame2_13_0));
    Odrv4 I__11007 (
            .O(N__45828),
            .I(data_out_frame2_13_0));
    CascadeMux I__11006 (
            .O(N__45819),
            .I(\c0.n18897_cascade_ ));
    InMux I__11005 (
            .O(N__45816),
            .I(N__45811));
    InMux I__11004 (
            .O(N__45815),
            .I(N__45808));
    InMux I__11003 (
            .O(N__45814),
            .I(N__45805));
    LocalMux I__11002 (
            .O(N__45811),
            .I(N__45802));
    LocalMux I__11001 (
            .O(N__45808),
            .I(N__45798));
    LocalMux I__11000 (
            .O(N__45805),
            .I(N__45795));
    Span4Mux_v I__10999 (
            .O(N__45802),
            .I(N__45792));
    CascadeMux I__10998 (
            .O(N__45801),
            .I(N__45786));
    Span4Mux_s3_v I__10997 (
            .O(N__45798),
            .I(N__45781));
    Span4Mux_s3_v I__10996 (
            .O(N__45795),
            .I(N__45781));
    Span4Mux_v I__10995 (
            .O(N__45792),
            .I(N__45778));
    InMux I__10994 (
            .O(N__45791),
            .I(N__45773));
    InMux I__10993 (
            .O(N__45790),
            .I(N__45773));
    InMux I__10992 (
            .O(N__45789),
            .I(N__45770));
    InMux I__10991 (
            .O(N__45786),
            .I(N__45767));
    Span4Mux_h I__10990 (
            .O(N__45781),
            .I(N__45763));
    Span4Mux_s1_v I__10989 (
            .O(N__45778),
            .I(N__45758));
    LocalMux I__10988 (
            .O(N__45773),
            .I(N__45758));
    LocalMux I__10987 (
            .O(N__45770),
            .I(N__45755));
    LocalMux I__10986 (
            .O(N__45767),
            .I(N__45752));
    InMux I__10985 (
            .O(N__45766),
            .I(N__45749));
    Sp12to4 I__10984 (
            .O(N__45763),
            .I(N__45746));
    Span4Mux_h I__10983 (
            .O(N__45758),
            .I(N__45739));
    Span4Mux_h I__10982 (
            .O(N__45755),
            .I(N__45739));
    Span4Mux_h I__10981 (
            .O(N__45752),
            .I(N__45739));
    LocalMux I__10980 (
            .O(N__45749),
            .I(data_out_frame2_12_0));
    Odrv12 I__10979 (
            .O(N__45746),
            .I(data_out_frame2_12_0));
    Odrv4 I__10978 (
            .O(N__45739),
            .I(data_out_frame2_12_0));
    InMux I__10977 (
            .O(N__45732),
            .I(N__45729));
    LocalMux I__10976 (
            .O(N__45729),
            .I(\c0.n18060 ));
    CascadeMux I__10975 (
            .O(N__45726),
            .I(\c0.n18057_cascade_ ));
    InMux I__10974 (
            .O(N__45723),
            .I(N__45720));
    LocalMux I__10973 (
            .O(N__45720),
            .I(N__45717));
    Odrv12 I__10972 (
            .O(N__45717),
            .I(\c0.n18374 ));
    CascadeMux I__10971 (
            .O(N__45714),
            .I(\c0.n18723_cascade_ ));
    InMux I__10970 (
            .O(N__45711),
            .I(N__45708));
    LocalMux I__10969 (
            .O(N__45708),
            .I(N__45705));
    Span4Mux_v I__10968 (
            .O(N__45705),
            .I(N__45702));
    Span4Mux_h I__10967 (
            .O(N__45702),
            .I(N__45699));
    Odrv4 I__10966 (
            .O(N__45699),
            .I(\c0.n6_adj_2275 ));
    InMux I__10965 (
            .O(N__45696),
            .I(N__45692));
    InMux I__10964 (
            .O(N__45695),
            .I(N__45689));
    LocalMux I__10963 (
            .O(N__45692),
            .I(N__45684));
    LocalMux I__10962 (
            .O(N__45689),
            .I(N__45684));
    Span4Mux_s3_v I__10961 (
            .O(N__45684),
            .I(N__45679));
    InMux I__10960 (
            .O(N__45683),
            .I(N__45674));
    InMux I__10959 (
            .O(N__45682),
            .I(N__45674));
    Odrv4 I__10958 (
            .O(N__45679),
            .I(\c0.n17810 ));
    LocalMux I__10957 (
            .O(N__45674),
            .I(\c0.n17810 ));
    InMux I__10956 (
            .O(N__45669),
            .I(N__45664));
    InMux I__10955 (
            .O(N__45668),
            .I(N__45659));
    InMux I__10954 (
            .O(N__45667),
            .I(N__45659));
    LocalMux I__10953 (
            .O(N__45664),
            .I(N__45656));
    LocalMux I__10952 (
            .O(N__45659),
            .I(N__45651));
    Span4Mux_h I__10951 (
            .O(N__45656),
            .I(N__45647));
    InMux I__10950 (
            .O(N__45655),
            .I(N__45642));
    InMux I__10949 (
            .O(N__45654),
            .I(N__45642));
    Span4Mux_h I__10948 (
            .O(N__45651),
            .I(N__45639));
    InMux I__10947 (
            .O(N__45650),
            .I(N__45636));
    Odrv4 I__10946 (
            .O(N__45647),
            .I(data_out_frame2_11_2));
    LocalMux I__10945 (
            .O(N__45642),
            .I(data_out_frame2_11_2));
    Odrv4 I__10944 (
            .O(N__45639),
            .I(data_out_frame2_11_2));
    LocalMux I__10943 (
            .O(N__45636),
            .I(data_out_frame2_11_2));
    InMux I__10942 (
            .O(N__45627),
            .I(N__45622));
    CascadeMux I__10941 (
            .O(N__45626),
            .I(N__45618));
    InMux I__10940 (
            .O(N__45625),
            .I(N__45615));
    LocalMux I__10939 (
            .O(N__45622),
            .I(N__45610));
    InMux I__10938 (
            .O(N__45621),
            .I(N__45605));
    InMux I__10937 (
            .O(N__45618),
            .I(N__45605));
    LocalMux I__10936 (
            .O(N__45615),
            .I(N__45602));
    InMux I__10935 (
            .O(N__45614),
            .I(N__45599));
    InMux I__10934 (
            .O(N__45613),
            .I(N__45596));
    Span4Mux_s1_v I__10933 (
            .O(N__45610),
            .I(N__45593));
    LocalMux I__10932 (
            .O(N__45605),
            .I(N__45590));
    Span4Mux_h I__10931 (
            .O(N__45602),
            .I(N__45587));
    LocalMux I__10930 (
            .O(N__45599),
            .I(data_out_frame2_11_3));
    LocalMux I__10929 (
            .O(N__45596),
            .I(data_out_frame2_11_3));
    Odrv4 I__10928 (
            .O(N__45593),
            .I(data_out_frame2_11_3));
    Odrv12 I__10927 (
            .O(N__45590),
            .I(data_out_frame2_11_3));
    Odrv4 I__10926 (
            .O(N__45587),
            .I(data_out_frame2_11_3));
    InMux I__10925 (
            .O(N__45576),
            .I(N__45571));
    InMux I__10924 (
            .O(N__45575),
            .I(N__45567));
    InMux I__10923 (
            .O(N__45574),
            .I(N__45564));
    LocalMux I__10922 (
            .O(N__45571),
            .I(N__45561));
    InMux I__10921 (
            .O(N__45570),
            .I(N__45558));
    LocalMux I__10920 (
            .O(N__45567),
            .I(N__45555));
    LocalMux I__10919 (
            .O(N__45564),
            .I(data_out_frame2_11_1));
    Odrv12 I__10918 (
            .O(N__45561),
            .I(data_out_frame2_11_1));
    LocalMux I__10917 (
            .O(N__45558),
            .I(data_out_frame2_11_1));
    Odrv4 I__10916 (
            .O(N__45555),
            .I(data_out_frame2_11_1));
    InMux I__10915 (
            .O(N__45546),
            .I(N__45543));
    LocalMux I__10914 (
            .O(N__45543),
            .I(\c0.n17798 ));
    InMux I__10913 (
            .O(N__45540),
            .I(N__45537));
    LocalMux I__10912 (
            .O(N__45537),
            .I(N__45533));
    InMux I__10911 (
            .O(N__45536),
            .I(N__45530));
    Span4Mux_v I__10910 (
            .O(N__45533),
            .I(N__45527));
    LocalMux I__10909 (
            .O(N__45530),
            .I(N__45524));
    Span4Mux_h I__10908 (
            .O(N__45527),
            .I(N__45520));
    Span4Mux_s1_v I__10907 (
            .O(N__45524),
            .I(N__45517));
    InMux I__10906 (
            .O(N__45523),
            .I(N__45514));
    Odrv4 I__10905 (
            .O(N__45520),
            .I(\c0.n17751 ));
    Odrv4 I__10904 (
            .O(N__45517),
            .I(\c0.n17751 ));
    LocalMux I__10903 (
            .O(N__45514),
            .I(\c0.n17751 ));
    InMux I__10902 (
            .O(N__45507),
            .I(N__45503));
    InMux I__10901 (
            .O(N__45506),
            .I(N__45500));
    LocalMux I__10900 (
            .O(N__45503),
            .I(N__45497));
    LocalMux I__10899 (
            .O(N__45500),
            .I(N__45494));
    Odrv4 I__10898 (
            .O(N__45497),
            .I(\c0.n17868 ));
    Odrv12 I__10897 (
            .O(N__45494),
            .I(\c0.n17868 ));
    CascadeMux I__10896 (
            .O(N__45489),
            .I(\c0.n17798_cascade_ ));
    InMux I__10895 (
            .O(N__45486),
            .I(N__45483));
    LocalMux I__10894 (
            .O(N__45483),
            .I(N__45479));
    InMux I__10893 (
            .O(N__45482),
            .I(N__45476));
    Span4Mux_h I__10892 (
            .O(N__45479),
            .I(N__45473));
    LocalMux I__10891 (
            .O(N__45476),
            .I(\c0.n17902 ));
    Odrv4 I__10890 (
            .O(N__45473),
            .I(\c0.n17902 ));
    InMux I__10889 (
            .O(N__45468),
            .I(N__45465));
    LocalMux I__10888 (
            .O(N__45465),
            .I(\c0.n18_adj_2393 ));
    InMux I__10887 (
            .O(N__45462),
            .I(N__45459));
    LocalMux I__10886 (
            .O(N__45459),
            .I(N__45456));
    Span4Mux_v I__10885 (
            .O(N__45456),
            .I(N__45451));
    InMux I__10884 (
            .O(N__45455),
            .I(N__45448));
    InMux I__10883 (
            .O(N__45454),
            .I(N__45445));
    Span4Mux_h I__10882 (
            .O(N__45451),
            .I(N__45439));
    LocalMux I__10881 (
            .O(N__45448),
            .I(N__45439));
    LocalMux I__10880 (
            .O(N__45445),
            .I(N__45436));
    InMux I__10879 (
            .O(N__45444),
            .I(N__45432));
    Span4Mux_s1_v I__10878 (
            .O(N__45439),
            .I(N__45427));
    Span4Mux_h I__10877 (
            .O(N__45436),
            .I(N__45427));
    InMux I__10876 (
            .O(N__45435),
            .I(N__45424));
    LocalMux I__10875 (
            .O(N__45432),
            .I(data_out_frame2_16_5));
    Odrv4 I__10874 (
            .O(N__45427),
            .I(data_out_frame2_16_5));
    LocalMux I__10873 (
            .O(N__45424),
            .I(data_out_frame2_16_5));
    CascadeMux I__10872 (
            .O(N__45417),
            .I(\c0.n24_adj_2394_cascade_ ));
    InMux I__10871 (
            .O(N__45414),
            .I(N__45411));
    LocalMux I__10870 (
            .O(N__45411),
            .I(N__45407));
    InMux I__10869 (
            .O(N__45410),
            .I(N__45404));
    Span4Mux_v I__10868 (
            .O(N__45407),
            .I(N__45398));
    LocalMux I__10867 (
            .O(N__45404),
            .I(N__45398));
    CascadeMux I__10866 (
            .O(N__45403),
            .I(N__45395));
    Span4Mux_h I__10865 (
            .O(N__45398),
            .I(N__45391));
    InMux I__10864 (
            .O(N__45395),
            .I(N__45386));
    InMux I__10863 (
            .O(N__45394),
            .I(N__45386));
    Odrv4 I__10862 (
            .O(N__45391),
            .I(data_out_frame2_15_5));
    LocalMux I__10861 (
            .O(N__45386),
            .I(data_out_frame2_15_5));
    InMux I__10860 (
            .O(N__45381),
            .I(N__45375));
    InMux I__10859 (
            .O(N__45380),
            .I(N__45375));
    LocalMux I__10858 (
            .O(N__45375),
            .I(N__45372));
    Odrv4 I__10857 (
            .O(N__45372),
            .I(\c0.n17920 ));
    InMux I__10856 (
            .O(N__45369),
            .I(N__45366));
    LocalMux I__10855 (
            .O(N__45366),
            .I(N__45363));
    Odrv12 I__10854 (
            .O(N__45363),
            .I(\c0.n22_adj_2395 ));
    CascadeMux I__10853 (
            .O(N__45360),
            .I(\c0.n26_adj_2396_cascade_ ));
    InMux I__10852 (
            .O(N__45357),
            .I(N__45354));
    LocalMux I__10851 (
            .O(N__45354),
            .I(N__45350));
    InMux I__10850 (
            .O(N__45353),
            .I(N__45347));
    Span4Mux_h I__10849 (
            .O(N__45350),
            .I(N__45344));
    LocalMux I__10848 (
            .O(N__45347),
            .I(N__45339));
    Span4Mux_h I__10847 (
            .O(N__45344),
            .I(N__45339));
    Odrv4 I__10846 (
            .O(N__45339),
            .I(\c0.n17917 ));
    CascadeMux I__10845 (
            .O(N__45336),
            .I(N__45333));
    InMux I__10844 (
            .O(N__45333),
            .I(N__45330));
    LocalMux I__10843 (
            .O(N__45330),
            .I(N__45327));
    Span4Mux_h I__10842 (
            .O(N__45327),
            .I(N__45324));
    Span4Mux_h I__10841 (
            .O(N__45324),
            .I(N__45321));
    Sp12to4 I__10840 (
            .O(N__45321),
            .I(N__45318));
    Odrv12 I__10839 (
            .O(N__45318),
            .I(\c0.data_out_frame2_20_7 ));
    InMux I__10838 (
            .O(N__45315),
            .I(N__45312));
    LocalMux I__10837 (
            .O(N__45312),
            .I(N__45309));
    Span4Mux_v I__10836 (
            .O(N__45309),
            .I(N__45306));
    Span4Mux_v I__10835 (
            .O(N__45306),
            .I(N__45302));
    InMux I__10834 (
            .O(N__45305),
            .I(N__45299));
    Sp12to4 I__10833 (
            .O(N__45302),
            .I(N__45296));
    LocalMux I__10832 (
            .O(N__45299),
            .I(N__45293));
    Odrv12 I__10831 (
            .O(N__45296),
            .I(\c0.n10778 ));
    Odrv4 I__10830 (
            .O(N__45293),
            .I(\c0.n10778 ));
    InMux I__10829 (
            .O(N__45288),
            .I(N__45284));
    InMux I__10828 (
            .O(N__45287),
            .I(N__45281));
    LocalMux I__10827 (
            .O(N__45284),
            .I(N__45278));
    LocalMux I__10826 (
            .O(N__45281),
            .I(N__45275));
    Odrv4 I__10825 (
            .O(N__45278),
            .I(\c0.n17871 ));
    Odrv4 I__10824 (
            .O(N__45275),
            .I(\c0.n17871 ));
    CascadeMux I__10823 (
            .O(N__45270),
            .I(\c0.n14_adj_2406_cascade_ ));
    InMux I__10822 (
            .O(N__45267),
            .I(N__45264));
    LocalMux I__10821 (
            .O(N__45264),
            .I(N__45260));
    InMux I__10820 (
            .O(N__45263),
            .I(N__45257));
    Span4Mux_s1_v I__10819 (
            .O(N__45260),
            .I(N__45254));
    LocalMux I__10818 (
            .O(N__45257),
            .I(\c0.n10583 ));
    Odrv4 I__10817 (
            .O(N__45254),
            .I(\c0.n10583 ));
    InMux I__10816 (
            .O(N__45249),
            .I(N__45245));
    InMux I__10815 (
            .O(N__45248),
            .I(N__45241));
    LocalMux I__10814 (
            .O(N__45245),
            .I(N__45238));
    InMux I__10813 (
            .O(N__45244),
            .I(N__45235));
    LocalMux I__10812 (
            .O(N__45241),
            .I(N__45230));
    Span4Mux_v I__10811 (
            .O(N__45238),
            .I(N__45225));
    LocalMux I__10810 (
            .O(N__45235),
            .I(N__45225));
    InMux I__10809 (
            .O(N__45234),
            .I(N__45222));
    InMux I__10808 (
            .O(N__45233),
            .I(N__45219));
    Span4Mux_h I__10807 (
            .O(N__45230),
            .I(N__45214));
    Span4Mux_h I__10806 (
            .O(N__45225),
            .I(N__45214));
    LocalMux I__10805 (
            .O(N__45222),
            .I(data_out_frame2_11_5));
    LocalMux I__10804 (
            .O(N__45219),
            .I(data_out_frame2_11_5));
    Odrv4 I__10803 (
            .O(N__45214),
            .I(data_out_frame2_11_5));
    CascadeMux I__10802 (
            .O(N__45207),
            .I(N__45203));
    InMux I__10801 (
            .O(N__45206),
            .I(N__45198));
    InMux I__10800 (
            .O(N__45203),
            .I(N__45195));
    InMux I__10799 (
            .O(N__45202),
            .I(N__45192));
    InMux I__10798 (
            .O(N__45201),
            .I(N__45189));
    LocalMux I__10797 (
            .O(N__45198),
            .I(N__45186));
    LocalMux I__10796 (
            .O(N__45195),
            .I(N__45182));
    LocalMux I__10795 (
            .O(N__45192),
            .I(N__45179));
    LocalMux I__10794 (
            .O(N__45189),
            .I(N__45176));
    Span4Mux_h I__10793 (
            .O(N__45186),
            .I(N__45173));
    InMux I__10792 (
            .O(N__45185),
            .I(N__45170));
    Span4Mux_h I__10791 (
            .O(N__45182),
            .I(N__45167));
    Span12Mux_s11_h I__10790 (
            .O(N__45179),
            .I(N__45164));
    Span4Mux_h I__10789 (
            .O(N__45176),
            .I(N__45161));
    Span4Mux_v I__10788 (
            .O(N__45173),
            .I(N__45158));
    LocalMux I__10787 (
            .O(N__45170),
            .I(data_out_frame2_12_4));
    Odrv4 I__10786 (
            .O(N__45167),
            .I(data_out_frame2_12_4));
    Odrv12 I__10785 (
            .O(N__45164),
            .I(data_out_frame2_12_4));
    Odrv4 I__10784 (
            .O(N__45161),
            .I(data_out_frame2_12_4));
    Odrv4 I__10783 (
            .O(N__45158),
            .I(data_out_frame2_12_4));
    InMux I__10782 (
            .O(N__45147),
            .I(N__45143));
    InMux I__10781 (
            .O(N__45146),
            .I(N__45140));
    LocalMux I__10780 (
            .O(N__45143),
            .I(N__45137));
    LocalMux I__10779 (
            .O(N__45140),
            .I(N__45134));
    Span4Mux_h I__10778 (
            .O(N__45137),
            .I(N__45131));
    Span4Mux_s3_v I__10777 (
            .O(N__45134),
            .I(N__45128));
    Odrv4 I__10776 (
            .O(N__45131),
            .I(\c0.n17780 ));
    Odrv4 I__10775 (
            .O(N__45128),
            .I(\c0.n17780 ));
    InMux I__10774 (
            .O(N__45123),
            .I(N__45120));
    LocalMux I__10773 (
            .O(N__45120),
            .I(\c0.n15_adj_2407 ));
    InMux I__10772 (
            .O(N__45117),
            .I(N__45108));
    InMux I__10771 (
            .O(N__45116),
            .I(N__45108));
    InMux I__10770 (
            .O(N__45115),
            .I(N__45108));
    LocalMux I__10769 (
            .O(N__45108),
            .I(N__45104));
    InMux I__10768 (
            .O(N__45107),
            .I(N__45101));
    Span4Mux_s3_v I__10767 (
            .O(N__45104),
            .I(N__45098));
    LocalMux I__10766 (
            .O(N__45101),
            .I(data_out_frame2_7_3));
    Odrv4 I__10765 (
            .O(N__45098),
            .I(data_out_frame2_7_3));
    InMux I__10764 (
            .O(N__45093),
            .I(N__45089));
    CascadeMux I__10763 (
            .O(N__45092),
            .I(N__45085));
    LocalMux I__10762 (
            .O(N__45089),
            .I(N__45082));
    InMux I__10761 (
            .O(N__45088),
            .I(N__45079));
    InMux I__10760 (
            .O(N__45085),
            .I(N__45074));
    Span4Mux_v I__10759 (
            .O(N__45082),
            .I(N__45071));
    LocalMux I__10758 (
            .O(N__45079),
            .I(N__45068));
    InMux I__10757 (
            .O(N__45078),
            .I(N__45065));
    InMux I__10756 (
            .O(N__45077),
            .I(N__45062));
    LocalMux I__10755 (
            .O(N__45074),
            .I(N__45055));
    Span4Mux_h I__10754 (
            .O(N__45071),
            .I(N__45055));
    Span4Mux_v I__10753 (
            .O(N__45068),
            .I(N__45055));
    LocalMux I__10752 (
            .O(N__45065),
            .I(N__45052));
    LocalMux I__10751 (
            .O(N__45062),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__10750 (
            .O(N__45055),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv12 I__10749 (
            .O(N__45052),
            .I(\c0.data_out_frame2_0_3 ));
    InMux I__10748 (
            .O(N__45045),
            .I(N__45042));
    LocalMux I__10747 (
            .O(N__45042),
            .I(N__45036));
    InMux I__10746 (
            .O(N__45041),
            .I(N__45033));
    InMux I__10745 (
            .O(N__45040),
            .I(N__45030));
    InMux I__10744 (
            .O(N__45039),
            .I(N__45027));
    Span4Mux_h I__10743 (
            .O(N__45036),
            .I(N__45022));
    LocalMux I__10742 (
            .O(N__45033),
            .I(N__45022));
    LocalMux I__10741 (
            .O(N__45030),
            .I(data_out_frame2_14_3));
    LocalMux I__10740 (
            .O(N__45027),
            .I(data_out_frame2_14_3));
    Odrv4 I__10739 (
            .O(N__45022),
            .I(data_out_frame2_14_3));
    InMux I__10738 (
            .O(N__45015),
            .I(N__45010));
    InMux I__10737 (
            .O(N__45014),
            .I(N__45007));
    InMux I__10736 (
            .O(N__45013),
            .I(N__45004));
    LocalMux I__10735 (
            .O(N__45010),
            .I(N__44998));
    LocalMux I__10734 (
            .O(N__45007),
            .I(N__44998));
    LocalMux I__10733 (
            .O(N__45004),
            .I(N__44995));
    InMux I__10732 (
            .O(N__45003),
            .I(N__44991));
    Span4Mux_h I__10731 (
            .O(N__44998),
            .I(N__44988));
    Span4Mux_h I__10730 (
            .O(N__44995),
            .I(N__44985));
    InMux I__10729 (
            .O(N__44994),
            .I(N__44982));
    LocalMux I__10728 (
            .O(N__44991),
            .I(data_out_frame2_15_4));
    Odrv4 I__10727 (
            .O(N__44988),
            .I(data_out_frame2_15_4));
    Odrv4 I__10726 (
            .O(N__44985),
            .I(data_out_frame2_15_4));
    LocalMux I__10725 (
            .O(N__44982),
            .I(data_out_frame2_15_4));
    InMux I__10724 (
            .O(N__44973),
            .I(N__44968));
    CascadeMux I__10723 (
            .O(N__44972),
            .I(N__44964));
    CascadeMux I__10722 (
            .O(N__44971),
            .I(N__44961));
    LocalMux I__10721 (
            .O(N__44968),
            .I(N__44958));
    InMux I__10720 (
            .O(N__44967),
            .I(N__44953));
    InMux I__10719 (
            .O(N__44964),
            .I(N__44953));
    InMux I__10718 (
            .O(N__44961),
            .I(N__44950));
    Span4Mux_s3_v I__10717 (
            .O(N__44958),
            .I(N__44944));
    LocalMux I__10716 (
            .O(N__44953),
            .I(N__44944));
    LocalMux I__10715 (
            .O(N__44950),
            .I(N__44941));
    InMux I__10714 (
            .O(N__44949),
            .I(N__44938));
    Span4Mux_v I__10713 (
            .O(N__44944),
            .I(N__44933));
    Span4Mux_h I__10712 (
            .O(N__44941),
            .I(N__44933));
    LocalMux I__10711 (
            .O(N__44938),
            .I(data_out_frame2_7_4));
    Odrv4 I__10710 (
            .O(N__44933),
            .I(data_out_frame2_7_4));
    InMux I__10709 (
            .O(N__44928),
            .I(N__44925));
    LocalMux I__10708 (
            .O(N__44925),
            .I(\c0.n10710 ));
    CascadeMux I__10707 (
            .O(N__44922),
            .I(\c0.n10710_cascade_ ));
    InMux I__10706 (
            .O(N__44919),
            .I(N__44916));
    LocalMux I__10705 (
            .O(N__44916),
            .I(\c0.n18_adj_2402 ));
    InMux I__10704 (
            .O(N__44913),
            .I(N__44910));
    LocalMux I__10703 (
            .O(N__44910),
            .I(N__44907));
    Span4Mux_s3_v I__10702 (
            .O(N__44907),
            .I(N__44904));
    Odrv4 I__10701 (
            .O(N__44904),
            .I(\c0.n20_adj_2404 ));
    InMux I__10700 (
            .O(N__44901),
            .I(N__44895));
    InMux I__10699 (
            .O(N__44900),
            .I(N__44892));
    InMux I__10698 (
            .O(N__44899),
            .I(N__44889));
    InMux I__10697 (
            .O(N__44898),
            .I(N__44885));
    LocalMux I__10696 (
            .O(N__44895),
            .I(N__44880));
    LocalMux I__10695 (
            .O(N__44892),
            .I(N__44880));
    LocalMux I__10694 (
            .O(N__44889),
            .I(N__44877));
    InMux I__10693 (
            .O(N__44888),
            .I(N__44874));
    LocalMux I__10692 (
            .O(N__44885),
            .I(N__44871));
    Span4Mux_h I__10691 (
            .O(N__44880),
            .I(N__44866));
    Span4Mux_s3_v I__10690 (
            .O(N__44877),
            .I(N__44866));
    LocalMux I__10689 (
            .O(N__44874),
            .I(data_out_frame2_6_5));
    Odrv4 I__10688 (
            .O(N__44871),
            .I(data_out_frame2_6_5));
    Odrv4 I__10687 (
            .O(N__44866),
            .I(data_out_frame2_6_5));
    InMux I__10686 (
            .O(N__44859),
            .I(N__44854));
    InMux I__10685 (
            .O(N__44858),
            .I(N__44847));
    InMux I__10684 (
            .O(N__44857),
            .I(N__44847));
    LocalMux I__10683 (
            .O(N__44854),
            .I(N__44844));
    InMux I__10682 (
            .O(N__44853),
            .I(N__44841));
    InMux I__10681 (
            .O(N__44852),
            .I(N__44838));
    LocalMux I__10680 (
            .O(N__44847),
            .I(N__44835));
    Span4Mux_h I__10679 (
            .O(N__44844),
            .I(N__44832));
    LocalMux I__10678 (
            .O(N__44841),
            .I(N__44829));
    LocalMux I__10677 (
            .O(N__44838),
            .I(data_out_frame2_7_5));
    Odrv12 I__10676 (
            .O(N__44835),
            .I(data_out_frame2_7_5));
    Odrv4 I__10675 (
            .O(N__44832),
            .I(data_out_frame2_7_5));
    Odrv4 I__10674 (
            .O(N__44829),
            .I(data_out_frame2_7_5));
    InMux I__10673 (
            .O(N__44820),
            .I(N__44817));
    LocalMux I__10672 (
            .O(N__44817),
            .I(N__44814));
    Odrv12 I__10671 (
            .O(N__44814),
            .I(\c0.n5_adj_2386 ));
    InMux I__10670 (
            .O(N__44811),
            .I(N__44807));
    InMux I__10669 (
            .O(N__44810),
            .I(N__44802));
    LocalMux I__10668 (
            .O(N__44807),
            .I(N__44799));
    InMux I__10667 (
            .O(N__44806),
            .I(N__44796));
    CascadeMux I__10666 (
            .O(N__44805),
            .I(N__44793));
    LocalMux I__10665 (
            .O(N__44802),
            .I(N__44789));
    Span4Mux_v I__10664 (
            .O(N__44799),
            .I(N__44786));
    LocalMux I__10663 (
            .O(N__44796),
            .I(N__44783));
    InMux I__10662 (
            .O(N__44793),
            .I(N__44780));
    InMux I__10661 (
            .O(N__44792),
            .I(N__44777));
    Span4Mux_h I__10660 (
            .O(N__44789),
            .I(N__44774));
    Span4Mux_h I__10659 (
            .O(N__44786),
            .I(N__44771));
    Span4Mux_h I__10658 (
            .O(N__44783),
            .I(N__44768));
    LocalMux I__10657 (
            .O(N__44780),
            .I(N__44765));
    LocalMux I__10656 (
            .O(N__44777),
            .I(data_out_frame2_13_5));
    Odrv4 I__10655 (
            .O(N__44774),
            .I(data_out_frame2_13_5));
    Odrv4 I__10654 (
            .O(N__44771),
            .I(data_out_frame2_13_5));
    Odrv4 I__10653 (
            .O(N__44768),
            .I(data_out_frame2_13_5));
    Odrv4 I__10652 (
            .O(N__44765),
            .I(data_out_frame2_13_5));
    InMux I__10651 (
            .O(N__44754),
            .I(N__44750));
    InMux I__10650 (
            .O(N__44753),
            .I(N__44746));
    LocalMux I__10649 (
            .O(N__44750),
            .I(N__44743));
    InMux I__10648 (
            .O(N__44749),
            .I(N__44738));
    LocalMux I__10647 (
            .O(N__44746),
            .I(N__44735));
    Span4Mux_h I__10646 (
            .O(N__44743),
            .I(N__44732));
    InMux I__10645 (
            .O(N__44742),
            .I(N__44727));
    InMux I__10644 (
            .O(N__44741),
            .I(N__44727));
    LocalMux I__10643 (
            .O(N__44738),
            .I(data_out_frame2_10_7));
    Odrv12 I__10642 (
            .O(N__44735),
            .I(data_out_frame2_10_7));
    Odrv4 I__10641 (
            .O(N__44732),
            .I(data_out_frame2_10_7));
    LocalMux I__10640 (
            .O(N__44727),
            .I(data_out_frame2_10_7));
    InMux I__10639 (
            .O(N__44718),
            .I(N__44715));
    LocalMux I__10638 (
            .O(N__44715),
            .I(\c0.n10877 ));
    CascadeMux I__10637 (
            .O(N__44712),
            .I(\c0.n10593_cascade_ ));
    InMux I__10636 (
            .O(N__44709),
            .I(N__44706));
    LocalMux I__10635 (
            .O(N__44706),
            .I(N__44703));
    Span4Mux_h I__10634 (
            .O(N__44703),
            .I(N__44700));
    Odrv4 I__10633 (
            .O(N__44700),
            .I(\c0.n14 ));
    InMux I__10632 (
            .O(N__44697),
            .I(N__44691));
    InMux I__10631 (
            .O(N__44696),
            .I(N__44691));
    LocalMux I__10630 (
            .O(N__44691),
            .I(N__44687));
    InMux I__10629 (
            .O(N__44690),
            .I(N__44684));
    Span4Mux_v I__10628 (
            .O(N__44687),
            .I(N__44678));
    LocalMux I__10627 (
            .O(N__44684),
            .I(N__44678));
    InMux I__10626 (
            .O(N__44683),
            .I(N__44674));
    Span4Mux_h I__10625 (
            .O(N__44678),
            .I(N__44671));
    InMux I__10624 (
            .O(N__44677),
            .I(N__44668));
    LocalMux I__10623 (
            .O(N__44674),
            .I(data_out_frame2_7_6));
    Odrv4 I__10622 (
            .O(N__44671),
            .I(data_out_frame2_7_6));
    LocalMux I__10621 (
            .O(N__44668),
            .I(data_out_frame2_7_6));
    InMux I__10620 (
            .O(N__44661),
            .I(N__44656));
    InMux I__10619 (
            .O(N__44660),
            .I(N__44653));
    InMux I__10618 (
            .O(N__44659),
            .I(N__44650));
    LocalMux I__10617 (
            .O(N__44656),
            .I(N__44646));
    LocalMux I__10616 (
            .O(N__44653),
            .I(N__44641));
    LocalMux I__10615 (
            .O(N__44650),
            .I(N__44641));
    InMux I__10614 (
            .O(N__44649),
            .I(N__44638));
    Span4Mux_h I__10613 (
            .O(N__44646),
            .I(N__44635));
    Span4Mux_s3_v I__10612 (
            .O(N__44641),
            .I(N__44632));
    LocalMux I__10611 (
            .O(N__44638),
            .I(data_out_frame2_5_7));
    Odrv4 I__10610 (
            .O(N__44635),
            .I(data_out_frame2_5_7));
    Odrv4 I__10609 (
            .O(N__44632),
            .I(data_out_frame2_5_7));
    CascadeMux I__10608 (
            .O(N__44625),
            .I(N__44621));
    InMux I__10607 (
            .O(N__44624),
            .I(N__44618));
    InMux I__10606 (
            .O(N__44621),
            .I(N__44615));
    LocalMux I__10605 (
            .O(N__44618),
            .I(N__44610));
    LocalMux I__10604 (
            .O(N__44615),
            .I(N__44607));
    InMux I__10603 (
            .O(N__44614),
            .I(N__44604));
    InMux I__10602 (
            .O(N__44613),
            .I(N__44601));
    Span4Mux_h I__10601 (
            .O(N__44610),
            .I(N__44594));
    Span4Mux_v I__10600 (
            .O(N__44607),
            .I(N__44594));
    LocalMux I__10599 (
            .O(N__44604),
            .I(N__44594));
    LocalMux I__10598 (
            .O(N__44601),
            .I(data_out_frame2_9_5));
    Odrv4 I__10597 (
            .O(N__44594),
            .I(data_out_frame2_9_5));
    CascadeMux I__10596 (
            .O(N__44589),
            .I(N__44586));
    InMux I__10595 (
            .O(N__44586),
            .I(N__44583));
    LocalMux I__10594 (
            .O(N__44583),
            .I(N__44578));
    InMux I__10593 (
            .O(N__44582),
            .I(N__44575));
    CascadeMux I__10592 (
            .O(N__44581),
            .I(N__44572));
    Span4Mux_s1_v I__10591 (
            .O(N__44578),
            .I(N__44568));
    LocalMux I__10590 (
            .O(N__44575),
            .I(N__44565));
    InMux I__10589 (
            .O(N__44572),
            .I(N__44561));
    InMux I__10588 (
            .O(N__44571),
            .I(N__44558));
    Span4Mux_v I__10587 (
            .O(N__44568),
            .I(N__44555));
    Span4Mux_s3_v I__10586 (
            .O(N__44565),
            .I(N__44552));
    InMux I__10585 (
            .O(N__44564),
            .I(N__44549));
    LocalMux I__10584 (
            .O(N__44561),
            .I(N__44546));
    LocalMux I__10583 (
            .O(N__44558),
            .I(data_out_frame2_9_3));
    Odrv4 I__10582 (
            .O(N__44555),
            .I(data_out_frame2_9_3));
    Odrv4 I__10581 (
            .O(N__44552),
            .I(data_out_frame2_9_3));
    LocalMux I__10580 (
            .O(N__44549),
            .I(data_out_frame2_9_3));
    Odrv12 I__10579 (
            .O(N__44546),
            .I(data_out_frame2_9_3));
    CascadeMux I__10578 (
            .O(N__44535),
            .I(N__44532));
    InMux I__10577 (
            .O(N__44532),
            .I(N__44529));
    LocalMux I__10576 (
            .O(N__44529),
            .I(\c0.n10929 ));
    CascadeMux I__10575 (
            .O(N__44526),
            .I(\c0.n10929_cascade_ ));
    InMux I__10574 (
            .O(N__44523),
            .I(N__44520));
    LocalMux I__10573 (
            .O(N__44520),
            .I(\c0.n17823 ));
    InMux I__10572 (
            .O(N__44517),
            .I(N__44514));
    LocalMux I__10571 (
            .O(N__44514),
            .I(N__44510));
    InMux I__10570 (
            .O(N__44513),
            .I(N__44507));
    Odrv12 I__10569 (
            .O(N__44510),
            .I(\c0.n17853 ));
    LocalMux I__10568 (
            .O(N__44507),
            .I(\c0.n17853 ));
    CascadeMux I__10567 (
            .O(N__44502),
            .I(\c0.n17823_cascade_ ));
    InMux I__10566 (
            .O(N__44499),
            .I(N__44496));
    LocalMux I__10565 (
            .O(N__44496),
            .I(\c0.n17895 ));
    CascadeMux I__10564 (
            .O(N__44493),
            .I(\c0.n17_adj_2401_cascade_ ));
    InMux I__10563 (
            .O(N__44490),
            .I(N__44486));
    InMux I__10562 (
            .O(N__44489),
            .I(N__44483));
    LocalMux I__10561 (
            .O(N__44486),
            .I(N__44480));
    LocalMux I__10560 (
            .O(N__44483),
            .I(N__44477));
    Span4Mux_v I__10559 (
            .O(N__44480),
            .I(N__44474));
    Odrv4 I__10558 (
            .O(N__44477),
            .I(\c0.n17914 ));
    Odrv4 I__10557 (
            .O(N__44474),
            .I(\c0.n17914 ));
    InMux I__10556 (
            .O(N__44469),
            .I(N__44466));
    LocalMux I__10555 (
            .O(N__44466),
            .I(N__44463));
    Span4Mux_v I__10554 (
            .O(N__44463),
            .I(N__44460));
    Odrv4 I__10553 (
            .O(N__44460),
            .I(\c0.data_out_frame2_20_6 ));
    InMux I__10552 (
            .O(N__44457),
            .I(N__44454));
    LocalMux I__10551 (
            .O(N__44454),
            .I(N__44450));
    InMux I__10550 (
            .O(N__44453),
            .I(N__44447));
    Span4Mux_h I__10549 (
            .O(N__44450),
            .I(N__44444));
    LocalMux I__10548 (
            .O(N__44447),
            .I(\c0.n10703 ));
    Odrv4 I__10547 (
            .O(N__44444),
            .I(\c0.n10703 ));
    CascadeMux I__10546 (
            .O(N__44439),
            .I(N__44434));
    CascadeMux I__10545 (
            .O(N__44438),
            .I(N__44430));
    InMux I__10544 (
            .O(N__44437),
            .I(N__44427));
    InMux I__10543 (
            .O(N__44434),
            .I(N__44424));
    InMux I__10542 (
            .O(N__44433),
            .I(N__44419));
    InMux I__10541 (
            .O(N__44430),
            .I(N__44419));
    LocalMux I__10540 (
            .O(N__44427),
            .I(N__44415));
    LocalMux I__10539 (
            .O(N__44424),
            .I(N__44412));
    LocalMux I__10538 (
            .O(N__44419),
            .I(N__44409));
    InMux I__10537 (
            .O(N__44418),
            .I(N__44406));
    Span12Mux_s5_v I__10536 (
            .O(N__44415),
            .I(N__44403));
    Span4Mux_h I__10535 (
            .O(N__44412),
            .I(N__44400));
    Span4Mux_v I__10534 (
            .O(N__44409),
            .I(N__44397));
    LocalMux I__10533 (
            .O(N__44406),
            .I(data_out_frame2_14_4));
    Odrv12 I__10532 (
            .O(N__44403),
            .I(data_out_frame2_14_4));
    Odrv4 I__10531 (
            .O(N__44400),
            .I(data_out_frame2_14_4));
    Odrv4 I__10530 (
            .O(N__44397),
            .I(data_out_frame2_14_4));
    InMux I__10529 (
            .O(N__44388),
            .I(N__44385));
    LocalMux I__10528 (
            .O(N__44385),
            .I(N__44382));
    Span4Mux_h I__10527 (
            .O(N__44382),
            .I(N__44379));
    Odrv4 I__10526 (
            .O(N__44379),
            .I(\c0.n10825 ));
    InMux I__10525 (
            .O(N__44376),
            .I(N__44371));
    InMux I__10524 (
            .O(N__44375),
            .I(N__44368));
    InMux I__10523 (
            .O(N__44374),
            .I(N__44364));
    LocalMux I__10522 (
            .O(N__44371),
            .I(N__44361));
    LocalMux I__10521 (
            .O(N__44368),
            .I(N__44358));
    CascadeMux I__10520 (
            .O(N__44367),
            .I(N__44355));
    LocalMux I__10519 (
            .O(N__44364),
            .I(N__44352));
    Span4Mux_h I__10518 (
            .O(N__44361),
            .I(N__44347));
    Span4Mux_s2_v I__10517 (
            .O(N__44358),
            .I(N__44347));
    InMux I__10516 (
            .O(N__44355),
            .I(N__44344));
    Span4Mux_h I__10515 (
            .O(N__44352),
            .I(N__44341));
    Span4Mux_h I__10514 (
            .O(N__44347),
            .I(N__44338));
    LocalMux I__10513 (
            .O(N__44344),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv4 I__10512 (
            .O(N__44341),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv4 I__10511 (
            .O(N__44338),
            .I(\c0.data_out_frame2_0_5 ));
    InMux I__10510 (
            .O(N__44331),
            .I(N__44326));
    InMux I__10509 (
            .O(N__44330),
            .I(N__44321));
    InMux I__10508 (
            .O(N__44329),
            .I(N__44318));
    LocalMux I__10507 (
            .O(N__44326),
            .I(N__44315));
    InMux I__10506 (
            .O(N__44325),
            .I(N__44310));
    InMux I__10505 (
            .O(N__44324),
            .I(N__44310));
    LocalMux I__10504 (
            .O(N__44321),
            .I(N__44304));
    LocalMux I__10503 (
            .O(N__44318),
            .I(N__44304));
    Span4Mux_v I__10502 (
            .O(N__44315),
            .I(N__44299));
    LocalMux I__10501 (
            .O(N__44310),
            .I(N__44299));
    InMux I__10500 (
            .O(N__44309),
            .I(N__44296));
    Span4Mux_v I__10499 (
            .O(N__44304),
            .I(N__44291));
    Span4Mux_h I__10498 (
            .O(N__44299),
            .I(N__44291));
    LocalMux I__10497 (
            .O(N__44296),
            .I(data_out_frame2_8_1));
    Odrv4 I__10496 (
            .O(N__44291),
            .I(data_out_frame2_8_1));
    InMux I__10495 (
            .O(N__44286),
            .I(N__44281));
    CascadeMux I__10494 (
            .O(N__44285),
            .I(N__44278));
    InMux I__10493 (
            .O(N__44284),
            .I(N__44275));
    LocalMux I__10492 (
            .O(N__44281),
            .I(N__44272));
    InMux I__10491 (
            .O(N__44278),
            .I(N__44269));
    LocalMux I__10490 (
            .O(N__44275),
            .I(N__44264));
    Span4Mux_s2_v I__10489 (
            .O(N__44272),
            .I(N__44261));
    LocalMux I__10488 (
            .O(N__44269),
            .I(N__44258));
    InMux I__10487 (
            .O(N__44268),
            .I(N__44255));
    InMux I__10486 (
            .O(N__44267),
            .I(N__44252));
    Span4Mux_s2_v I__10485 (
            .O(N__44264),
            .I(N__44249));
    Span4Mux_h I__10484 (
            .O(N__44261),
            .I(N__44244));
    Span4Mux_h I__10483 (
            .O(N__44258),
            .I(N__44244));
    LocalMux I__10482 (
            .O(N__44255),
            .I(N__44241));
    LocalMux I__10481 (
            .O(N__44252),
            .I(data_out_frame2_12_7));
    Odrv4 I__10480 (
            .O(N__44249),
            .I(data_out_frame2_12_7));
    Odrv4 I__10479 (
            .O(N__44244),
            .I(data_out_frame2_12_7));
    Odrv12 I__10478 (
            .O(N__44241),
            .I(data_out_frame2_12_7));
    InMux I__10477 (
            .O(N__44232),
            .I(N__44225));
    InMux I__10476 (
            .O(N__44231),
            .I(N__44222));
    InMux I__10475 (
            .O(N__44230),
            .I(N__44219));
    InMux I__10474 (
            .O(N__44229),
            .I(N__44216));
    CascadeMux I__10473 (
            .O(N__44228),
            .I(N__44213));
    LocalMux I__10472 (
            .O(N__44225),
            .I(N__44210));
    LocalMux I__10471 (
            .O(N__44222),
            .I(N__44207));
    LocalMux I__10470 (
            .O(N__44219),
            .I(N__44204));
    LocalMux I__10469 (
            .O(N__44216),
            .I(N__44200));
    InMux I__10468 (
            .O(N__44213),
            .I(N__44197));
    Span4Mux_v I__10467 (
            .O(N__44210),
            .I(N__44194));
    Span4Mux_h I__10466 (
            .O(N__44207),
            .I(N__44189));
    Span4Mux_h I__10465 (
            .O(N__44204),
            .I(N__44189));
    InMux I__10464 (
            .O(N__44203),
            .I(N__44186));
    Span12Mux_h I__10463 (
            .O(N__44200),
            .I(N__44181));
    LocalMux I__10462 (
            .O(N__44197),
            .I(N__44181));
    Odrv4 I__10461 (
            .O(N__44194),
            .I(rand_data_5));
    Odrv4 I__10460 (
            .O(N__44189),
            .I(rand_data_5));
    LocalMux I__10459 (
            .O(N__44186),
            .I(rand_data_5));
    Odrv12 I__10458 (
            .O(N__44181),
            .I(rand_data_5));
    CascadeMux I__10457 (
            .O(N__44172),
            .I(N__44168));
    CascadeMux I__10456 (
            .O(N__44171),
            .I(N__44164));
    InMux I__10455 (
            .O(N__44168),
            .I(N__44161));
    InMux I__10454 (
            .O(N__44167),
            .I(N__44157));
    InMux I__10453 (
            .O(N__44164),
            .I(N__44154));
    LocalMux I__10452 (
            .O(N__44161),
            .I(N__44151));
    InMux I__10451 (
            .O(N__44160),
            .I(N__44147));
    LocalMux I__10450 (
            .O(N__44157),
            .I(N__44144));
    LocalMux I__10449 (
            .O(N__44154),
            .I(N__44141));
    Span4Mux_h I__10448 (
            .O(N__44151),
            .I(N__44137));
    InMux I__10447 (
            .O(N__44150),
            .I(N__44134));
    LocalMux I__10446 (
            .O(N__44147),
            .I(N__44131));
    Span4Mux_s3_v I__10445 (
            .O(N__44144),
            .I(N__44126));
    Span4Mux_s3_v I__10444 (
            .O(N__44141),
            .I(N__44126));
    InMux I__10443 (
            .O(N__44140),
            .I(N__44123));
    Span4Mux_h I__10442 (
            .O(N__44137),
            .I(N__44120));
    LocalMux I__10441 (
            .O(N__44134),
            .I(N__44117));
    Span4Mux_s3_v I__10440 (
            .O(N__44131),
            .I(N__44112));
    Span4Mux_h I__10439 (
            .O(N__44126),
            .I(N__44112));
    LocalMux I__10438 (
            .O(N__44123),
            .I(data_out_frame2_12_5));
    Odrv4 I__10437 (
            .O(N__44120),
            .I(data_out_frame2_12_5));
    Odrv4 I__10436 (
            .O(N__44117),
            .I(data_out_frame2_12_5));
    Odrv4 I__10435 (
            .O(N__44112),
            .I(data_out_frame2_12_5));
    InMux I__10434 (
            .O(N__44103),
            .I(N__44100));
    LocalMux I__10433 (
            .O(N__44100),
            .I(N__44096));
    InMux I__10432 (
            .O(N__44099),
            .I(N__44093));
    Span4Mux_v I__10431 (
            .O(N__44096),
            .I(N__44088));
    LocalMux I__10430 (
            .O(N__44093),
            .I(N__44088));
    Span4Mux_h I__10429 (
            .O(N__44088),
            .I(N__44083));
    InMux I__10428 (
            .O(N__44087),
            .I(N__44080));
    InMux I__10427 (
            .O(N__44086),
            .I(N__44077));
    Span4Mux_v I__10426 (
            .O(N__44083),
            .I(N__44074));
    LocalMux I__10425 (
            .O(N__44080),
            .I(data_out_frame2_6_3));
    LocalMux I__10424 (
            .O(N__44077),
            .I(data_out_frame2_6_3));
    Odrv4 I__10423 (
            .O(N__44074),
            .I(data_out_frame2_6_3));
    InMux I__10422 (
            .O(N__44067),
            .I(N__44064));
    LocalMux I__10421 (
            .O(N__44064),
            .I(\c0.n5_adj_2381 ));
    CascadeMux I__10420 (
            .O(N__44061),
            .I(N__44058));
    InMux I__10419 (
            .O(N__44058),
            .I(N__44054));
    InMux I__10418 (
            .O(N__44057),
            .I(N__44050));
    LocalMux I__10417 (
            .O(N__44054),
            .I(N__44047));
    InMux I__10416 (
            .O(N__44053),
            .I(N__44044));
    LocalMux I__10415 (
            .O(N__44050),
            .I(N__44041));
    Span4Mux_v I__10414 (
            .O(N__44047),
            .I(N__44037));
    LocalMux I__10413 (
            .O(N__44044),
            .I(N__44034));
    Span4Mux_h I__10412 (
            .O(N__44041),
            .I(N__44031));
    InMux I__10411 (
            .O(N__44040),
            .I(N__44028));
    Span4Mux_h I__10410 (
            .O(N__44037),
            .I(N__44025));
    Span4Mux_v I__10409 (
            .O(N__44034),
            .I(N__44022));
    Span4Mux_h I__10408 (
            .O(N__44031),
            .I(N__44019));
    LocalMux I__10407 (
            .O(N__44028),
            .I(data_out_frame2_6_1));
    Odrv4 I__10406 (
            .O(N__44025),
            .I(data_out_frame2_6_1));
    Odrv4 I__10405 (
            .O(N__44022),
            .I(data_out_frame2_6_1));
    Odrv4 I__10404 (
            .O(N__44019),
            .I(data_out_frame2_6_1));
    InMux I__10403 (
            .O(N__44010),
            .I(N__44007));
    LocalMux I__10402 (
            .O(N__44007),
            .I(N__44004));
    Span4Mux_s2_v I__10401 (
            .O(N__44004),
            .I(N__44001));
    Odrv4 I__10400 (
            .O(N__44001),
            .I(\c0.n30_adj_2434 ));
    InMux I__10399 (
            .O(N__43998),
            .I(N__43995));
    LocalMux I__10398 (
            .O(N__43995),
            .I(\c0.data_out_frame2_20_2 ));
    CascadeMux I__10397 (
            .O(N__43992),
            .I(\c0.n18636_cascade_ ));
    InMux I__10396 (
            .O(N__43989),
            .I(N__43986));
    LocalMux I__10395 (
            .O(N__43986),
            .I(\c0.n22_adj_2268 ));
    CascadeMux I__10394 (
            .O(N__43983),
            .I(N__43980));
    InMux I__10393 (
            .O(N__43980),
            .I(N__43976));
    InMux I__10392 (
            .O(N__43979),
            .I(N__43973));
    LocalMux I__10391 (
            .O(N__43976),
            .I(N__43970));
    LocalMux I__10390 (
            .O(N__43973),
            .I(N__43967));
    Span4Mux_s2_v I__10389 (
            .O(N__43970),
            .I(N__43964));
    Odrv12 I__10388 (
            .O(N__43967),
            .I(\c0.n17892 ));
    Odrv4 I__10387 (
            .O(N__43964),
            .I(\c0.n17892 ));
    InMux I__10386 (
            .O(N__43959),
            .I(N__43955));
    CascadeMux I__10385 (
            .O(N__43958),
            .I(N__43951));
    LocalMux I__10384 (
            .O(N__43955),
            .I(N__43946));
    InMux I__10383 (
            .O(N__43954),
            .I(N__43943));
    InMux I__10382 (
            .O(N__43951),
            .I(N__43940));
    InMux I__10381 (
            .O(N__43950),
            .I(N__43937));
    InMux I__10380 (
            .O(N__43949),
            .I(N__43934));
    Span4Mux_s2_v I__10379 (
            .O(N__43946),
            .I(N__43931));
    LocalMux I__10378 (
            .O(N__43943),
            .I(N__43928));
    LocalMux I__10377 (
            .O(N__43940),
            .I(N__43925));
    LocalMux I__10376 (
            .O(N__43937),
            .I(N__43922));
    LocalMux I__10375 (
            .O(N__43934),
            .I(data_out_frame2_9_1));
    Odrv4 I__10374 (
            .O(N__43931),
            .I(data_out_frame2_9_1));
    Odrv12 I__10373 (
            .O(N__43928),
            .I(data_out_frame2_9_1));
    Odrv4 I__10372 (
            .O(N__43925),
            .I(data_out_frame2_9_1));
    Odrv4 I__10371 (
            .O(N__43922),
            .I(data_out_frame2_9_1));
    InMux I__10370 (
            .O(N__43911),
            .I(N__43908));
    LocalMux I__10369 (
            .O(N__43908),
            .I(N__43905));
    Odrv12 I__10368 (
            .O(N__43905),
            .I(\c0.n10893 ));
    CascadeMux I__10367 (
            .O(N__43902),
            .I(\c0.n20_adj_2438_cascade_ ));
    InMux I__10366 (
            .O(N__43899),
            .I(N__43896));
    LocalMux I__10365 (
            .O(N__43896),
            .I(N__43893));
    Span4Mux_h I__10364 (
            .O(N__43893),
            .I(N__43889));
    InMux I__10363 (
            .O(N__43892),
            .I(N__43886));
    Odrv4 I__10362 (
            .O(N__43889),
            .I(\c0.n17755 ));
    LocalMux I__10361 (
            .O(N__43886),
            .I(\c0.n17755 ));
    CascadeMux I__10360 (
            .O(N__43881),
            .I(N__43878));
    InMux I__10359 (
            .O(N__43878),
            .I(N__43875));
    LocalMux I__10358 (
            .O(N__43875),
            .I(N__43872));
    Span4Mux_v I__10357 (
            .O(N__43872),
            .I(N__43869));
    Odrv4 I__10356 (
            .O(N__43869),
            .I(\c0.data_out_frame2_19_6 ));
    InMux I__10355 (
            .O(N__43866),
            .I(N__43862));
    InMux I__10354 (
            .O(N__43865),
            .I(N__43859));
    LocalMux I__10353 (
            .O(N__43862),
            .I(N__43856));
    LocalMux I__10352 (
            .O(N__43859),
            .I(N__43852));
    Span4Mux_v I__10351 (
            .O(N__43856),
            .I(N__43849));
    InMux I__10350 (
            .O(N__43855),
            .I(N__43846));
    Span4Mux_v I__10349 (
            .O(N__43852),
            .I(N__43842));
    Sp12to4 I__10348 (
            .O(N__43849),
            .I(N__43837));
    LocalMux I__10347 (
            .O(N__43846),
            .I(N__43837));
    InMux I__10346 (
            .O(N__43845),
            .I(N__43834));
    Span4Mux_v I__10345 (
            .O(N__43842),
            .I(N__43831));
    Span12Mux_h I__10344 (
            .O(N__43837),
            .I(N__43828));
    LocalMux I__10343 (
            .O(N__43834),
            .I(data_out_frame2_5_3));
    Odrv4 I__10342 (
            .O(N__43831),
            .I(data_out_frame2_5_3));
    Odrv12 I__10341 (
            .O(N__43828),
            .I(data_out_frame2_5_3));
    CascadeMux I__10340 (
            .O(N__43821),
            .I(N__43815));
    InMux I__10339 (
            .O(N__43820),
            .I(N__43812));
    InMux I__10338 (
            .O(N__43819),
            .I(N__43807));
    InMux I__10337 (
            .O(N__43818),
            .I(N__43807));
    InMux I__10336 (
            .O(N__43815),
            .I(N__43804));
    LocalMux I__10335 (
            .O(N__43812),
            .I(N__43801));
    LocalMux I__10334 (
            .O(N__43807),
            .I(N__43798));
    LocalMux I__10333 (
            .O(N__43804),
            .I(N__43794));
    Span4Mux_h I__10332 (
            .O(N__43801),
            .I(N__43789));
    Span4Mux_h I__10331 (
            .O(N__43798),
            .I(N__43789));
    InMux I__10330 (
            .O(N__43797),
            .I(N__43786));
    Span4Mux_h I__10329 (
            .O(N__43794),
            .I(N__43781));
    Span4Mux_v I__10328 (
            .O(N__43789),
            .I(N__43781));
    LocalMux I__10327 (
            .O(N__43786),
            .I(data_out_frame2_12_3));
    Odrv4 I__10326 (
            .O(N__43781),
            .I(data_out_frame2_12_3));
    InMux I__10325 (
            .O(N__43776),
            .I(N__43773));
    LocalMux I__10324 (
            .O(N__43773),
            .I(\c0.n10905 ));
    CascadeMux I__10323 (
            .O(N__43770),
            .I(\c0.n10905_cascade_ ));
    InMux I__10322 (
            .O(N__43767),
            .I(N__43764));
    LocalMux I__10321 (
            .O(N__43764),
            .I(\c0.n16_adj_2391 ));
    InMux I__10320 (
            .O(N__43761),
            .I(N__43756));
    InMux I__10319 (
            .O(N__43760),
            .I(N__43753));
    InMux I__10318 (
            .O(N__43759),
            .I(N__43749));
    LocalMux I__10317 (
            .O(N__43756),
            .I(N__43746));
    LocalMux I__10316 (
            .O(N__43753),
            .I(N__43742));
    InMux I__10315 (
            .O(N__43752),
            .I(N__43739));
    LocalMux I__10314 (
            .O(N__43749),
            .I(N__43734));
    Span4Mux_v I__10313 (
            .O(N__43746),
            .I(N__43734));
    InMux I__10312 (
            .O(N__43745),
            .I(N__43731));
    Span4Mux_h I__10311 (
            .O(N__43742),
            .I(N__43726));
    LocalMux I__10310 (
            .O(N__43739),
            .I(N__43726));
    Sp12to4 I__10309 (
            .O(N__43734),
            .I(N__43723));
    LocalMux I__10308 (
            .O(N__43731),
            .I(N__43720));
    Span4Mux_v I__10307 (
            .O(N__43726),
            .I(N__43717));
    Odrv12 I__10306 (
            .O(N__43723),
            .I(data_out_frame2_8_2));
    Odrv4 I__10305 (
            .O(N__43720),
            .I(data_out_frame2_8_2));
    Odrv4 I__10304 (
            .O(N__43717),
            .I(data_out_frame2_8_2));
    InMux I__10303 (
            .O(N__43710),
            .I(N__43703));
    InMux I__10302 (
            .O(N__43709),
            .I(N__43703));
    InMux I__10301 (
            .O(N__43708),
            .I(N__43700));
    LocalMux I__10300 (
            .O(N__43703),
            .I(N__43696));
    LocalMux I__10299 (
            .O(N__43700),
            .I(N__43693));
    InMux I__10298 (
            .O(N__43699),
            .I(N__43690));
    Span4Mux_h I__10297 (
            .O(N__43696),
            .I(N__43685));
    Span4Mux_s1_v I__10296 (
            .O(N__43693),
            .I(N__43685));
    LocalMux I__10295 (
            .O(N__43690),
            .I(data_out_frame2_14_6));
    Odrv4 I__10294 (
            .O(N__43685),
            .I(data_out_frame2_14_6));
    InMux I__10293 (
            .O(N__43680),
            .I(N__43676));
    CascadeMux I__10292 (
            .O(N__43679),
            .I(N__43672));
    LocalMux I__10291 (
            .O(N__43676),
            .I(N__43669));
    InMux I__10290 (
            .O(N__43675),
            .I(N__43666));
    InMux I__10289 (
            .O(N__43672),
            .I(N__43663));
    Span4Mux_h I__10288 (
            .O(N__43669),
            .I(N__43657));
    LocalMux I__10287 (
            .O(N__43666),
            .I(N__43650));
    LocalMux I__10286 (
            .O(N__43663),
            .I(N__43650));
    InMux I__10285 (
            .O(N__43662),
            .I(N__43645));
    InMux I__10284 (
            .O(N__43661),
            .I(N__43645));
    InMux I__10283 (
            .O(N__43660),
            .I(N__43642));
    Span4Mux_h I__10282 (
            .O(N__43657),
            .I(N__43639));
    InMux I__10281 (
            .O(N__43656),
            .I(N__43636));
    InMux I__10280 (
            .O(N__43655),
            .I(N__43633));
    Span4Mux_v I__10279 (
            .O(N__43650),
            .I(N__43630));
    LocalMux I__10278 (
            .O(N__43645),
            .I(N__43627));
    LocalMux I__10277 (
            .O(N__43642),
            .I(data_out_frame2_11_7));
    Odrv4 I__10276 (
            .O(N__43639),
            .I(data_out_frame2_11_7));
    LocalMux I__10275 (
            .O(N__43636),
            .I(data_out_frame2_11_7));
    LocalMux I__10274 (
            .O(N__43633),
            .I(data_out_frame2_11_7));
    Odrv4 I__10273 (
            .O(N__43630),
            .I(data_out_frame2_11_7));
    Odrv4 I__10272 (
            .O(N__43627),
            .I(data_out_frame2_11_7));
    InMux I__10271 (
            .O(N__43614),
            .I(N__43611));
    LocalMux I__10270 (
            .O(N__43611),
            .I(N__43607));
    InMux I__10269 (
            .O(N__43610),
            .I(N__43604));
    Span4Mux_h I__10268 (
            .O(N__43607),
            .I(N__43599));
    LocalMux I__10267 (
            .O(N__43604),
            .I(N__43596));
    InMux I__10266 (
            .O(N__43603),
            .I(N__43591));
    InMux I__10265 (
            .O(N__43602),
            .I(N__43591));
    Odrv4 I__10264 (
            .O(N__43599),
            .I(data_out_frame2_14_5));
    Odrv4 I__10263 (
            .O(N__43596),
            .I(data_out_frame2_14_5));
    LocalMux I__10262 (
            .O(N__43591),
            .I(data_out_frame2_14_5));
    CascadeMux I__10261 (
            .O(N__43584),
            .I(N__43580));
    InMux I__10260 (
            .O(N__43583),
            .I(N__43576));
    InMux I__10259 (
            .O(N__43580),
            .I(N__43571));
    InMux I__10258 (
            .O(N__43579),
            .I(N__43568));
    LocalMux I__10257 (
            .O(N__43576),
            .I(N__43565));
    InMux I__10256 (
            .O(N__43575),
            .I(N__43562));
    InMux I__10255 (
            .O(N__43574),
            .I(N__43559));
    LocalMux I__10254 (
            .O(N__43571),
            .I(N__43556));
    LocalMux I__10253 (
            .O(N__43568),
            .I(data_out_frame2_12_6));
    Odrv4 I__10252 (
            .O(N__43565),
            .I(data_out_frame2_12_6));
    LocalMux I__10251 (
            .O(N__43562),
            .I(data_out_frame2_12_6));
    LocalMux I__10250 (
            .O(N__43559),
            .I(data_out_frame2_12_6));
    Odrv4 I__10249 (
            .O(N__43556),
            .I(data_out_frame2_12_6));
    InMux I__10248 (
            .O(N__43545),
            .I(N__43541));
    InMux I__10247 (
            .O(N__43544),
            .I(N__43538));
    LocalMux I__10246 (
            .O(N__43541),
            .I(rand_setpoint_31));
    LocalMux I__10245 (
            .O(N__43538),
            .I(rand_setpoint_31));
    CascadeMux I__10244 (
            .O(N__43533),
            .I(N__43530));
    InMux I__10243 (
            .O(N__43530),
            .I(N__43524));
    InMux I__10242 (
            .O(N__43529),
            .I(N__43521));
    InMux I__10241 (
            .O(N__43528),
            .I(N__43518));
    InMux I__10240 (
            .O(N__43527),
            .I(N__43515));
    LocalMux I__10239 (
            .O(N__43524),
            .I(N__43511));
    LocalMux I__10238 (
            .O(N__43521),
            .I(N__43508));
    LocalMux I__10237 (
            .O(N__43518),
            .I(N__43505));
    LocalMux I__10236 (
            .O(N__43515),
            .I(N__43502));
    InMux I__10235 (
            .O(N__43514),
            .I(N__43499));
    Span4Mux_h I__10234 (
            .O(N__43511),
            .I(N__43494));
    Span4Mux_v I__10233 (
            .O(N__43508),
            .I(N__43494));
    Span4Mux_h I__10232 (
            .O(N__43505),
            .I(N__43491));
    Span4Mux_v I__10231 (
            .O(N__43502),
            .I(N__43488));
    LocalMux I__10230 (
            .O(N__43499),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv4 I__10229 (
            .O(N__43494),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv4 I__10228 (
            .O(N__43491),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv4 I__10227 (
            .O(N__43488),
            .I(\c0.data_out_7__3__N_441 ));
    SRMux I__10226 (
            .O(N__43479),
            .I(N__43474));
    SRMux I__10225 (
            .O(N__43478),
            .I(N__43471));
    SRMux I__10224 (
            .O(N__43477),
            .I(N__43468));
    LocalMux I__10223 (
            .O(N__43474),
            .I(N__43463));
    LocalMux I__10222 (
            .O(N__43471),
            .I(N__43463));
    LocalMux I__10221 (
            .O(N__43468),
            .I(N__43459));
    Span4Mux_h I__10220 (
            .O(N__43463),
            .I(N__43456));
    SRMux I__10219 (
            .O(N__43462),
            .I(N__43453));
    Span4Mux_v I__10218 (
            .O(N__43459),
            .I(N__43450));
    Span4Mux_h I__10217 (
            .O(N__43456),
            .I(N__43447));
    LocalMux I__10216 (
            .O(N__43453),
            .I(N__43444));
    Odrv4 I__10215 (
            .O(N__43450),
            .I(\c0.n11277 ));
    Odrv4 I__10214 (
            .O(N__43447),
            .I(\c0.n11277 ));
    Odrv12 I__10213 (
            .O(N__43444),
            .I(\c0.n11277 ));
    InMux I__10212 (
            .O(N__43437),
            .I(N__43434));
    LocalMux I__10211 (
            .O(N__43434),
            .I(N__43431));
    Span4Mux_h I__10210 (
            .O(N__43431),
            .I(N__43428));
    Odrv4 I__10209 (
            .O(N__43428),
            .I(\c0.data_out_1_1 ));
    CEMux I__10208 (
            .O(N__43425),
            .I(N__43420));
    CEMux I__10207 (
            .O(N__43424),
            .I(N__43414));
    CEMux I__10206 (
            .O(N__43423),
            .I(N__43406));
    LocalMux I__10205 (
            .O(N__43420),
            .I(N__43403));
    CEMux I__10204 (
            .O(N__43419),
            .I(N__43400));
    CEMux I__10203 (
            .O(N__43418),
            .I(N__43397));
    CEMux I__10202 (
            .O(N__43417),
            .I(N__43390));
    LocalMux I__10201 (
            .O(N__43414),
            .I(N__43387));
    CEMux I__10200 (
            .O(N__43413),
            .I(N__43384));
    InMux I__10199 (
            .O(N__43412),
            .I(N__43377));
    InMux I__10198 (
            .O(N__43411),
            .I(N__43377));
    CascadeMux I__10197 (
            .O(N__43410),
            .I(N__43373));
    CascadeMux I__10196 (
            .O(N__43409),
            .I(N__43369));
    LocalMux I__10195 (
            .O(N__43406),
            .I(N__43365));
    Span4Mux_v I__10194 (
            .O(N__43403),
            .I(N__43362));
    LocalMux I__10193 (
            .O(N__43400),
            .I(N__43357));
    LocalMux I__10192 (
            .O(N__43397),
            .I(N__43357));
    CEMux I__10191 (
            .O(N__43396),
            .I(N__43354));
    InMux I__10190 (
            .O(N__43395),
            .I(N__43351));
    InMux I__10189 (
            .O(N__43394),
            .I(N__43348));
    CascadeMux I__10188 (
            .O(N__43393),
            .I(N__43343));
    LocalMux I__10187 (
            .O(N__43390),
            .I(N__43336));
    Span4Mux_v I__10186 (
            .O(N__43387),
            .I(N__43336));
    LocalMux I__10185 (
            .O(N__43384),
            .I(N__43336));
    CEMux I__10184 (
            .O(N__43383),
            .I(N__43333));
    InMux I__10183 (
            .O(N__43382),
            .I(N__43330));
    LocalMux I__10182 (
            .O(N__43377),
            .I(N__43327));
    InMux I__10181 (
            .O(N__43376),
            .I(N__43320));
    InMux I__10180 (
            .O(N__43373),
            .I(N__43320));
    InMux I__10179 (
            .O(N__43372),
            .I(N__43320));
    InMux I__10178 (
            .O(N__43369),
            .I(N__43314));
    InMux I__10177 (
            .O(N__43368),
            .I(N__43311));
    Span4Mux_v I__10176 (
            .O(N__43365),
            .I(N__43308));
    Span4Mux_v I__10175 (
            .O(N__43362),
            .I(N__43301));
    Span4Mux_v I__10174 (
            .O(N__43357),
            .I(N__43301));
    LocalMux I__10173 (
            .O(N__43354),
            .I(N__43301));
    LocalMux I__10172 (
            .O(N__43351),
            .I(N__43296));
    LocalMux I__10171 (
            .O(N__43348),
            .I(N__43296));
    InMux I__10170 (
            .O(N__43347),
            .I(N__43293));
    InMux I__10169 (
            .O(N__43346),
            .I(N__43290));
    InMux I__10168 (
            .O(N__43343),
            .I(N__43287));
    Span4Mux_h I__10167 (
            .O(N__43336),
            .I(N__43282));
    LocalMux I__10166 (
            .O(N__43333),
            .I(N__43282));
    LocalMux I__10165 (
            .O(N__43330),
            .I(N__43279));
    Span4Mux_v I__10164 (
            .O(N__43327),
            .I(N__43274));
    LocalMux I__10163 (
            .O(N__43320),
            .I(N__43274));
    InMux I__10162 (
            .O(N__43319),
            .I(N__43271));
    CascadeMux I__10161 (
            .O(N__43318),
            .I(N__43266));
    CascadeMux I__10160 (
            .O(N__43317),
            .I(N__43261));
    LocalMux I__10159 (
            .O(N__43314),
            .I(N__43254));
    LocalMux I__10158 (
            .O(N__43311),
            .I(N__43254));
    Span4Mux_h I__10157 (
            .O(N__43308),
            .I(N__43249));
    Span4Mux_h I__10156 (
            .O(N__43301),
            .I(N__43249));
    Span4Mux_h I__10155 (
            .O(N__43296),
            .I(N__43244));
    LocalMux I__10154 (
            .O(N__43293),
            .I(N__43244));
    LocalMux I__10153 (
            .O(N__43290),
            .I(N__43239));
    LocalMux I__10152 (
            .O(N__43287),
            .I(N__43239));
    Span4Mux_v I__10151 (
            .O(N__43282),
            .I(N__43230));
    Span4Mux_v I__10150 (
            .O(N__43279),
            .I(N__43230));
    Span4Mux_v I__10149 (
            .O(N__43274),
            .I(N__43230));
    LocalMux I__10148 (
            .O(N__43271),
            .I(N__43230));
    InMux I__10147 (
            .O(N__43270),
            .I(N__43227));
    InMux I__10146 (
            .O(N__43269),
            .I(N__43222));
    InMux I__10145 (
            .O(N__43266),
            .I(N__43222));
    InMux I__10144 (
            .O(N__43265),
            .I(N__43217));
    InMux I__10143 (
            .O(N__43264),
            .I(N__43217));
    InMux I__10142 (
            .O(N__43261),
            .I(N__43212));
    InMux I__10141 (
            .O(N__43260),
            .I(N__43212));
    InMux I__10140 (
            .O(N__43259),
            .I(N__43209));
    Span4Mux_h I__10139 (
            .O(N__43254),
            .I(N__43206));
    Odrv4 I__10138 (
            .O(N__43249),
            .I(n11017));
    Odrv4 I__10137 (
            .O(N__43244),
            .I(n11017));
    Odrv4 I__10136 (
            .O(N__43239),
            .I(n11017));
    Odrv4 I__10135 (
            .O(N__43230),
            .I(n11017));
    LocalMux I__10134 (
            .O(N__43227),
            .I(n11017));
    LocalMux I__10133 (
            .O(N__43222),
            .I(n11017));
    LocalMux I__10132 (
            .O(N__43217),
            .I(n11017));
    LocalMux I__10131 (
            .O(N__43212),
            .I(n11017));
    LocalMux I__10130 (
            .O(N__43209),
            .I(n11017));
    Odrv4 I__10129 (
            .O(N__43206),
            .I(n11017));
    InMux I__10128 (
            .O(N__43185),
            .I(N__43182));
    LocalMux I__10127 (
            .O(N__43182),
            .I(N__43179));
    Odrv4 I__10126 (
            .O(N__43179),
            .I(\c0.n18250 ));
    CascadeMux I__10125 (
            .O(N__43176),
            .I(N__43173));
    InMux I__10124 (
            .O(N__43173),
            .I(N__43170));
    LocalMux I__10123 (
            .O(N__43170),
            .I(N__43166));
    CascadeMux I__10122 (
            .O(N__43169),
            .I(N__43163));
    Span4Mux_v I__10121 (
            .O(N__43166),
            .I(N__43160));
    InMux I__10120 (
            .O(N__43163),
            .I(N__43157));
    Odrv4 I__10119 (
            .O(N__43160),
            .I(rand_setpoint_8));
    LocalMux I__10118 (
            .O(N__43157),
            .I(rand_setpoint_8));
    InMux I__10117 (
            .O(N__43152),
            .I(N__43149));
    LocalMux I__10116 (
            .O(N__43149),
            .I(N__43144));
    InMux I__10115 (
            .O(N__43148),
            .I(N__43141));
    InMux I__10114 (
            .O(N__43147),
            .I(N__43138));
    Span4Mux_v I__10113 (
            .O(N__43144),
            .I(N__43133));
    LocalMux I__10112 (
            .O(N__43141),
            .I(N__43133));
    LocalMux I__10111 (
            .O(N__43138),
            .I(N__43130));
    Span4Mux_h I__10110 (
            .O(N__43133),
            .I(N__43127));
    Odrv12 I__10109 (
            .O(N__43130),
            .I(\c0.data_out_7_0 ));
    Odrv4 I__10108 (
            .O(N__43127),
            .I(\c0.data_out_7_0 ));
    InMux I__10107 (
            .O(N__43122),
            .I(N__43119));
    LocalMux I__10106 (
            .O(N__43119),
            .I(N__43116));
    Odrv4 I__10105 (
            .O(N__43116),
            .I(\c0.n18648 ));
    CascadeMux I__10104 (
            .O(N__43113),
            .I(N__43110));
    InMux I__10103 (
            .O(N__43110),
            .I(N__43107));
    LocalMux I__10102 (
            .O(N__43107),
            .I(N__43104));
    Odrv12 I__10101 (
            .O(N__43104),
            .I(\c0.n18642 ));
    InMux I__10100 (
            .O(N__43101),
            .I(N__43098));
    LocalMux I__10099 (
            .O(N__43098),
            .I(N__43095));
    Span4Mux_h I__10098 (
            .O(N__43095),
            .I(N__43092));
    Odrv4 I__10097 (
            .O(N__43092),
            .I(\c0.n18221 ));
    CascadeMux I__10096 (
            .O(N__43089),
            .I(\c0.n18765_cascade_ ));
    InMux I__10095 (
            .O(N__43086),
            .I(N__43083));
    LocalMux I__10094 (
            .O(N__43083),
            .I(N__43080));
    Odrv4 I__10093 (
            .O(N__43080),
            .I(\c0.n6_adj_2227 ));
    CascadeMux I__10092 (
            .O(N__43077),
            .I(\c0.n18768_cascade_ ));
    InMux I__10091 (
            .O(N__43074),
            .I(N__43071));
    LocalMux I__10090 (
            .O(N__43071),
            .I(N__43068));
    Span4Mux_h I__10089 (
            .O(N__43068),
            .I(N__43065));
    Span4Mux_h I__10088 (
            .O(N__43065),
            .I(N__43062));
    Span4Mux_v I__10087 (
            .O(N__43062),
            .I(N__43059));
    Odrv4 I__10086 (
            .O(N__43059),
            .I(\c0.tx2.r_Tx_Data_2 ));
    InMux I__10085 (
            .O(N__43056),
            .I(N__43053));
    LocalMux I__10084 (
            .O(N__43053),
            .I(N__43049));
    InMux I__10083 (
            .O(N__43052),
            .I(N__43046));
    Span4Mux_s2_v I__10082 (
            .O(N__43049),
            .I(N__43043));
    LocalMux I__10081 (
            .O(N__43046),
            .I(data_out_frame2_18_2));
    Odrv4 I__10080 (
            .O(N__43043),
            .I(data_out_frame2_18_2));
    CascadeMux I__10079 (
            .O(N__43038),
            .I(N__43035));
    InMux I__10078 (
            .O(N__43035),
            .I(N__43032));
    LocalMux I__10077 (
            .O(N__43032),
            .I(N__43029));
    Odrv12 I__10076 (
            .O(N__43029),
            .I(\c0.data_out_frame2_19_2 ));
    InMux I__10075 (
            .O(N__43026),
            .I(N__43023));
    LocalMux I__10074 (
            .O(N__43023),
            .I(N__43020));
    Sp12to4 I__10073 (
            .O(N__43020),
            .I(N__43016));
    InMux I__10072 (
            .O(N__43019),
            .I(N__43013));
    Span12Mux_s2_v I__10071 (
            .O(N__43016),
            .I(N__43010));
    LocalMux I__10070 (
            .O(N__43013),
            .I(data_out_frame2_17_2));
    Odrv12 I__10069 (
            .O(N__43010),
            .I(data_out_frame2_17_2));
    CascadeMux I__10068 (
            .O(N__43005),
            .I(\c0.n18633_cascade_ ));
    InMux I__10067 (
            .O(N__43002),
            .I(N__42999));
    LocalMux I__10066 (
            .O(N__42999),
            .I(\c0.n18780 ));
    CascadeMux I__10065 (
            .O(N__42996),
            .I(\c0.n22_adj_2240_cascade_ ));
    InMux I__10064 (
            .O(N__42993),
            .I(N__42990));
    LocalMux I__10063 (
            .O(N__42990),
            .I(N__42987));
    Span12Mux_s5_h I__10062 (
            .O(N__42987),
            .I(N__42984));
    Odrv12 I__10061 (
            .O(N__42984),
            .I(\c0.tx2.r_Tx_Data_6 ));
    CascadeMux I__10060 (
            .O(N__42981),
            .I(\c0.n18783_cascade_ ));
    InMux I__10059 (
            .O(N__42978),
            .I(N__42973));
    InMux I__10058 (
            .O(N__42977),
            .I(N__42970));
    InMux I__10057 (
            .O(N__42976),
            .I(N__42966));
    LocalMux I__10056 (
            .O(N__42973),
            .I(N__42963));
    LocalMux I__10055 (
            .O(N__42970),
            .I(N__42960));
    InMux I__10054 (
            .O(N__42969),
            .I(N__42957));
    LocalMux I__10053 (
            .O(N__42966),
            .I(N__42952));
    Span12Mux_h I__10052 (
            .O(N__42963),
            .I(N__42952));
    Span4Mux_h I__10051 (
            .O(N__42960),
            .I(N__42949));
    LocalMux I__10050 (
            .O(N__42957),
            .I(data_out_frame2_13_4));
    Odrv12 I__10049 (
            .O(N__42952),
            .I(data_out_frame2_13_4));
    Odrv4 I__10048 (
            .O(N__42949),
            .I(data_out_frame2_13_4));
    InMux I__10047 (
            .O(N__42942),
            .I(N__42938));
    InMux I__10046 (
            .O(N__42941),
            .I(N__42934));
    LocalMux I__10045 (
            .O(N__42938),
            .I(N__42930));
    InMux I__10044 (
            .O(N__42937),
            .I(N__42926));
    LocalMux I__10043 (
            .O(N__42934),
            .I(N__42923));
    InMux I__10042 (
            .O(N__42933),
            .I(N__42920));
    Span4Mux_v I__10041 (
            .O(N__42930),
            .I(N__42917));
    InMux I__10040 (
            .O(N__42929),
            .I(N__42914));
    LocalMux I__10039 (
            .O(N__42926),
            .I(N__42911));
    Span4Mux_h I__10038 (
            .O(N__42923),
            .I(N__42906));
    LocalMux I__10037 (
            .O(N__42920),
            .I(N__42906));
    Odrv4 I__10036 (
            .O(N__42917),
            .I(\c0.data_out_7__2__N_447 ));
    LocalMux I__10035 (
            .O(N__42914),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__10034 (
            .O(N__42911),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__10033 (
            .O(N__42906),
            .I(\c0.data_out_7__2__N_447 ));
    InMux I__10032 (
            .O(N__42897),
            .I(N__42894));
    LocalMux I__10031 (
            .O(N__42894),
            .I(N__42891));
    Odrv12 I__10030 (
            .O(N__42891),
            .I(\c0.n18311 ));
    CascadeMux I__10029 (
            .O(N__42888),
            .I(N__42884));
    InMux I__10028 (
            .O(N__42887),
            .I(N__42881));
    InMux I__10027 (
            .O(N__42884),
            .I(N__42878));
    LocalMux I__10026 (
            .O(N__42881),
            .I(rand_setpoint_11));
    LocalMux I__10025 (
            .O(N__42878),
            .I(rand_setpoint_11));
    InMux I__10024 (
            .O(N__42873),
            .I(N__42852));
    InMux I__10023 (
            .O(N__42872),
            .I(N__42852));
    InMux I__10022 (
            .O(N__42871),
            .I(N__42843));
    InMux I__10021 (
            .O(N__42870),
            .I(N__42843));
    InMux I__10020 (
            .O(N__42869),
            .I(N__42843));
    InMux I__10019 (
            .O(N__42868),
            .I(N__42843));
    InMux I__10018 (
            .O(N__42867),
            .I(N__42836));
    InMux I__10017 (
            .O(N__42866),
            .I(N__42836));
    InMux I__10016 (
            .O(N__42865),
            .I(N__42836));
    InMux I__10015 (
            .O(N__42864),
            .I(N__42831));
    InMux I__10014 (
            .O(N__42863),
            .I(N__42831));
    InMux I__10013 (
            .O(N__42862),
            .I(N__42827));
    InMux I__10012 (
            .O(N__42861),
            .I(N__42824));
    InMux I__10011 (
            .O(N__42860),
            .I(N__42805));
    InMux I__10010 (
            .O(N__42859),
            .I(N__42792));
    InMux I__10009 (
            .O(N__42858),
            .I(N__42792));
    InMux I__10008 (
            .O(N__42857),
            .I(N__42789));
    LocalMux I__10007 (
            .O(N__42852),
            .I(N__42782));
    LocalMux I__10006 (
            .O(N__42843),
            .I(N__42782));
    LocalMux I__10005 (
            .O(N__42836),
            .I(N__42782));
    LocalMux I__10004 (
            .O(N__42831),
            .I(N__42776));
    InMux I__10003 (
            .O(N__42830),
            .I(N__42773));
    LocalMux I__10002 (
            .O(N__42827),
            .I(N__42770));
    LocalMux I__10001 (
            .O(N__42824),
            .I(N__42767));
    InMux I__10000 (
            .O(N__42823),
            .I(N__42758));
    InMux I__9999 (
            .O(N__42822),
            .I(N__42758));
    InMux I__9998 (
            .O(N__42821),
            .I(N__42758));
    InMux I__9997 (
            .O(N__42820),
            .I(N__42758));
    InMux I__9996 (
            .O(N__42819),
            .I(N__42749));
    InMux I__9995 (
            .O(N__42818),
            .I(N__42749));
    InMux I__9994 (
            .O(N__42817),
            .I(N__42749));
    InMux I__9993 (
            .O(N__42816),
            .I(N__42749));
    InMux I__9992 (
            .O(N__42815),
            .I(N__42742));
    InMux I__9991 (
            .O(N__42814),
            .I(N__42742));
    InMux I__9990 (
            .O(N__42813),
            .I(N__42742));
    InMux I__9989 (
            .O(N__42812),
            .I(N__42739));
    InMux I__9988 (
            .O(N__42811),
            .I(N__42736));
    InMux I__9987 (
            .O(N__42810),
            .I(N__42731));
    InMux I__9986 (
            .O(N__42809),
            .I(N__42731));
    InMux I__9985 (
            .O(N__42808),
            .I(N__42728));
    LocalMux I__9984 (
            .O(N__42805),
            .I(N__42725));
    InMux I__9983 (
            .O(N__42804),
            .I(N__42718));
    InMux I__9982 (
            .O(N__42803),
            .I(N__42718));
    InMux I__9981 (
            .O(N__42802),
            .I(N__42718));
    InMux I__9980 (
            .O(N__42801),
            .I(N__42713));
    InMux I__9979 (
            .O(N__42800),
            .I(N__42713));
    CascadeMux I__9978 (
            .O(N__42799),
            .I(N__42709));
    InMux I__9977 (
            .O(N__42798),
            .I(N__42704));
    InMux I__9976 (
            .O(N__42797),
            .I(N__42701));
    LocalMux I__9975 (
            .O(N__42792),
            .I(N__42694));
    LocalMux I__9974 (
            .O(N__42789),
            .I(N__42694));
    Span4Mux_v I__9973 (
            .O(N__42782),
            .I(N__42694));
    InMux I__9972 (
            .O(N__42781),
            .I(N__42691));
    InMux I__9971 (
            .O(N__42780),
            .I(N__42686));
    InMux I__9970 (
            .O(N__42779),
            .I(N__42686));
    Span4Mux_v I__9969 (
            .O(N__42776),
            .I(N__42683));
    LocalMux I__9968 (
            .O(N__42773),
            .I(N__42670));
    Span4Mux_h I__9967 (
            .O(N__42770),
            .I(N__42670));
    Span4Mux_v I__9966 (
            .O(N__42767),
            .I(N__42670));
    LocalMux I__9965 (
            .O(N__42758),
            .I(N__42670));
    LocalMux I__9964 (
            .O(N__42749),
            .I(N__42670));
    LocalMux I__9963 (
            .O(N__42742),
            .I(N__42670));
    LocalMux I__9962 (
            .O(N__42739),
            .I(N__42655));
    LocalMux I__9961 (
            .O(N__42736),
            .I(N__42655));
    LocalMux I__9960 (
            .O(N__42731),
            .I(N__42655));
    LocalMux I__9959 (
            .O(N__42728),
            .I(N__42655));
    Span4Mux_v I__9958 (
            .O(N__42725),
            .I(N__42655));
    LocalMux I__9957 (
            .O(N__42718),
            .I(N__42655));
    LocalMux I__9956 (
            .O(N__42713),
            .I(N__42655));
    InMux I__9955 (
            .O(N__42712),
            .I(N__42652));
    InMux I__9954 (
            .O(N__42709),
            .I(N__42649));
    InMux I__9953 (
            .O(N__42708),
            .I(N__42646));
    InMux I__9952 (
            .O(N__42707),
            .I(N__42643));
    LocalMux I__9951 (
            .O(N__42704),
            .I(N__42636));
    LocalMux I__9950 (
            .O(N__42701),
            .I(N__42636));
    Span4Mux_v I__9949 (
            .O(N__42694),
            .I(N__42636));
    LocalMux I__9948 (
            .O(N__42691),
            .I(N__42627));
    LocalMux I__9947 (
            .O(N__42686),
            .I(N__42627));
    Span4Mux_h I__9946 (
            .O(N__42683),
            .I(N__42627));
    Span4Mux_v I__9945 (
            .O(N__42670),
            .I(N__42627));
    Sp12to4 I__9944 (
            .O(N__42655),
            .I(N__42622));
    LocalMux I__9943 (
            .O(N__42652),
            .I(N__42622));
    LocalMux I__9942 (
            .O(N__42649),
            .I(N__42619));
    LocalMux I__9941 (
            .O(N__42646),
            .I(byte_transmit_counter_0));
    LocalMux I__9940 (
            .O(N__42643),
            .I(byte_transmit_counter_0));
    Odrv4 I__9939 (
            .O(N__42636),
            .I(byte_transmit_counter_0));
    Odrv4 I__9938 (
            .O(N__42627),
            .I(byte_transmit_counter_0));
    Odrv12 I__9937 (
            .O(N__42622),
            .I(byte_transmit_counter_0));
    Odrv4 I__9936 (
            .O(N__42619),
            .I(byte_transmit_counter_0));
    InMux I__9935 (
            .O(N__42606),
            .I(N__42601));
    InMux I__9934 (
            .O(N__42605),
            .I(N__42597));
    InMux I__9933 (
            .O(N__42604),
            .I(N__42594));
    LocalMux I__9932 (
            .O(N__42601),
            .I(N__42591));
    InMux I__9931 (
            .O(N__42600),
            .I(N__42588));
    LocalMux I__9930 (
            .O(N__42597),
            .I(N__42585));
    LocalMux I__9929 (
            .O(N__42594),
            .I(N__42582));
    Span4Mux_h I__9928 (
            .O(N__42591),
            .I(N__42577));
    LocalMux I__9927 (
            .O(N__42588),
            .I(N__42577));
    Span4Mux_h I__9926 (
            .O(N__42585),
            .I(N__42574));
    Span4Mux_h I__9925 (
            .O(N__42582),
            .I(N__42571));
    Span4Mux_v I__9924 (
            .O(N__42577),
            .I(N__42568));
    Odrv4 I__9923 (
            .O(N__42574),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__9922 (
            .O(N__42571),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__9921 (
            .O(N__42568),
            .I(\c0.data_out_6_3 ));
    CascadeMux I__9920 (
            .O(N__42561),
            .I(N__42558));
    InMux I__9919 (
            .O(N__42558),
            .I(N__42555));
    LocalMux I__9918 (
            .O(N__42555),
            .I(N__42552));
    Odrv12 I__9917 (
            .O(N__42552),
            .I(\c0.n5_adj_2217 ));
    CascadeMux I__9916 (
            .O(N__42549),
            .I(N__42546));
    InMux I__9915 (
            .O(N__42546),
            .I(N__42543));
    LocalMux I__9914 (
            .O(N__42543),
            .I(\c0.n18201 ));
    InMux I__9913 (
            .O(N__42540),
            .I(N__42537));
    LocalMux I__9912 (
            .O(N__42537),
            .I(N__42533));
    InMux I__9911 (
            .O(N__42536),
            .I(N__42530));
    Span4Mux_v I__9910 (
            .O(N__42533),
            .I(N__42525));
    LocalMux I__9909 (
            .O(N__42530),
            .I(N__42525));
    Span4Mux_h I__9908 (
            .O(N__42525),
            .I(N__42521));
    InMux I__9907 (
            .O(N__42524),
            .I(N__42518));
    Odrv4 I__9906 (
            .O(N__42521),
            .I(\c0.data_out_7_3 ));
    LocalMux I__9905 (
            .O(N__42518),
            .I(\c0.data_out_7_3 ));
    CascadeMux I__9904 (
            .O(N__42513),
            .I(N__42509));
    InMux I__9903 (
            .O(N__42512),
            .I(N__42506));
    InMux I__9902 (
            .O(N__42509),
            .I(N__42503));
    LocalMux I__9901 (
            .O(N__42506),
            .I(rand_setpoint_24));
    LocalMux I__9900 (
            .O(N__42503),
            .I(rand_setpoint_24));
    InMux I__9899 (
            .O(N__42498),
            .I(N__42495));
    LocalMux I__9898 (
            .O(N__42495),
            .I(N__42490));
    InMux I__9897 (
            .O(N__42494),
            .I(N__42486));
    InMux I__9896 (
            .O(N__42493),
            .I(N__42482));
    Span4Mux_v I__9895 (
            .O(N__42490),
            .I(N__42479));
    InMux I__9894 (
            .O(N__42489),
            .I(N__42476));
    LocalMux I__9893 (
            .O(N__42486),
            .I(N__42473));
    InMux I__9892 (
            .O(N__42485),
            .I(N__42470));
    LocalMux I__9891 (
            .O(N__42482),
            .I(N__42466));
    Span4Mux_h I__9890 (
            .O(N__42479),
            .I(N__42461));
    LocalMux I__9889 (
            .O(N__42476),
            .I(N__42461));
    Sp12to4 I__9888 (
            .O(N__42473),
            .I(N__42456));
    LocalMux I__9887 (
            .O(N__42470),
            .I(N__42456));
    InMux I__9886 (
            .O(N__42469),
            .I(N__42453));
    Span4Mux_h I__9885 (
            .O(N__42466),
            .I(N__42448));
    Span4Mux_h I__9884 (
            .O(N__42461),
            .I(N__42448));
    Span12Mux_v I__9883 (
            .O(N__42456),
            .I(N__42443));
    LocalMux I__9882 (
            .O(N__42453),
            .I(N__42443));
    Odrv4 I__9881 (
            .O(N__42448),
            .I(\c0.data_out_6__1__N_537 ));
    Odrv12 I__9880 (
            .O(N__42443),
            .I(\c0.data_out_6__1__N_537 ));
    InMux I__9879 (
            .O(N__42438),
            .I(N__42435));
    LocalMux I__9878 (
            .O(N__42435),
            .I(N__42432));
    Odrv12 I__9877 (
            .O(N__42432),
            .I(\c0.n18666 ));
    CascadeMux I__9876 (
            .O(N__42429),
            .I(N__42426));
    InMux I__9875 (
            .O(N__42426),
            .I(N__42423));
    LocalMux I__9874 (
            .O(N__42423),
            .I(N__42420));
    Odrv4 I__9873 (
            .O(N__42420),
            .I(\c0.n18660 ));
    InMux I__9872 (
            .O(N__42417),
            .I(N__42414));
    LocalMux I__9871 (
            .O(N__42414),
            .I(N__42411));
    Odrv12 I__9870 (
            .O(N__42411),
            .I(\c0.n18371 ));
    CascadeMux I__9869 (
            .O(N__42408),
            .I(\c0.n18735_cascade_ ));
    InMux I__9868 (
            .O(N__42405),
            .I(N__42402));
    LocalMux I__9867 (
            .O(N__42402),
            .I(N__42399));
    Odrv4 I__9866 (
            .O(N__42399),
            .I(\c0.n6_adj_2360 ));
    InMux I__9865 (
            .O(N__42396),
            .I(N__42393));
    LocalMux I__9864 (
            .O(N__42393),
            .I(\c0.n22_adj_2259 ));
    CascadeMux I__9863 (
            .O(N__42390),
            .I(\c0.n18738_cascade_ ));
    InMux I__9862 (
            .O(N__42387),
            .I(N__42384));
    LocalMux I__9861 (
            .O(N__42384),
            .I(N__42381));
    Span4Mux_h I__9860 (
            .O(N__42381),
            .I(N__42378));
    Span4Mux_h I__9859 (
            .O(N__42378),
            .I(N__42375));
    Odrv4 I__9858 (
            .O(N__42375),
            .I(\c0.tx2.r_Tx_Data_3 ));
    InMux I__9857 (
            .O(N__42372),
            .I(N__42369));
    LocalMux I__9856 (
            .O(N__42369),
            .I(N__42365));
    InMux I__9855 (
            .O(N__42368),
            .I(N__42362));
    Span4Mux_h I__9854 (
            .O(N__42365),
            .I(N__42359));
    LocalMux I__9853 (
            .O(N__42362),
            .I(data_out_frame2_18_6));
    Odrv4 I__9852 (
            .O(N__42359),
            .I(data_out_frame2_18_6));
    InMux I__9851 (
            .O(N__42354),
            .I(N__42351));
    LocalMux I__9850 (
            .O(N__42351),
            .I(N__42348));
    Odrv4 I__9849 (
            .O(N__42348),
            .I(\c0.n18708 ));
    CascadeMux I__9848 (
            .O(N__42345),
            .I(N__42342));
    InMux I__9847 (
            .O(N__42342),
            .I(N__42339));
    LocalMux I__9846 (
            .O(N__42339),
            .I(N__42336));
    Span4Mux_h I__9845 (
            .O(N__42336),
            .I(N__42333));
    Span4Mux_v I__9844 (
            .O(N__42333),
            .I(N__42330));
    Odrv4 I__9843 (
            .O(N__42330),
            .I(\c0.n18762 ));
    InMux I__9842 (
            .O(N__42327),
            .I(N__42324));
    LocalMux I__9841 (
            .O(N__42324),
            .I(N__42321));
    Span4Mux_h I__9840 (
            .O(N__42321),
            .I(N__42318));
    Odrv4 I__9839 (
            .O(N__42318),
            .I(\c0.n18308 ));
    CascadeMux I__9838 (
            .O(N__42315),
            .I(\c0.n18777_cascade_ ));
    InMux I__9837 (
            .O(N__42312),
            .I(N__42309));
    LocalMux I__9836 (
            .O(N__42309),
            .I(N__42306));
    Odrv12 I__9835 (
            .O(N__42306),
            .I(\c0.n6_adj_2218 ));
    InMux I__9834 (
            .O(N__42303),
            .I(N__42300));
    LocalMux I__9833 (
            .O(N__42300),
            .I(\c0.n18699 ));
    CascadeMux I__9832 (
            .O(N__42297),
            .I(N__42294));
    InMux I__9831 (
            .O(N__42294),
            .I(N__42291));
    LocalMux I__9830 (
            .O(N__42291),
            .I(N__42287));
    InMux I__9829 (
            .O(N__42290),
            .I(N__42284));
    Span4Mux_h I__9828 (
            .O(N__42287),
            .I(N__42281));
    LocalMux I__9827 (
            .O(N__42284),
            .I(data_out_frame2_17_6));
    Odrv4 I__9826 (
            .O(N__42281),
            .I(data_out_frame2_17_6));
    InMux I__9825 (
            .O(N__42276),
            .I(N__42272));
    CascadeMux I__9824 (
            .O(N__42275),
            .I(N__42269));
    LocalMux I__9823 (
            .O(N__42272),
            .I(N__42266));
    InMux I__9822 (
            .O(N__42269),
            .I(N__42262));
    Span4Mux_v I__9821 (
            .O(N__42266),
            .I(N__42258));
    InMux I__9820 (
            .O(N__42265),
            .I(N__42255));
    LocalMux I__9819 (
            .O(N__42262),
            .I(N__42252));
    InMux I__9818 (
            .O(N__42261),
            .I(N__42249));
    Span4Mux_v I__9817 (
            .O(N__42258),
            .I(N__42246));
    LocalMux I__9816 (
            .O(N__42255),
            .I(N__42241));
    Span4Mux_s0_v I__9815 (
            .O(N__42252),
            .I(N__42241));
    LocalMux I__9814 (
            .O(N__42249),
            .I(data_out_frame2_16_6));
    Odrv4 I__9813 (
            .O(N__42246),
            .I(data_out_frame2_16_6));
    Odrv4 I__9812 (
            .O(N__42241),
            .I(data_out_frame2_16_6));
    CascadeMux I__9811 (
            .O(N__42234),
            .I(\c0.n18702_cascade_ ));
    InMux I__9810 (
            .O(N__42231),
            .I(N__42227));
    InMux I__9809 (
            .O(N__42230),
            .I(N__42224));
    LocalMux I__9808 (
            .O(N__42227),
            .I(N__42220));
    LocalMux I__9807 (
            .O(N__42224),
            .I(N__42217));
    InMux I__9806 (
            .O(N__42223),
            .I(N__42214));
    Span4Mux_s2_v I__9805 (
            .O(N__42220),
            .I(N__42211));
    Span4Mux_h I__9804 (
            .O(N__42217),
            .I(N__42208));
    LocalMux I__9803 (
            .O(N__42214),
            .I(data_out_frame2_13_7));
    Odrv4 I__9802 (
            .O(N__42211),
            .I(data_out_frame2_13_7));
    Odrv4 I__9801 (
            .O(N__42208),
            .I(data_out_frame2_13_7));
    InMux I__9800 (
            .O(N__42201),
            .I(N__42198));
    LocalMux I__9799 (
            .O(N__42198),
            .I(N__42195));
    Odrv12 I__9798 (
            .O(N__42195),
            .I(\c0.n10_adj_2411 ));
    InMux I__9797 (
            .O(N__42192),
            .I(N__42189));
    LocalMux I__9796 (
            .O(N__42189),
            .I(N__42186));
    Span4Mux_v I__9795 (
            .O(N__42186),
            .I(N__42183));
    Odrv4 I__9794 (
            .O(N__42183),
            .I(\c0.n18705 ));
    InMux I__9793 (
            .O(N__42180),
            .I(N__42177));
    LocalMux I__9792 (
            .O(N__42177),
            .I(N__42174));
    Span4Mux_s1_v I__9791 (
            .O(N__42174),
            .I(N__42170));
    InMux I__9790 (
            .O(N__42173),
            .I(N__42167));
    Span4Mux_v I__9789 (
            .O(N__42170),
            .I(N__42160));
    LocalMux I__9788 (
            .O(N__42167),
            .I(N__42160));
    InMux I__9787 (
            .O(N__42166),
            .I(N__42155));
    InMux I__9786 (
            .O(N__42165),
            .I(N__42155));
    Odrv4 I__9785 (
            .O(N__42160),
            .I(data_out_frame2_13_6));
    LocalMux I__9784 (
            .O(N__42155),
            .I(data_out_frame2_13_6));
    InMux I__9783 (
            .O(N__42150),
            .I(N__42145));
    InMux I__9782 (
            .O(N__42149),
            .I(N__42142));
    CascadeMux I__9781 (
            .O(N__42148),
            .I(N__42139));
    LocalMux I__9780 (
            .O(N__42145),
            .I(N__42135));
    LocalMux I__9779 (
            .O(N__42142),
            .I(N__42132));
    InMux I__9778 (
            .O(N__42139),
            .I(N__42129));
    InMux I__9777 (
            .O(N__42138),
            .I(N__42125));
    Span4Mux_h I__9776 (
            .O(N__42135),
            .I(N__42122));
    Span4Mux_v I__9775 (
            .O(N__42132),
            .I(N__42119));
    LocalMux I__9774 (
            .O(N__42129),
            .I(N__42116));
    InMux I__9773 (
            .O(N__42128),
            .I(N__42113));
    LocalMux I__9772 (
            .O(N__42125),
            .I(N__42110));
    Odrv4 I__9771 (
            .O(N__42122),
            .I(rand_data_27));
    Odrv4 I__9770 (
            .O(N__42119),
            .I(rand_data_27));
    Odrv4 I__9769 (
            .O(N__42116),
            .I(rand_data_27));
    LocalMux I__9768 (
            .O(N__42113),
            .I(rand_data_27));
    Odrv12 I__9767 (
            .O(N__42110),
            .I(rand_data_27));
    InMux I__9766 (
            .O(N__42099),
            .I(N__42092));
    InMux I__9765 (
            .O(N__42098),
            .I(N__42092));
    CascadeMux I__9764 (
            .O(N__42097),
            .I(N__42088));
    LocalMux I__9763 (
            .O(N__42092),
            .I(N__42084));
    InMux I__9762 (
            .O(N__42091),
            .I(N__42081));
    InMux I__9761 (
            .O(N__42088),
            .I(N__42077));
    InMux I__9760 (
            .O(N__42087),
            .I(N__42074));
    Span12Mux_s4_v I__9759 (
            .O(N__42084),
            .I(N__42069));
    LocalMux I__9758 (
            .O(N__42081),
            .I(N__42069));
    InMux I__9757 (
            .O(N__42080),
            .I(N__42066));
    LocalMux I__9756 (
            .O(N__42077),
            .I(N__42063));
    LocalMux I__9755 (
            .O(N__42074),
            .I(rand_data_7));
    Odrv12 I__9754 (
            .O(N__42069),
            .I(rand_data_7));
    LocalMux I__9753 (
            .O(N__42066),
            .I(rand_data_7));
    Odrv12 I__9752 (
            .O(N__42063),
            .I(rand_data_7));
    InMux I__9751 (
            .O(N__42054),
            .I(N__42049));
    InMux I__9750 (
            .O(N__42053),
            .I(N__42046));
    InMux I__9749 (
            .O(N__42052),
            .I(N__42043));
    LocalMux I__9748 (
            .O(N__42049),
            .I(N__42040));
    LocalMux I__9747 (
            .O(N__42046),
            .I(N__42036));
    LocalMux I__9746 (
            .O(N__42043),
            .I(N__42031));
    Span4Mux_h I__9745 (
            .O(N__42040),
            .I(N__42031));
    InMux I__9744 (
            .O(N__42039),
            .I(N__42028));
    Span4Mux_h I__9743 (
            .O(N__42036),
            .I(N__42025));
    Span4Mux_v I__9742 (
            .O(N__42031),
            .I(N__42022));
    LocalMux I__9741 (
            .O(N__42028),
            .I(data_out_frame2_13_3));
    Odrv4 I__9740 (
            .O(N__42025),
            .I(data_out_frame2_13_3));
    Odrv4 I__9739 (
            .O(N__42022),
            .I(data_out_frame2_13_3));
    InMux I__9738 (
            .O(N__42015),
            .I(N__42012));
    LocalMux I__9737 (
            .O(N__42012),
            .I(N__42009));
    Span4Mux_h I__9736 (
            .O(N__42009),
            .I(N__42006));
    Odrv4 I__9735 (
            .O(N__42006),
            .I(\c0.n18657 ));
    InMux I__9734 (
            .O(N__42003),
            .I(N__42000));
    LocalMux I__9733 (
            .O(N__42000),
            .I(N__41996));
    InMux I__9732 (
            .O(N__41999),
            .I(N__41993));
    Span4Mux_h I__9731 (
            .O(N__41996),
            .I(N__41990));
    LocalMux I__9730 (
            .O(N__41993),
            .I(data_out_frame2_18_3));
    Odrv4 I__9729 (
            .O(N__41990),
            .I(data_out_frame2_18_3));
    CascadeMux I__9728 (
            .O(N__41985),
            .I(N__41982));
    InMux I__9727 (
            .O(N__41982),
            .I(N__41979));
    LocalMux I__9726 (
            .O(N__41979),
            .I(N__41976));
    Odrv4 I__9725 (
            .O(N__41976),
            .I(\c0.data_out_frame2_19_3 ));
    InMux I__9724 (
            .O(N__41973),
            .I(N__41969));
    InMux I__9723 (
            .O(N__41972),
            .I(N__41966));
    LocalMux I__9722 (
            .O(N__41969),
            .I(data_out_frame2_17_3));
    LocalMux I__9721 (
            .O(N__41966),
            .I(data_out_frame2_17_3));
    CascadeMux I__9720 (
            .O(N__41961),
            .I(\c0.n18651_cascade_ ));
    InMux I__9719 (
            .O(N__41958),
            .I(N__41955));
    LocalMux I__9718 (
            .O(N__41955),
            .I(N__41951));
    InMux I__9717 (
            .O(N__41954),
            .I(N__41947));
    Span4Mux_h I__9716 (
            .O(N__41951),
            .I(N__41943));
    InMux I__9715 (
            .O(N__41950),
            .I(N__41940));
    LocalMux I__9714 (
            .O(N__41947),
            .I(N__41937));
    InMux I__9713 (
            .O(N__41946),
            .I(N__41934));
    Span4Mux_h I__9712 (
            .O(N__41943),
            .I(N__41931));
    LocalMux I__9711 (
            .O(N__41940),
            .I(N__41928));
    Span4Mux_h I__9710 (
            .O(N__41937),
            .I(N__41925));
    LocalMux I__9709 (
            .O(N__41934),
            .I(data_out_frame2_16_3));
    Odrv4 I__9708 (
            .O(N__41931),
            .I(data_out_frame2_16_3));
    Odrv4 I__9707 (
            .O(N__41928),
            .I(data_out_frame2_16_3));
    Odrv4 I__9706 (
            .O(N__41925),
            .I(data_out_frame2_16_3));
    InMux I__9705 (
            .O(N__41916),
            .I(N__41913));
    LocalMux I__9704 (
            .O(N__41913),
            .I(N__41910));
    Span4Mux_v I__9703 (
            .O(N__41910),
            .I(N__41907));
    Odrv4 I__9702 (
            .O(N__41907),
            .I(\c0.data_out_frame2_20_3 ));
    CascadeMux I__9701 (
            .O(N__41904),
            .I(\c0.n18654_cascade_ ));
    InMux I__9700 (
            .O(N__41901),
            .I(N__41898));
    LocalMux I__9699 (
            .O(N__41898),
            .I(N__41894));
    InMux I__9698 (
            .O(N__41897),
            .I(N__41891));
    Span4Mux_v I__9697 (
            .O(N__41894),
            .I(N__41888));
    LocalMux I__9696 (
            .O(N__41891),
            .I(\c0.n17880 ));
    Odrv4 I__9695 (
            .O(N__41888),
            .I(\c0.n17880 ));
    InMux I__9694 (
            .O(N__41883),
            .I(N__41879));
    InMux I__9693 (
            .O(N__41882),
            .I(N__41876));
    LocalMux I__9692 (
            .O(N__41879),
            .I(N__41873));
    LocalMux I__9691 (
            .O(N__41876),
            .I(N__41868));
    Span4Mux_s1_v I__9690 (
            .O(N__41873),
            .I(N__41868));
    Odrv4 I__9689 (
            .O(N__41868),
            .I(\c0.n17789 ));
    InMux I__9688 (
            .O(N__41865),
            .I(N__41860));
    InMux I__9687 (
            .O(N__41864),
            .I(N__41854));
    InMux I__9686 (
            .O(N__41863),
            .I(N__41854));
    LocalMux I__9685 (
            .O(N__41860),
            .I(N__41850));
    InMux I__9684 (
            .O(N__41859),
            .I(N__41847));
    LocalMux I__9683 (
            .O(N__41854),
            .I(N__41844));
    InMux I__9682 (
            .O(N__41853),
            .I(N__41841));
    Span4Mux_v I__9681 (
            .O(N__41850),
            .I(N__41836));
    LocalMux I__9680 (
            .O(N__41847),
            .I(N__41836));
    Span4Mux_h I__9679 (
            .O(N__41844),
            .I(N__41833));
    LocalMux I__9678 (
            .O(N__41841),
            .I(data_out_frame2_5_6));
    Odrv4 I__9677 (
            .O(N__41836),
            .I(data_out_frame2_5_6));
    Odrv4 I__9676 (
            .O(N__41833),
            .I(data_out_frame2_5_6));
    CascadeMux I__9675 (
            .O(N__41826),
            .I(N__41823));
    InMux I__9674 (
            .O(N__41823),
            .I(N__41820));
    LocalMux I__9673 (
            .O(N__41820),
            .I(\c0.n5_adj_2439 ));
    InMux I__9672 (
            .O(N__41817),
            .I(N__41812));
    InMux I__9671 (
            .O(N__41816),
            .I(N__41808));
    InMux I__9670 (
            .O(N__41815),
            .I(N__41805));
    LocalMux I__9669 (
            .O(N__41812),
            .I(N__41802));
    CascadeMux I__9668 (
            .O(N__41811),
            .I(N__41799));
    LocalMux I__9667 (
            .O(N__41808),
            .I(N__41796));
    LocalMux I__9666 (
            .O(N__41805),
            .I(N__41793));
    Span4Mux_h I__9665 (
            .O(N__41802),
            .I(N__41790));
    InMux I__9664 (
            .O(N__41799),
            .I(N__41787));
    Span4Mux_h I__9663 (
            .O(N__41796),
            .I(N__41782));
    Span4Mux_v I__9662 (
            .O(N__41793),
            .I(N__41782));
    Span4Mux_h I__9661 (
            .O(N__41790),
            .I(N__41779));
    LocalMux I__9660 (
            .O(N__41787),
            .I(N__41774));
    Sp12to4 I__9659 (
            .O(N__41782),
            .I(N__41774));
    Span4Mux_h I__9658 (
            .O(N__41779),
            .I(N__41771));
    Odrv12 I__9657 (
            .O(N__41774),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv4 I__9656 (
            .O(N__41771),
            .I(\c0.data_out_frame2_0_6 ));
    InMux I__9655 (
            .O(N__41766),
            .I(N__41760));
    InMux I__9654 (
            .O(N__41765),
            .I(N__41755));
    InMux I__9653 (
            .O(N__41764),
            .I(N__41755));
    InMux I__9652 (
            .O(N__41763),
            .I(N__41752));
    LocalMux I__9651 (
            .O(N__41760),
            .I(N__41748));
    LocalMux I__9650 (
            .O(N__41755),
            .I(N__41745));
    LocalMux I__9649 (
            .O(N__41752),
            .I(N__41742));
    InMux I__9648 (
            .O(N__41751),
            .I(N__41739));
    Span4Mux_h I__9647 (
            .O(N__41748),
            .I(N__41736));
    Span4Mux_h I__9646 (
            .O(N__41745),
            .I(N__41731));
    Span4Mux_h I__9645 (
            .O(N__41742),
            .I(N__41731));
    LocalMux I__9644 (
            .O(N__41739),
            .I(data_out_frame2_15_6));
    Odrv4 I__9643 (
            .O(N__41736),
            .I(data_out_frame2_15_6));
    Odrv4 I__9642 (
            .O(N__41731),
            .I(data_out_frame2_15_6));
    InMux I__9641 (
            .O(N__41724),
            .I(N__41719));
    InMux I__9640 (
            .O(N__41723),
            .I(N__41716));
    CascadeMux I__9639 (
            .O(N__41722),
            .I(N__41713));
    LocalMux I__9638 (
            .O(N__41719),
            .I(N__41710));
    LocalMux I__9637 (
            .O(N__41716),
            .I(N__41707));
    InMux I__9636 (
            .O(N__41713),
            .I(N__41704));
    Span4Mux_s2_v I__9635 (
            .O(N__41710),
            .I(N__41698));
    Span4Mux_v I__9634 (
            .O(N__41707),
            .I(N__41698));
    LocalMux I__9633 (
            .O(N__41704),
            .I(N__41695));
    InMux I__9632 (
            .O(N__41703),
            .I(N__41692));
    Span4Mux_h I__9631 (
            .O(N__41698),
            .I(N__41689));
    Span4Mux_s3_v I__9630 (
            .O(N__41695),
            .I(N__41686));
    LocalMux I__9629 (
            .O(N__41692),
            .I(data_out_frame2_13_1));
    Odrv4 I__9628 (
            .O(N__41689),
            .I(data_out_frame2_13_1));
    Odrv4 I__9627 (
            .O(N__41686),
            .I(data_out_frame2_13_1));
    InMux I__9626 (
            .O(N__41679),
            .I(N__41675));
    CascadeMux I__9625 (
            .O(N__41678),
            .I(N__41671));
    LocalMux I__9624 (
            .O(N__41675),
            .I(N__41667));
    InMux I__9623 (
            .O(N__41674),
            .I(N__41664));
    InMux I__9622 (
            .O(N__41671),
            .I(N__41661));
    InMux I__9621 (
            .O(N__41670),
            .I(N__41658));
    Span4Mux_h I__9620 (
            .O(N__41667),
            .I(N__41654));
    LocalMux I__9619 (
            .O(N__41664),
            .I(N__41651));
    LocalMux I__9618 (
            .O(N__41661),
            .I(N__41648));
    LocalMux I__9617 (
            .O(N__41658),
            .I(N__41645));
    InMux I__9616 (
            .O(N__41657),
            .I(N__41642));
    Span4Mux_s1_v I__9615 (
            .O(N__41654),
            .I(N__41639));
    Span4Mux_v I__9614 (
            .O(N__41651),
            .I(N__41632));
    Span4Mux_v I__9613 (
            .O(N__41648),
            .I(N__41632));
    Span4Mux_h I__9612 (
            .O(N__41645),
            .I(N__41632));
    LocalMux I__9611 (
            .O(N__41642),
            .I(data_out_frame2_8_7));
    Odrv4 I__9610 (
            .O(N__41639),
            .I(data_out_frame2_8_7));
    Odrv4 I__9609 (
            .O(N__41632),
            .I(data_out_frame2_8_7));
    CascadeMux I__9608 (
            .O(N__41625),
            .I(N__41621));
    InMux I__9607 (
            .O(N__41624),
            .I(N__41617));
    InMux I__9606 (
            .O(N__41621),
            .I(N__41614));
    InMux I__9605 (
            .O(N__41620),
            .I(N__41610));
    LocalMux I__9604 (
            .O(N__41617),
            .I(N__41607));
    LocalMux I__9603 (
            .O(N__41614),
            .I(N__41604));
    CascadeMux I__9602 (
            .O(N__41613),
            .I(N__41601));
    LocalMux I__9601 (
            .O(N__41610),
            .I(N__41598));
    Span4Mux_v I__9600 (
            .O(N__41607),
            .I(N__41593));
    Span4Mux_h I__9599 (
            .O(N__41604),
            .I(N__41593));
    InMux I__9598 (
            .O(N__41601),
            .I(N__41590));
    Span12Mux_h I__9597 (
            .O(N__41598),
            .I(N__41587));
    Span4Mux_h I__9596 (
            .O(N__41593),
            .I(N__41584));
    LocalMux I__9595 (
            .O(N__41590),
            .I(\c0.data_out_frame2_0_0 ));
    Odrv12 I__9594 (
            .O(N__41587),
            .I(\c0.data_out_frame2_0_0 ));
    Odrv4 I__9593 (
            .O(N__41584),
            .I(\c0.data_out_frame2_0_0 ));
    InMux I__9592 (
            .O(N__41577),
            .I(N__41574));
    LocalMux I__9591 (
            .O(N__41574),
            .I(N__41571));
    Odrv4 I__9590 (
            .O(N__41571),
            .I(\c0.n10_adj_2431 ));
    InMux I__9589 (
            .O(N__41568),
            .I(N__41561));
    InMux I__9588 (
            .O(N__41567),
            .I(N__41556));
    InMux I__9587 (
            .O(N__41566),
            .I(N__41556));
    InMux I__9586 (
            .O(N__41565),
            .I(N__41552));
    InMux I__9585 (
            .O(N__41564),
            .I(N__41549));
    LocalMux I__9584 (
            .O(N__41561),
            .I(N__41546));
    LocalMux I__9583 (
            .O(N__41556),
            .I(N__41543));
    InMux I__9582 (
            .O(N__41555),
            .I(N__41540));
    LocalMux I__9581 (
            .O(N__41552),
            .I(N__41537));
    LocalMux I__9580 (
            .O(N__41549),
            .I(N__41530));
    Span4Mux_h I__9579 (
            .O(N__41546),
            .I(N__41530));
    Span4Mux_h I__9578 (
            .O(N__41543),
            .I(N__41530));
    LocalMux I__9577 (
            .O(N__41540),
            .I(data_out_frame2_5_2));
    Odrv4 I__9576 (
            .O(N__41537),
            .I(data_out_frame2_5_2));
    Odrv4 I__9575 (
            .O(N__41530),
            .I(data_out_frame2_5_2));
    CascadeMux I__9574 (
            .O(N__41523),
            .I(N__41520));
    InMux I__9573 (
            .O(N__41520),
            .I(N__41517));
    LocalMux I__9572 (
            .O(N__41517),
            .I(N__41514));
    Sp12to4 I__9571 (
            .O(N__41514),
            .I(N__41511));
    Odrv12 I__9570 (
            .O(N__41511),
            .I(\c0.n17865 ));
    CascadeMux I__9569 (
            .O(N__41508),
            .I(N__41504));
    InMux I__9568 (
            .O(N__41507),
            .I(N__41501));
    InMux I__9567 (
            .O(N__41504),
            .I(N__41496));
    LocalMux I__9566 (
            .O(N__41501),
            .I(N__41493));
    InMux I__9565 (
            .O(N__41500),
            .I(N__41490));
    InMux I__9564 (
            .O(N__41499),
            .I(N__41487));
    LocalMux I__9563 (
            .O(N__41496),
            .I(N__41484));
    Span4Mux_v I__9562 (
            .O(N__41493),
            .I(N__41479));
    LocalMux I__9561 (
            .O(N__41490),
            .I(N__41479));
    LocalMux I__9560 (
            .O(N__41487),
            .I(N__41475));
    Span4Mux_v I__9559 (
            .O(N__41484),
            .I(N__41472));
    Span4Mux_h I__9558 (
            .O(N__41479),
            .I(N__41469));
    InMux I__9557 (
            .O(N__41478),
            .I(N__41466));
    Span4Mux_v I__9556 (
            .O(N__41475),
            .I(N__41463));
    Odrv4 I__9555 (
            .O(N__41472),
            .I(rand_data_28));
    Odrv4 I__9554 (
            .O(N__41469),
            .I(rand_data_28));
    LocalMux I__9553 (
            .O(N__41466),
            .I(rand_data_28));
    Odrv4 I__9552 (
            .O(N__41463),
            .I(rand_data_28));
    InMux I__9551 (
            .O(N__41454),
            .I(N__41448));
    InMux I__9550 (
            .O(N__41453),
            .I(N__41443));
    InMux I__9549 (
            .O(N__41452),
            .I(N__41438));
    InMux I__9548 (
            .O(N__41451),
            .I(N__41438));
    LocalMux I__9547 (
            .O(N__41448),
            .I(N__41435));
    InMux I__9546 (
            .O(N__41447),
            .I(N__41432));
    InMux I__9545 (
            .O(N__41446),
            .I(N__41429));
    LocalMux I__9544 (
            .O(N__41443),
            .I(N__41426));
    LocalMux I__9543 (
            .O(N__41438),
            .I(rand_data_11));
    Odrv4 I__9542 (
            .O(N__41435),
            .I(rand_data_11));
    LocalMux I__9541 (
            .O(N__41432),
            .I(rand_data_11));
    LocalMux I__9540 (
            .O(N__41429),
            .I(rand_data_11));
    Odrv12 I__9539 (
            .O(N__41426),
            .I(rand_data_11));
    InMux I__9538 (
            .O(N__41415),
            .I(N__41410));
    InMux I__9537 (
            .O(N__41414),
            .I(N__41407));
    InMux I__9536 (
            .O(N__41413),
            .I(N__41402));
    LocalMux I__9535 (
            .O(N__41410),
            .I(N__41399));
    LocalMux I__9534 (
            .O(N__41407),
            .I(N__41396));
    InMux I__9533 (
            .O(N__41406),
            .I(N__41393));
    InMux I__9532 (
            .O(N__41405),
            .I(N__41390));
    LocalMux I__9531 (
            .O(N__41402),
            .I(N__41383));
    Span4Mux_s3_v I__9530 (
            .O(N__41399),
            .I(N__41383));
    Span4Mux_h I__9529 (
            .O(N__41396),
            .I(N__41383));
    LocalMux I__9528 (
            .O(N__41393),
            .I(data_out_frame2_10_3));
    LocalMux I__9527 (
            .O(N__41390),
            .I(data_out_frame2_10_3));
    Odrv4 I__9526 (
            .O(N__41383),
            .I(data_out_frame2_10_3));
    InMux I__9525 (
            .O(N__41376),
            .I(N__41373));
    LocalMux I__9524 (
            .O(N__41373),
            .I(\c0.n18663 ));
    InMux I__9523 (
            .O(N__41370),
            .I(N__41367));
    LocalMux I__9522 (
            .O(N__41367),
            .I(N__41361));
    InMux I__9521 (
            .O(N__41366),
            .I(N__41358));
    InMux I__9520 (
            .O(N__41365),
            .I(N__41354));
    InMux I__9519 (
            .O(N__41364),
            .I(N__41351));
    Span12Mux_s7_v I__9518 (
            .O(N__41361),
            .I(N__41348));
    LocalMux I__9517 (
            .O(N__41358),
            .I(N__41345));
    InMux I__9516 (
            .O(N__41357),
            .I(N__41342));
    LocalMux I__9515 (
            .O(N__41354),
            .I(data_out_frame2_5_0));
    LocalMux I__9514 (
            .O(N__41351),
            .I(data_out_frame2_5_0));
    Odrv12 I__9513 (
            .O(N__41348),
            .I(data_out_frame2_5_0));
    Odrv12 I__9512 (
            .O(N__41345),
            .I(data_out_frame2_5_0));
    LocalMux I__9511 (
            .O(N__41342),
            .I(data_out_frame2_5_0));
    InMux I__9510 (
            .O(N__41331),
            .I(N__41328));
    LocalMux I__9509 (
            .O(N__41328),
            .I(\c0.n10911 ));
    InMux I__9508 (
            .O(N__41325),
            .I(N__41319));
    InMux I__9507 (
            .O(N__41324),
            .I(N__41316));
    InMux I__9506 (
            .O(N__41323),
            .I(N__41313));
    InMux I__9505 (
            .O(N__41322),
            .I(N__41309));
    LocalMux I__9504 (
            .O(N__41319),
            .I(N__41306));
    LocalMux I__9503 (
            .O(N__41316),
            .I(N__41301));
    LocalMux I__9502 (
            .O(N__41313),
            .I(N__41301));
    InMux I__9501 (
            .O(N__41312),
            .I(N__41298));
    LocalMux I__9500 (
            .O(N__41309),
            .I(data_out_frame2_11_6));
    Odrv4 I__9499 (
            .O(N__41306),
            .I(data_out_frame2_11_6));
    Odrv4 I__9498 (
            .O(N__41301),
            .I(data_out_frame2_11_6));
    LocalMux I__9497 (
            .O(N__41298),
            .I(data_out_frame2_11_6));
    InMux I__9496 (
            .O(N__41289),
            .I(N__41285));
    InMux I__9495 (
            .O(N__41288),
            .I(N__41281));
    LocalMux I__9494 (
            .O(N__41285),
            .I(N__41277));
    InMux I__9493 (
            .O(N__41284),
            .I(N__41274));
    LocalMux I__9492 (
            .O(N__41281),
            .I(N__41271));
    CascadeMux I__9491 (
            .O(N__41280),
            .I(N__41268));
    Span4Mux_h I__9490 (
            .O(N__41277),
            .I(N__41263));
    LocalMux I__9489 (
            .O(N__41274),
            .I(N__41263));
    Span4Mux_h I__9488 (
            .O(N__41271),
            .I(N__41259));
    InMux I__9487 (
            .O(N__41268),
            .I(N__41255));
    Span4Mux_v I__9486 (
            .O(N__41263),
            .I(N__41252));
    InMux I__9485 (
            .O(N__41262),
            .I(N__41249));
    Span4Mux_s2_v I__9484 (
            .O(N__41259),
            .I(N__41246));
    InMux I__9483 (
            .O(N__41258),
            .I(N__41243));
    LocalMux I__9482 (
            .O(N__41255),
            .I(N__41240));
    Odrv4 I__9481 (
            .O(N__41252),
            .I(rand_data_6));
    LocalMux I__9480 (
            .O(N__41249),
            .I(rand_data_6));
    Odrv4 I__9479 (
            .O(N__41246),
            .I(rand_data_6));
    LocalMux I__9478 (
            .O(N__41243),
            .I(rand_data_6));
    Odrv12 I__9477 (
            .O(N__41240),
            .I(rand_data_6));
    InMux I__9476 (
            .O(N__41229),
            .I(N__41224));
    InMux I__9475 (
            .O(N__41228),
            .I(N__41219));
    InMux I__9474 (
            .O(N__41227),
            .I(N__41219));
    LocalMux I__9473 (
            .O(N__41224),
            .I(N__41214));
    LocalMux I__9472 (
            .O(N__41219),
            .I(N__41211));
    InMux I__9471 (
            .O(N__41218),
            .I(N__41208));
    InMux I__9470 (
            .O(N__41217),
            .I(N__41205));
    Span4Mux_s2_v I__9469 (
            .O(N__41214),
            .I(N__41200));
    Span4Mux_h I__9468 (
            .O(N__41211),
            .I(N__41200));
    LocalMux I__9467 (
            .O(N__41208),
            .I(N__41197));
    LocalMux I__9466 (
            .O(N__41205),
            .I(data_out_frame2_9_4));
    Odrv4 I__9465 (
            .O(N__41200),
            .I(data_out_frame2_9_4));
    Odrv4 I__9464 (
            .O(N__41197),
            .I(data_out_frame2_9_4));
    InMux I__9463 (
            .O(N__41190),
            .I(N__41186));
    InMux I__9462 (
            .O(N__41189),
            .I(N__41181));
    LocalMux I__9461 (
            .O(N__41186),
            .I(N__41178));
    InMux I__9460 (
            .O(N__41185),
            .I(N__41175));
    InMux I__9459 (
            .O(N__41184),
            .I(N__41172));
    LocalMux I__9458 (
            .O(N__41181),
            .I(N__41169));
    Span4Mux_h I__9457 (
            .O(N__41178),
            .I(N__41166));
    LocalMux I__9456 (
            .O(N__41175),
            .I(N__41163));
    LocalMux I__9455 (
            .O(N__41172),
            .I(data_out_frame2_7_7));
    Odrv4 I__9454 (
            .O(N__41169),
            .I(data_out_frame2_7_7));
    Odrv4 I__9453 (
            .O(N__41166),
            .I(data_out_frame2_7_7));
    Odrv4 I__9452 (
            .O(N__41163),
            .I(data_out_frame2_7_7));
    InMux I__9451 (
            .O(N__41154),
            .I(N__41151));
    LocalMux I__9450 (
            .O(N__41151),
            .I(N__41146));
    CascadeMux I__9449 (
            .O(N__41150),
            .I(N__41142));
    InMux I__9448 (
            .O(N__41149),
            .I(N__41139));
    Span12Mux_h I__9447 (
            .O(N__41146),
            .I(N__41136));
    InMux I__9446 (
            .O(N__41145),
            .I(N__41133));
    InMux I__9445 (
            .O(N__41142),
            .I(N__41130));
    LocalMux I__9444 (
            .O(N__41139),
            .I(data_out_frame2_9_7));
    Odrv12 I__9443 (
            .O(N__41136),
            .I(data_out_frame2_9_7));
    LocalMux I__9442 (
            .O(N__41133),
            .I(data_out_frame2_9_7));
    LocalMux I__9441 (
            .O(N__41130),
            .I(data_out_frame2_9_7));
    CascadeMux I__9440 (
            .O(N__41121),
            .I(N__41118));
    InMux I__9439 (
            .O(N__41118),
            .I(N__41115));
    LocalMux I__9438 (
            .O(N__41115),
            .I(N__41112));
    Odrv4 I__9437 (
            .O(N__41112),
            .I(\c0.n10617 ));
    InMux I__9436 (
            .O(N__41109),
            .I(N__41106));
    LocalMux I__9435 (
            .O(N__41106),
            .I(N__41103));
    Span4Mux_s2_v I__9434 (
            .O(N__41103),
            .I(N__41100));
    Span4Mux_h I__9433 (
            .O(N__41100),
            .I(N__41097));
    Odrv4 I__9432 (
            .O(N__41097),
            .I(\c0.n14_adj_2362 ));
    CascadeMux I__9431 (
            .O(N__41094),
            .I(N__41091));
    InMux I__9430 (
            .O(N__41091),
            .I(N__41086));
    InMux I__9429 (
            .O(N__41090),
            .I(N__41083));
    InMux I__9428 (
            .O(N__41089),
            .I(N__41079));
    LocalMux I__9427 (
            .O(N__41086),
            .I(N__41073));
    LocalMux I__9426 (
            .O(N__41083),
            .I(N__41070));
    InMux I__9425 (
            .O(N__41082),
            .I(N__41067));
    LocalMux I__9424 (
            .O(N__41079),
            .I(N__41064));
    InMux I__9423 (
            .O(N__41078),
            .I(N__41059));
    InMux I__9422 (
            .O(N__41077),
            .I(N__41059));
    InMux I__9421 (
            .O(N__41076),
            .I(N__41056));
    Span4Mux_h I__9420 (
            .O(N__41073),
            .I(N__41051));
    Span4Mux_v I__9419 (
            .O(N__41070),
            .I(N__41051));
    LocalMux I__9418 (
            .O(N__41067),
            .I(N__41044));
    Span4Mux_h I__9417 (
            .O(N__41064),
            .I(N__41044));
    LocalMux I__9416 (
            .O(N__41059),
            .I(N__41044));
    LocalMux I__9415 (
            .O(N__41056),
            .I(data_out_frame2_12_2));
    Odrv4 I__9414 (
            .O(N__41051),
            .I(data_out_frame2_12_2));
    Odrv4 I__9413 (
            .O(N__41044),
            .I(data_out_frame2_12_2));
    InMux I__9412 (
            .O(N__41037),
            .I(N__41032));
    InMux I__9411 (
            .O(N__41036),
            .I(N__41029));
    InMux I__9410 (
            .O(N__41035),
            .I(N__41026));
    LocalMux I__9409 (
            .O(N__41032),
            .I(N__41022));
    LocalMux I__9408 (
            .O(N__41029),
            .I(N__41019));
    LocalMux I__9407 (
            .O(N__41026),
            .I(N__41016));
    InMux I__9406 (
            .O(N__41025),
            .I(N__41012));
    Span4Mux_v I__9405 (
            .O(N__41022),
            .I(N__41009));
    Span4Mux_h I__9404 (
            .O(N__41019),
            .I(N__41004));
    Span4Mux_s1_v I__9403 (
            .O(N__41016),
            .I(N__41004));
    InMux I__9402 (
            .O(N__41015),
            .I(N__41001));
    LocalMux I__9401 (
            .O(N__41012),
            .I(data_out_frame2_10_4));
    Odrv4 I__9400 (
            .O(N__41009),
            .I(data_out_frame2_10_4));
    Odrv4 I__9399 (
            .O(N__41004),
            .I(data_out_frame2_10_4));
    LocalMux I__9398 (
            .O(N__41001),
            .I(data_out_frame2_10_4));
    InMux I__9397 (
            .O(N__40992),
            .I(N__40988));
    InMux I__9396 (
            .O(N__40991),
            .I(N__40985));
    LocalMux I__9395 (
            .O(N__40988),
            .I(N__40980));
    LocalMux I__9394 (
            .O(N__40985),
            .I(N__40977));
    InMux I__9393 (
            .O(N__40984),
            .I(N__40973));
    InMux I__9392 (
            .O(N__40983),
            .I(N__40970));
    Span4Mux_s2_v I__9391 (
            .O(N__40980),
            .I(N__40967));
    Span4Mux_s2_v I__9390 (
            .O(N__40977),
            .I(N__40964));
    InMux I__9389 (
            .O(N__40976),
            .I(N__40961));
    LocalMux I__9388 (
            .O(N__40973),
            .I(data_out_frame2_16_7));
    LocalMux I__9387 (
            .O(N__40970),
            .I(data_out_frame2_16_7));
    Odrv4 I__9386 (
            .O(N__40967),
            .I(data_out_frame2_16_7));
    Odrv4 I__9385 (
            .O(N__40964),
            .I(data_out_frame2_16_7));
    LocalMux I__9384 (
            .O(N__40961),
            .I(data_out_frame2_16_7));
    InMux I__9383 (
            .O(N__40950),
            .I(N__40946));
    InMux I__9382 (
            .O(N__40949),
            .I(N__40943));
    LocalMux I__9381 (
            .O(N__40946),
            .I(N__40937));
    LocalMux I__9380 (
            .O(N__40943),
            .I(N__40934));
    InMux I__9379 (
            .O(N__40942),
            .I(N__40929));
    InMux I__9378 (
            .O(N__40941),
            .I(N__40929));
    InMux I__9377 (
            .O(N__40940),
            .I(N__40925));
    Span4Mux_v I__9376 (
            .O(N__40937),
            .I(N__40918));
    Span4Mux_s0_v I__9375 (
            .O(N__40934),
            .I(N__40918));
    LocalMux I__9374 (
            .O(N__40929),
            .I(N__40918));
    InMux I__9373 (
            .O(N__40928),
            .I(N__40915));
    LocalMux I__9372 (
            .O(N__40925),
            .I(N__40910));
    Span4Mux_h I__9371 (
            .O(N__40918),
            .I(N__40910));
    LocalMux I__9370 (
            .O(N__40915),
            .I(data_out_frame2_15_7));
    Odrv4 I__9369 (
            .O(N__40910),
            .I(data_out_frame2_15_7));
    InMux I__9368 (
            .O(N__40905),
            .I(N__40902));
    LocalMux I__9367 (
            .O(N__40902),
            .I(\c0.n17889 ));
    InMux I__9366 (
            .O(N__40899),
            .I(N__40896));
    LocalMux I__9365 (
            .O(N__40896),
            .I(N__40893));
    Span4Mux_h I__9364 (
            .O(N__40893),
            .I(N__40888));
    InMux I__9363 (
            .O(N__40892),
            .I(N__40885));
    InMux I__9362 (
            .O(N__40891),
            .I(N__40882));
    Span4Mux_s2_v I__9361 (
            .O(N__40888),
            .I(N__40877));
    LocalMux I__9360 (
            .O(N__40885),
            .I(N__40877));
    LocalMux I__9359 (
            .O(N__40882),
            .I(N__40873));
    Span4Mux_h I__9358 (
            .O(N__40877),
            .I(N__40870));
    InMux I__9357 (
            .O(N__40876),
            .I(N__40866));
    Span4Mux_h I__9356 (
            .O(N__40873),
            .I(N__40863));
    Span4Mux_v I__9355 (
            .O(N__40870),
            .I(N__40860));
    InMux I__9354 (
            .O(N__40869),
            .I(N__40857));
    LocalMux I__9353 (
            .O(N__40866),
            .I(N__40854));
    Odrv4 I__9352 (
            .O(N__40863),
            .I(rand_data_18));
    Odrv4 I__9351 (
            .O(N__40860),
            .I(rand_data_18));
    LocalMux I__9350 (
            .O(N__40857),
            .I(rand_data_18));
    Odrv12 I__9349 (
            .O(N__40854),
            .I(rand_data_18));
    CascadeMux I__9348 (
            .O(N__40845),
            .I(N__40841));
    InMux I__9347 (
            .O(N__40844),
            .I(N__40836));
    InMux I__9346 (
            .O(N__40841),
            .I(N__40831));
    InMux I__9345 (
            .O(N__40840),
            .I(N__40831));
    InMux I__9344 (
            .O(N__40839),
            .I(N__40828));
    LocalMux I__9343 (
            .O(N__40836),
            .I(N__40825));
    LocalMux I__9342 (
            .O(N__40831),
            .I(N__40822));
    LocalMux I__9341 (
            .O(N__40828),
            .I(data_out_frame2_6_2));
    Odrv12 I__9340 (
            .O(N__40825),
            .I(data_out_frame2_6_2));
    Odrv4 I__9339 (
            .O(N__40822),
            .I(data_out_frame2_6_2));
    InMux I__9338 (
            .O(N__40815),
            .I(N__40812));
    LocalMux I__9337 (
            .O(N__40812),
            .I(N__40809));
    Span4Mux_h I__9336 (
            .O(N__40809),
            .I(N__40806));
    Odrv4 I__9335 (
            .O(N__40806),
            .I(\c0.n18645 ));
    InMux I__9334 (
            .O(N__40803),
            .I(N__40800));
    LocalMux I__9333 (
            .O(N__40800),
            .I(N__40797));
    Span12Mux_h I__9332 (
            .O(N__40797),
            .I(N__40794));
    Odrv12 I__9331 (
            .O(N__40794),
            .I(\c0.n18_adj_2441 ));
    InMux I__9330 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__9329 (
            .O(N__40788),
            .I(N__40783));
    InMux I__9328 (
            .O(N__40787),
            .I(N__40778));
    InMux I__9327 (
            .O(N__40786),
            .I(N__40778));
    Span4Mux_s2_v I__9326 (
            .O(N__40783),
            .I(N__40772));
    LocalMux I__9325 (
            .O(N__40778),
            .I(N__40769));
    InMux I__9324 (
            .O(N__40777),
            .I(N__40766));
    InMux I__9323 (
            .O(N__40776),
            .I(N__40761));
    InMux I__9322 (
            .O(N__40775),
            .I(N__40761));
    Odrv4 I__9321 (
            .O(N__40772),
            .I(data_out_frame2_8_3));
    Odrv12 I__9320 (
            .O(N__40769),
            .I(data_out_frame2_8_3));
    LocalMux I__9319 (
            .O(N__40766),
            .I(data_out_frame2_8_3));
    LocalMux I__9318 (
            .O(N__40761),
            .I(data_out_frame2_8_3));
    InMux I__9317 (
            .O(N__40752),
            .I(N__40747));
    InMux I__9316 (
            .O(N__40751),
            .I(N__40743));
    CascadeMux I__9315 (
            .O(N__40750),
            .I(N__40740));
    LocalMux I__9314 (
            .O(N__40747),
            .I(N__40736));
    InMux I__9313 (
            .O(N__40746),
            .I(N__40733));
    LocalMux I__9312 (
            .O(N__40743),
            .I(N__40730));
    InMux I__9311 (
            .O(N__40740),
            .I(N__40725));
    InMux I__9310 (
            .O(N__40739),
            .I(N__40725));
    Span4Mux_h I__9309 (
            .O(N__40736),
            .I(N__40722));
    LocalMux I__9308 (
            .O(N__40733),
            .I(N__40719));
    Span4Mux_s2_v I__9307 (
            .O(N__40730),
            .I(N__40716));
    LocalMux I__9306 (
            .O(N__40725),
            .I(data_out_frame2_10_1));
    Odrv4 I__9305 (
            .O(N__40722),
            .I(data_out_frame2_10_1));
    Odrv4 I__9304 (
            .O(N__40719),
            .I(data_out_frame2_10_1));
    Odrv4 I__9303 (
            .O(N__40716),
            .I(data_out_frame2_10_1));
    InMux I__9302 (
            .O(N__40707),
            .I(N__40704));
    LocalMux I__9301 (
            .O(N__40704),
            .I(N__40700));
    InMux I__9300 (
            .O(N__40703),
            .I(N__40697));
    Span4Mux_h I__9299 (
            .O(N__40700),
            .I(N__40694));
    LocalMux I__9298 (
            .O(N__40697),
            .I(\c0.n17838 ));
    Odrv4 I__9297 (
            .O(N__40694),
            .I(\c0.n17838 ));
    InMux I__9296 (
            .O(N__40689),
            .I(N__40685));
    InMux I__9295 (
            .O(N__40688),
            .I(N__40682));
    LocalMux I__9294 (
            .O(N__40685),
            .I(N__40679));
    LocalMux I__9293 (
            .O(N__40682),
            .I(N__40676));
    Odrv12 I__9292 (
            .O(N__40679),
            .I(\c0.n17792 ));
    Odrv4 I__9291 (
            .O(N__40676),
            .I(\c0.n17792 ));
    InMux I__9290 (
            .O(N__40671),
            .I(N__40668));
    LocalMux I__9289 (
            .O(N__40668),
            .I(\c0.n33 ));
    InMux I__9288 (
            .O(N__40665),
            .I(N__40661));
    InMux I__9287 (
            .O(N__40664),
            .I(N__40658));
    LocalMux I__9286 (
            .O(N__40661),
            .I(N__40653));
    LocalMux I__9285 (
            .O(N__40658),
            .I(N__40650));
    InMux I__9284 (
            .O(N__40657),
            .I(N__40647));
    InMux I__9283 (
            .O(N__40656),
            .I(N__40644));
    Span12Mux_s9_v I__9282 (
            .O(N__40653),
            .I(N__40641));
    Span12Mux_s2_v I__9281 (
            .O(N__40650),
            .I(N__40638));
    LocalMux I__9280 (
            .O(N__40647),
            .I(data_out_frame2_6_6));
    LocalMux I__9279 (
            .O(N__40644),
            .I(data_out_frame2_6_6));
    Odrv12 I__9278 (
            .O(N__40641),
            .I(data_out_frame2_6_6));
    Odrv12 I__9277 (
            .O(N__40638),
            .I(data_out_frame2_6_6));
    CascadeMux I__9276 (
            .O(N__40629),
            .I(N__40626));
    InMux I__9275 (
            .O(N__40626),
            .I(N__40623));
    LocalMux I__9274 (
            .O(N__40623),
            .I(N__40620));
    Span4Mux_h I__9273 (
            .O(N__40620),
            .I(N__40617));
    Sp12to4 I__9272 (
            .O(N__40617),
            .I(N__40614));
    Odrv12 I__9271 (
            .O(N__40614),
            .I(\c0.n17736 ));
    CascadeMux I__9270 (
            .O(N__40611),
            .I(\c0.n17736_cascade_ ));
    InMux I__9269 (
            .O(N__40608),
            .I(N__40605));
    LocalMux I__9268 (
            .O(N__40605),
            .I(\c0.n18813 ));
    CascadeMux I__9267 (
            .O(N__40602),
            .I(N__40599));
    InMux I__9266 (
            .O(N__40599),
            .I(N__40596));
    LocalMux I__9265 (
            .O(N__40596),
            .I(N__40593));
    Odrv12 I__9264 (
            .O(N__40593),
            .I(\c0.n18816 ));
    InMux I__9263 (
            .O(N__40590),
            .I(N__40582));
    InMux I__9262 (
            .O(N__40589),
            .I(N__40582));
    InMux I__9261 (
            .O(N__40588),
            .I(N__40577));
    InMux I__9260 (
            .O(N__40587),
            .I(N__40577));
    LocalMux I__9259 (
            .O(N__40582),
            .I(N__40571));
    LocalMux I__9258 (
            .O(N__40577),
            .I(N__40571));
    InMux I__9257 (
            .O(N__40576),
            .I(N__40568));
    Span4Mux_s1_v I__9256 (
            .O(N__40571),
            .I(N__40565));
    LocalMux I__9255 (
            .O(N__40568),
            .I(data_out_frame2_9_6));
    Odrv4 I__9254 (
            .O(N__40565),
            .I(data_out_frame2_9_6));
    InMux I__9253 (
            .O(N__40560),
            .I(N__40557));
    LocalMux I__9252 (
            .O(N__40557),
            .I(N__40554));
    Odrv12 I__9251 (
            .O(N__40554),
            .I(\c0.n10725 ));
    InMux I__9250 (
            .O(N__40551),
            .I(N__40546));
    InMux I__9249 (
            .O(N__40550),
            .I(N__40543));
    InMux I__9248 (
            .O(N__40549),
            .I(N__40540));
    LocalMux I__9247 (
            .O(N__40546),
            .I(N__40537));
    LocalMux I__9246 (
            .O(N__40543),
            .I(N__40530));
    LocalMux I__9245 (
            .O(N__40540),
            .I(N__40530));
    Span4Mux_v I__9244 (
            .O(N__40537),
            .I(N__40527));
    InMux I__9243 (
            .O(N__40536),
            .I(N__40524));
    InMux I__9242 (
            .O(N__40535),
            .I(N__40521));
    Span4Mux_h I__9241 (
            .O(N__40530),
            .I(N__40516));
    Span4Mux_v I__9240 (
            .O(N__40527),
            .I(N__40516));
    LocalMux I__9239 (
            .O(N__40524),
            .I(data_out_frame2_7_0));
    LocalMux I__9238 (
            .O(N__40521),
            .I(data_out_frame2_7_0));
    Odrv4 I__9237 (
            .O(N__40516),
            .I(data_out_frame2_7_0));
    CascadeMux I__9236 (
            .O(N__40509),
            .I(N__40506));
    InMux I__9235 (
            .O(N__40506),
            .I(N__40503));
    LocalMux I__9234 (
            .O(N__40503),
            .I(N__40500));
    Span4Mux_h I__9233 (
            .O(N__40500),
            .I(N__40497));
    IoSpan4Mux I__9232 (
            .O(N__40497),
            .I(N__40494));
    Odrv4 I__9231 (
            .O(N__40494),
            .I(\c0.n10700 ));
    InMux I__9230 (
            .O(N__40491),
            .I(N__40488));
    LocalMux I__9229 (
            .O(N__40488),
            .I(N__40485));
    Span12Mux_h I__9228 (
            .O(N__40485),
            .I(N__40482));
    Odrv12 I__9227 (
            .O(N__40482),
            .I(\c0.n16_adj_2412 ));
    CascadeMux I__9226 (
            .O(N__40479),
            .I(\c0.n17_adj_2413_cascade_ ));
    InMux I__9225 (
            .O(N__40476),
            .I(N__40472));
    InMux I__9224 (
            .O(N__40475),
            .I(N__40469));
    LocalMux I__9223 (
            .O(N__40472),
            .I(N__40463));
    LocalMux I__9222 (
            .O(N__40469),
            .I(N__40463));
    InMux I__9221 (
            .O(N__40468),
            .I(N__40459));
    Span4Mux_v I__9220 (
            .O(N__40463),
            .I(N__40456));
    CascadeMux I__9219 (
            .O(N__40462),
            .I(N__40453));
    LocalMux I__9218 (
            .O(N__40459),
            .I(N__40448));
    Sp12to4 I__9217 (
            .O(N__40456),
            .I(N__40448));
    InMux I__9216 (
            .O(N__40453),
            .I(N__40445));
    Span12Mux_h I__9215 (
            .O(N__40448),
            .I(N__40442));
    LocalMux I__9214 (
            .O(N__40445),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv12 I__9213 (
            .O(N__40442),
            .I(\c0.data_out_frame2_0_1 ));
    InMux I__9212 (
            .O(N__40437),
            .I(N__40433));
    CascadeMux I__9211 (
            .O(N__40436),
            .I(N__40430));
    LocalMux I__9210 (
            .O(N__40433),
            .I(N__40427));
    InMux I__9209 (
            .O(N__40430),
            .I(N__40424));
    Span4Mux_h I__9208 (
            .O(N__40427),
            .I(N__40421));
    LocalMux I__9207 (
            .O(N__40424),
            .I(N__40418));
    Span4Mux_v I__9206 (
            .O(N__40421),
            .I(N__40415));
    Span12Mux_s8_v I__9205 (
            .O(N__40418),
            .I(N__40412));
    Odrv4 I__9204 (
            .O(N__40415),
            .I(\c0.n10782 ));
    Odrv12 I__9203 (
            .O(N__40412),
            .I(\c0.n10782 ));
    InMux I__9202 (
            .O(N__40407),
            .I(N__40403));
    CascadeMux I__9201 (
            .O(N__40406),
            .I(N__40400));
    LocalMux I__9200 (
            .O(N__40403),
            .I(N__40397));
    InMux I__9199 (
            .O(N__40400),
            .I(N__40393));
    IoSpan4Mux I__9198 (
            .O(N__40397),
            .I(N__40390));
    InMux I__9197 (
            .O(N__40396),
            .I(N__40386));
    LocalMux I__9196 (
            .O(N__40393),
            .I(N__40381));
    IoSpan4Mux I__9195 (
            .O(N__40390),
            .I(N__40381));
    InMux I__9194 (
            .O(N__40389),
            .I(N__40378));
    LocalMux I__9193 (
            .O(N__40386),
            .I(data_out_frame2_14_1));
    Odrv4 I__9192 (
            .O(N__40381),
            .I(data_out_frame2_14_1));
    LocalMux I__9191 (
            .O(N__40378),
            .I(data_out_frame2_14_1));
    InMux I__9190 (
            .O(N__40371),
            .I(N__40368));
    LocalMux I__9189 (
            .O(N__40368),
            .I(\c0.n17862 ));
    CascadeMux I__9188 (
            .O(N__40365),
            .I(\c0.n17862_cascade_ ));
    InMux I__9187 (
            .O(N__40362),
            .I(N__40359));
    LocalMux I__9186 (
            .O(N__40359),
            .I(N__40356));
    Span4Mux_h I__9185 (
            .O(N__40356),
            .I(N__40352));
    InMux I__9184 (
            .O(N__40355),
            .I(N__40349));
    Odrv4 I__9183 (
            .O(N__40352),
            .I(\c0.n17841 ));
    LocalMux I__9182 (
            .O(N__40349),
            .I(\c0.n17841 ));
    CascadeMux I__9181 (
            .O(N__40344),
            .I(\c0.n12_adj_2410_cascade_ ));
    InMux I__9180 (
            .O(N__40341),
            .I(N__40338));
    LocalMux I__9179 (
            .O(N__40338),
            .I(N__40335));
    Span4Mux_h I__9178 (
            .O(N__40335),
            .I(N__40331));
    InMux I__9177 (
            .O(N__40334),
            .I(N__40328));
    Odrv4 I__9176 (
            .O(N__40331),
            .I(\c0.n17718 ));
    LocalMux I__9175 (
            .O(N__40328),
            .I(\c0.n17718 ));
    InMux I__9174 (
            .O(N__40323),
            .I(N__40319));
    InMux I__9173 (
            .O(N__40322),
            .I(N__40316));
    LocalMux I__9172 (
            .O(N__40319),
            .I(\c0.n17829 ));
    LocalMux I__9171 (
            .O(N__40316),
            .I(\c0.n17829 ));
    InMux I__9170 (
            .O(N__40311),
            .I(N__40306));
    InMux I__9169 (
            .O(N__40310),
            .I(N__40303));
    InMux I__9168 (
            .O(N__40309),
            .I(N__40300));
    LocalMux I__9167 (
            .O(N__40306),
            .I(N__40297));
    LocalMux I__9166 (
            .O(N__40303),
            .I(N__40294));
    LocalMux I__9165 (
            .O(N__40300),
            .I(N__40291));
    Span4Mux_v I__9164 (
            .O(N__40297),
            .I(N__40286));
    Span4Mux_h I__9163 (
            .O(N__40294),
            .I(N__40286));
    Odrv4 I__9162 (
            .O(N__40291),
            .I(\c0.data_out_10_4 ));
    Odrv4 I__9161 (
            .O(N__40286),
            .I(\c0.data_out_10_4 ));
    InMux I__9160 (
            .O(N__40281),
            .I(N__40278));
    LocalMux I__9159 (
            .O(N__40278),
            .I(N__40274));
    InMux I__9158 (
            .O(N__40277),
            .I(N__40271));
    Span4Mux_v I__9157 (
            .O(N__40274),
            .I(N__40267));
    LocalMux I__9156 (
            .O(N__40271),
            .I(N__40264));
    InMux I__9155 (
            .O(N__40270),
            .I(N__40261));
    Span4Mux_h I__9154 (
            .O(N__40267),
            .I(N__40258));
    Span4Mux_h I__9153 (
            .O(N__40264),
            .I(N__40255));
    LocalMux I__9152 (
            .O(N__40261),
            .I(N__40252));
    Odrv4 I__9151 (
            .O(N__40258),
            .I(n2837));
    Odrv4 I__9150 (
            .O(N__40255),
            .I(n2837));
    Odrv4 I__9149 (
            .O(N__40252),
            .I(n2837));
    InMux I__9148 (
            .O(N__40245),
            .I(N__40239));
    InMux I__9147 (
            .O(N__40244),
            .I(N__40239));
    LocalMux I__9146 (
            .O(N__40239),
            .I(data_out_3_0));
    InMux I__9145 (
            .O(N__40236),
            .I(N__40233));
    LocalMux I__9144 (
            .O(N__40233),
            .I(N__40230));
    Odrv4 I__9143 (
            .O(N__40230),
            .I(\c0.n2_adj_2221 ));
    InMux I__9142 (
            .O(N__40227),
            .I(N__40221));
    InMux I__9141 (
            .O(N__40226),
            .I(N__40221));
    LocalMux I__9140 (
            .O(N__40221),
            .I(data_out_2_0));
    InMux I__9139 (
            .O(N__40218),
            .I(N__40215));
    LocalMux I__9138 (
            .O(N__40215),
            .I(N__40212));
    Span4Mux_s0_v I__9137 (
            .O(N__40212),
            .I(N__40209));
    Span4Mux_h I__9136 (
            .O(N__40209),
            .I(N__40206));
    Odrv4 I__9135 (
            .O(N__40206),
            .I(\c0.n5_adj_2433 ));
    InMux I__9134 (
            .O(N__40203),
            .I(N__40200));
    LocalMux I__9133 (
            .O(N__40200),
            .I(N__40194));
    InMux I__9132 (
            .O(N__40199),
            .I(N__40189));
    InMux I__9131 (
            .O(N__40198),
            .I(N__40189));
    InMux I__9130 (
            .O(N__40197),
            .I(N__40186));
    Span4Mux_s2_v I__9129 (
            .O(N__40194),
            .I(N__40183));
    LocalMux I__9128 (
            .O(N__40189),
            .I(N__40180));
    LocalMux I__9127 (
            .O(N__40186),
            .I(data_out_frame2_14_7));
    Odrv4 I__9126 (
            .O(N__40183),
            .I(data_out_frame2_14_7));
    Odrv4 I__9125 (
            .O(N__40180),
            .I(data_out_frame2_14_7));
    InMux I__9124 (
            .O(N__40173),
            .I(N__40170));
    LocalMux I__9123 (
            .O(N__40170),
            .I(\c0.n17899 ));
    CascadeMux I__9122 (
            .O(N__40167),
            .I(\c0.n17899_cascade_ ));
    InMux I__9121 (
            .O(N__40164),
            .I(N__40161));
    LocalMux I__9120 (
            .O(N__40161),
            .I(N__40158));
    Span4Mux_v I__9119 (
            .O(N__40158),
            .I(N__40155));
    Span4Mux_s0_v I__9118 (
            .O(N__40155),
            .I(N__40152));
    Odrv4 I__9117 (
            .O(N__40152),
            .I(\c0.n34 ));
    InMux I__9116 (
            .O(N__40149),
            .I(N__40143));
    InMux I__9115 (
            .O(N__40148),
            .I(N__40140));
    InMux I__9114 (
            .O(N__40147),
            .I(N__40137));
    InMux I__9113 (
            .O(N__40146),
            .I(N__40134));
    LocalMux I__9112 (
            .O(N__40143),
            .I(N__40131));
    LocalMux I__9111 (
            .O(N__40140),
            .I(N__40126));
    LocalMux I__9110 (
            .O(N__40137),
            .I(N__40126));
    LocalMux I__9109 (
            .O(N__40134),
            .I(N__40122));
    Span4Mux_h I__9108 (
            .O(N__40131),
            .I(N__40119));
    Span4Mux_v I__9107 (
            .O(N__40126),
            .I(N__40116));
    InMux I__9106 (
            .O(N__40125),
            .I(N__40113));
    Span4Mux_v I__9105 (
            .O(N__40122),
            .I(N__40110));
    Odrv4 I__9104 (
            .O(N__40119),
            .I(rand_data_30));
    Odrv4 I__9103 (
            .O(N__40116),
            .I(rand_data_30));
    LocalMux I__9102 (
            .O(N__40113),
            .I(rand_data_30));
    Odrv4 I__9101 (
            .O(N__40110),
            .I(rand_data_30));
    InMux I__9100 (
            .O(N__40101),
            .I(n16607));
    InMux I__9099 (
            .O(N__40098),
            .I(N__40093));
    InMux I__9098 (
            .O(N__40097),
            .I(N__40089));
    InMux I__9097 (
            .O(N__40096),
            .I(N__40086));
    LocalMux I__9096 (
            .O(N__40093),
            .I(N__40083));
    InMux I__9095 (
            .O(N__40092),
            .I(N__40080));
    LocalMux I__9094 (
            .O(N__40089),
            .I(N__40077));
    LocalMux I__9093 (
            .O(N__40086),
            .I(N__40073));
    Span4Mux_h I__9092 (
            .O(N__40083),
            .I(N__40070));
    LocalMux I__9091 (
            .O(N__40080),
            .I(N__40067));
    Span4Mux_s3_v I__9090 (
            .O(N__40077),
            .I(N__40064));
    InMux I__9089 (
            .O(N__40076),
            .I(N__40061));
    Span4Mux_v I__9088 (
            .O(N__40073),
            .I(N__40058));
    Span4Mux_v I__9087 (
            .O(N__40070),
            .I(N__40051));
    Span4Mux_v I__9086 (
            .O(N__40067),
            .I(N__40051));
    Span4Mux_v I__9085 (
            .O(N__40064),
            .I(N__40051));
    LocalMux I__9084 (
            .O(N__40061),
            .I(rand_data_31));
    Odrv4 I__9083 (
            .O(N__40058),
            .I(rand_data_31));
    Odrv4 I__9082 (
            .O(N__40051),
            .I(rand_data_31));
    InMux I__9081 (
            .O(N__40044),
            .I(n16608));
    InMux I__9080 (
            .O(N__40041),
            .I(N__40037));
    CascadeMux I__9079 (
            .O(N__40040),
            .I(N__40034));
    LocalMux I__9078 (
            .O(N__40037),
            .I(N__40031));
    InMux I__9077 (
            .O(N__40034),
            .I(N__40028));
    Odrv4 I__9076 (
            .O(N__40031),
            .I(rand_setpoint_13));
    LocalMux I__9075 (
            .O(N__40028),
            .I(rand_setpoint_13));
    CascadeMux I__9074 (
            .O(N__40023),
            .I(N__40020));
    InMux I__9073 (
            .O(N__40020),
            .I(N__40017));
    LocalMux I__9072 (
            .O(N__40017),
            .I(N__40014));
    Odrv4 I__9071 (
            .O(N__40014),
            .I(\c0.n18234 ));
    InMux I__9070 (
            .O(N__40011),
            .I(N__40007));
    CascadeMux I__9069 (
            .O(N__40010),
            .I(N__40004));
    LocalMux I__9068 (
            .O(N__40007),
            .I(N__40001));
    InMux I__9067 (
            .O(N__40004),
            .I(N__39998));
    Odrv12 I__9066 (
            .O(N__40001),
            .I(rand_setpoint_1));
    LocalMux I__9065 (
            .O(N__39998),
            .I(rand_setpoint_1));
    CascadeMux I__9064 (
            .O(N__39993),
            .I(N__39990));
    InMux I__9063 (
            .O(N__39990),
            .I(N__39987));
    LocalMux I__9062 (
            .O(N__39987),
            .I(N__39981));
    InMux I__9061 (
            .O(N__39986),
            .I(N__39978));
    InMux I__9060 (
            .O(N__39985),
            .I(N__39973));
    InMux I__9059 (
            .O(N__39984),
            .I(N__39973));
    Span4Mux_v I__9058 (
            .O(N__39981),
            .I(N__39969));
    LocalMux I__9057 (
            .O(N__39978),
            .I(N__39966));
    LocalMux I__9056 (
            .O(N__39973),
            .I(N__39963));
    InMux I__9055 (
            .O(N__39972),
            .I(N__39960));
    Span4Mux_v I__9054 (
            .O(N__39969),
            .I(N__39957));
    Span4Mux_h I__9053 (
            .O(N__39966),
            .I(N__39954));
    Span4Mux_h I__9052 (
            .O(N__39963),
            .I(N__39951));
    LocalMux I__9051 (
            .O(N__39960),
            .I(\c0.data_out_8_1 ));
    Odrv4 I__9050 (
            .O(N__39957),
            .I(\c0.data_out_8_1 ));
    Odrv4 I__9049 (
            .O(N__39954),
            .I(\c0.data_out_8_1 ));
    Odrv4 I__9048 (
            .O(N__39951),
            .I(\c0.data_out_8_1 ));
    InMux I__9047 (
            .O(N__39942),
            .I(N__39938));
    InMux I__9046 (
            .O(N__39941),
            .I(N__39935));
    LocalMux I__9045 (
            .O(N__39938),
            .I(N__39932));
    LocalMux I__9044 (
            .O(N__39935),
            .I(N__39927));
    Span4Mux_h I__9043 (
            .O(N__39932),
            .I(N__39924));
    InMux I__9042 (
            .O(N__39931),
            .I(N__39919));
    InMux I__9041 (
            .O(N__39930),
            .I(N__39919));
    Span4Mux_h I__9040 (
            .O(N__39927),
            .I(N__39916));
    Odrv4 I__9039 (
            .O(N__39924),
            .I(\c0.data_out_7_5 ));
    LocalMux I__9038 (
            .O(N__39919),
            .I(\c0.data_out_7_5 ));
    Odrv4 I__9037 (
            .O(N__39916),
            .I(\c0.data_out_7_5 ));
    InMux I__9036 (
            .O(N__39909),
            .I(N__39904));
    InMux I__9035 (
            .O(N__39908),
            .I(N__39901));
    InMux I__9034 (
            .O(N__39907),
            .I(N__39897));
    LocalMux I__9033 (
            .O(N__39904),
            .I(N__39894));
    LocalMux I__9032 (
            .O(N__39901),
            .I(N__39890));
    InMux I__9031 (
            .O(N__39900),
            .I(N__39887));
    LocalMux I__9030 (
            .O(N__39897),
            .I(N__39884));
    Span4Mux_h I__9029 (
            .O(N__39894),
            .I(N__39881));
    InMux I__9028 (
            .O(N__39893),
            .I(N__39878));
    Span4Mux_h I__9027 (
            .O(N__39890),
            .I(N__39875));
    LocalMux I__9026 (
            .O(N__39887),
            .I(\c0.data_out_7_7 ));
    Odrv12 I__9025 (
            .O(N__39884),
            .I(\c0.data_out_7_7 ));
    Odrv4 I__9024 (
            .O(N__39881),
            .I(\c0.data_out_7_7 ));
    LocalMux I__9023 (
            .O(N__39878),
            .I(\c0.data_out_7_7 ));
    Odrv4 I__9022 (
            .O(N__39875),
            .I(\c0.data_out_7_7 ));
    InMux I__9021 (
            .O(N__39864),
            .I(N__39861));
    LocalMux I__9020 (
            .O(N__39861),
            .I(N__39858));
    Odrv4 I__9019 (
            .O(N__39858),
            .I(\c0.n10533 ));
    InMux I__9018 (
            .O(N__39855),
            .I(N__39851));
    CascadeMux I__9017 (
            .O(N__39854),
            .I(N__39848));
    LocalMux I__9016 (
            .O(N__39851),
            .I(N__39845));
    InMux I__9015 (
            .O(N__39848),
            .I(N__39842));
    Odrv4 I__9014 (
            .O(N__39845),
            .I(rand_setpoint_26));
    LocalMux I__9013 (
            .O(N__39842),
            .I(rand_setpoint_26));
    InMux I__9012 (
            .O(N__39837),
            .I(N__39831));
    InMux I__9011 (
            .O(N__39836),
            .I(N__39826));
    InMux I__9010 (
            .O(N__39835),
            .I(N__39826));
    InMux I__9009 (
            .O(N__39834),
            .I(N__39823));
    LocalMux I__9008 (
            .O(N__39831),
            .I(N__39816));
    LocalMux I__9007 (
            .O(N__39826),
            .I(N__39816));
    LocalMux I__9006 (
            .O(N__39823),
            .I(N__39813));
    InMux I__9005 (
            .O(N__39822),
            .I(N__39810));
    InMux I__9004 (
            .O(N__39821),
            .I(N__39807));
    Span4Mux_h I__9003 (
            .O(N__39816),
            .I(N__39804));
    Span4Mux_h I__9002 (
            .O(N__39813),
            .I(N__39801));
    LocalMux I__9001 (
            .O(N__39810),
            .I(\c0.data_out_5_2 ));
    LocalMux I__9000 (
            .O(N__39807),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__8999 (
            .O(N__39804),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__8998 (
            .O(N__39801),
            .I(\c0.data_out_5_2 ));
    InMux I__8997 (
            .O(N__39792),
            .I(N__39788));
    CascadeMux I__8996 (
            .O(N__39791),
            .I(N__39785));
    LocalMux I__8995 (
            .O(N__39788),
            .I(N__39782));
    InMux I__8994 (
            .O(N__39785),
            .I(N__39779));
    Odrv4 I__8993 (
            .O(N__39782),
            .I(rand_setpoint_30));
    LocalMux I__8992 (
            .O(N__39779),
            .I(rand_setpoint_30));
    InMux I__8991 (
            .O(N__39774),
            .I(N__39770));
    CascadeMux I__8990 (
            .O(N__39773),
            .I(N__39767));
    LocalMux I__8989 (
            .O(N__39770),
            .I(N__39764));
    InMux I__8988 (
            .O(N__39767),
            .I(N__39761));
    Odrv4 I__8987 (
            .O(N__39764),
            .I(rand_setpoint_27));
    LocalMux I__8986 (
            .O(N__39761),
            .I(rand_setpoint_27));
    InMux I__8985 (
            .O(N__39756),
            .I(N__39752));
    InMux I__8984 (
            .O(N__39755),
            .I(N__39747));
    LocalMux I__8983 (
            .O(N__39752),
            .I(N__39744));
    InMux I__8982 (
            .O(N__39751),
            .I(N__39736));
    InMux I__8981 (
            .O(N__39750),
            .I(N__39736));
    LocalMux I__8980 (
            .O(N__39747),
            .I(N__39733));
    Span4Mux_v I__8979 (
            .O(N__39744),
            .I(N__39730));
    InMux I__8978 (
            .O(N__39743),
            .I(N__39727));
    InMux I__8977 (
            .O(N__39742),
            .I(N__39722));
    InMux I__8976 (
            .O(N__39741),
            .I(N__39722));
    LocalMux I__8975 (
            .O(N__39736),
            .I(N__39719));
    Span4Mux_h I__8974 (
            .O(N__39733),
            .I(N__39716));
    Odrv4 I__8973 (
            .O(N__39730),
            .I(\c0.data_out_5_3 ));
    LocalMux I__8972 (
            .O(N__39727),
            .I(\c0.data_out_5_3 ));
    LocalMux I__8971 (
            .O(N__39722),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__8970 (
            .O(N__39719),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__8969 (
            .O(N__39716),
            .I(\c0.data_out_5_3 ));
    InMux I__8968 (
            .O(N__39705),
            .I(N__39701));
    InMux I__8967 (
            .O(N__39704),
            .I(N__39696));
    LocalMux I__8966 (
            .O(N__39701),
            .I(N__39693));
    InMux I__8965 (
            .O(N__39700),
            .I(N__39690));
    InMux I__8964 (
            .O(N__39699),
            .I(N__39687));
    LocalMux I__8963 (
            .O(N__39696),
            .I(N__39684));
    Span4Mux_v I__8962 (
            .O(N__39693),
            .I(N__39681));
    LocalMux I__8961 (
            .O(N__39690),
            .I(N__39677));
    LocalMux I__8960 (
            .O(N__39687),
            .I(N__39674));
    Span4Mux_h I__8959 (
            .O(N__39684),
            .I(N__39669));
    Span4Mux_h I__8958 (
            .O(N__39681),
            .I(N__39669));
    InMux I__8957 (
            .O(N__39680),
            .I(N__39666));
    Span4Mux_h I__8956 (
            .O(N__39677),
            .I(N__39661));
    Span4Mux_v I__8955 (
            .O(N__39674),
            .I(N__39661));
    Odrv4 I__8954 (
            .O(N__39669),
            .I(rand_data_22));
    LocalMux I__8953 (
            .O(N__39666),
            .I(rand_data_22));
    Odrv4 I__8952 (
            .O(N__39661),
            .I(rand_data_22));
    InMux I__8951 (
            .O(N__39654),
            .I(N__39650));
    CascadeMux I__8950 (
            .O(N__39653),
            .I(N__39647));
    LocalMux I__8949 (
            .O(N__39650),
            .I(N__39644));
    InMux I__8948 (
            .O(N__39647),
            .I(N__39641));
    Odrv4 I__8947 (
            .O(N__39644),
            .I(rand_setpoint_22));
    LocalMux I__8946 (
            .O(N__39641),
            .I(rand_setpoint_22));
    InMux I__8945 (
            .O(N__39636),
            .I(n16599));
    CascadeMux I__8944 (
            .O(N__39633),
            .I(N__39629));
    InMux I__8943 (
            .O(N__39632),
            .I(N__39626));
    InMux I__8942 (
            .O(N__39629),
            .I(N__39621));
    LocalMux I__8941 (
            .O(N__39626),
            .I(N__39618));
    InMux I__8940 (
            .O(N__39625),
            .I(N__39615));
    InMux I__8939 (
            .O(N__39624),
            .I(N__39612));
    LocalMux I__8938 (
            .O(N__39621),
            .I(N__39609));
    Span4Mux_h I__8937 (
            .O(N__39618),
            .I(N__39606));
    LocalMux I__8936 (
            .O(N__39615),
            .I(N__39603));
    LocalMux I__8935 (
            .O(N__39612),
            .I(N__39599));
    Span4Mux_v I__8934 (
            .O(N__39609),
            .I(N__39596));
    Span4Mux_v I__8933 (
            .O(N__39606),
            .I(N__39591));
    Span4Mux_v I__8932 (
            .O(N__39603),
            .I(N__39591));
    InMux I__8931 (
            .O(N__39602),
            .I(N__39588));
    Span4Mux_v I__8930 (
            .O(N__39599),
            .I(N__39585));
    Odrv4 I__8929 (
            .O(N__39596),
            .I(rand_data_23));
    Odrv4 I__8928 (
            .O(N__39591),
            .I(rand_data_23));
    LocalMux I__8927 (
            .O(N__39588),
            .I(rand_data_23));
    Odrv4 I__8926 (
            .O(N__39585),
            .I(rand_data_23));
    CascadeMux I__8925 (
            .O(N__39576),
            .I(N__39572));
    CascadeMux I__8924 (
            .O(N__39575),
            .I(N__39569));
    InMux I__8923 (
            .O(N__39572),
            .I(N__39566));
    InMux I__8922 (
            .O(N__39569),
            .I(N__39563));
    LocalMux I__8921 (
            .O(N__39566),
            .I(rand_setpoint_23));
    LocalMux I__8920 (
            .O(N__39563),
            .I(rand_setpoint_23));
    InMux I__8919 (
            .O(N__39558),
            .I(n16600));
    InMux I__8918 (
            .O(N__39555),
            .I(N__39549));
    InMux I__8917 (
            .O(N__39554),
            .I(N__39546));
    InMux I__8916 (
            .O(N__39553),
            .I(N__39543));
    CascadeMux I__8915 (
            .O(N__39552),
            .I(N__39540));
    LocalMux I__8914 (
            .O(N__39549),
            .I(N__39534));
    LocalMux I__8913 (
            .O(N__39546),
            .I(N__39534));
    LocalMux I__8912 (
            .O(N__39543),
            .I(N__39531));
    InMux I__8911 (
            .O(N__39540),
            .I(N__39528));
    InMux I__8910 (
            .O(N__39539),
            .I(N__39525));
    Span4Mux_h I__8909 (
            .O(N__39534),
            .I(N__39520));
    Span4Mux_v I__8908 (
            .O(N__39531),
            .I(N__39520));
    LocalMux I__8907 (
            .O(N__39528),
            .I(rand_data_24));
    LocalMux I__8906 (
            .O(N__39525),
            .I(rand_data_24));
    Odrv4 I__8905 (
            .O(N__39520),
            .I(rand_data_24));
    InMux I__8904 (
            .O(N__39513),
            .I(bfn_14_12_0_));
    InMux I__8903 (
            .O(N__39510),
            .I(N__39507));
    LocalMux I__8902 (
            .O(N__39507),
            .I(N__39504));
    Span4Mux_h I__8901 (
            .O(N__39504),
            .I(N__39499));
    InMux I__8900 (
            .O(N__39503),
            .I(N__39496));
    InMux I__8899 (
            .O(N__39502),
            .I(N__39493));
    Span4Mux_v I__8898 (
            .O(N__39499),
            .I(N__39489));
    LocalMux I__8897 (
            .O(N__39496),
            .I(N__39484));
    LocalMux I__8896 (
            .O(N__39493),
            .I(N__39484));
    InMux I__8895 (
            .O(N__39492),
            .I(N__39481));
    Sp12to4 I__8894 (
            .O(N__39489),
            .I(N__39478));
    Span4Mux_h I__8893 (
            .O(N__39484),
            .I(N__39474));
    LocalMux I__8892 (
            .O(N__39481),
            .I(N__39471));
    Span12Mux_v I__8891 (
            .O(N__39478),
            .I(N__39468));
    InMux I__8890 (
            .O(N__39477),
            .I(N__39465));
    Span4Mux_v I__8889 (
            .O(N__39474),
            .I(N__39460));
    Span4Mux_v I__8888 (
            .O(N__39471),
            .I(N__39460));
    Odrv12 I__8887 (
            .O(N__39468),
            .I(rand_data_25));
    LocalMux I__8886 (
            .O(N__39465),
            .I(rand_data_25));
    Odrv4 I__8885 (
            .O(N__39460),
            .I(rand_data_25));
    CascadeMux I__8884 (
            .O(N__39453),
            .I(N__39450));
    InMux I__8883 (
            .O(N__39450),
            .I(N__39447));
    LocalMux I__8882 (
            .O(N__39447),
            .I(N__39443));
    CascadeMux I__8881 (
            .O(N__39446),
            .I(N__39440));
    Span4Mux_v I__8880 (
            .O(N__39443),
            .I(N__39437));
    InMux I__8879 (
            .O(N__39440),
            .I(N__39434));
    Odrv4 I__8878 (
            .O(N__39437),
            .I(rand_setpoint_25));
    LocalMux I__8877 (
            .O(N__39434),
            .I(rand_setpoint_25));
    InMux I__8876 (
            .O(N__39429),
            .I(n16602));
    InMux I__8875 (
            .O(N__39426),
            .I(N__39419));
    InMux I__8874 (
            .O(N__39425),
            .I(N__39419));
    InMux I__8873 (
            .O(N__39424),
            .I(N__39416));
    LocalMux I__8872 (
            .O(N__39419),
            .I(N__39412));
    LocalMux I__8871 (
            .O(N__39416),
            .I(N__39408));
    InMux I__8870 (
            .O(N__39415),
            .I(N__39405));
    Span4Mux_h I__8869 (
            .O(N__39412),
            .I(N__39402));
    InMux I__8868 (
            .O(N__39411),
            .I(N__39399));
    Span12Mux_s5_v I__8867 (
            .O(N__39408),
            .I(N__39394));
    LocalMux I__8866 (
            .O(N__39405),
            .I(N__39394));
    Odrv4 I__8865 (
            .O(N__39402),
            .I(rand_data_26));
    LocalMux I__8864 (
            .O(N__39399),
            .I(rand_data_26));
    Odrv12 I__8863 (
            .O(N__39394),
            .I(rand_data_26));
    InMux I__8862 (
            .O(N__39387),
            .I(n16603));
    InMux I__8861 (
            .O(N__39384),
            .I(n16604));
    InMux I__8860 (
            .O(N__39381),
            .I(N__39378));
    LocalMux I__8859 (
            .O(N__39378),
            .I(N__39375));
    Span4Mux_v I__8858 (
            .O(N__39375),
            .I(N__39371));
    CascadeMux I__8857 (
            .O(N__39374),
            .I(N__39368));
    Span4Mux_v I__8856 (
            .O(N__39371),
            .I(N__39365));
    InMux I__8855 (
            .O(N__39368),
            .I(N__39362));
    Odrv4 I__8854 (
            .O(N__39365),
            .I(rand_setpoint_28));
    LocalMux I__8853 (
            .O(N__39362),
            .I(rand_setpoint_28));
    InMux I__8852 (
            .O(N__39357),
            .I(n16605));
    InMux I__8851 (
            .O(N__39354),
            .I(N__39351));
    LocalMux I__8850 (
            .O(N__39351),
            .I(N__39347));
    InMux I__8849 (
            .O(N__39350),
            .I(N__39344));
    Span4Mux_h I__8848 (
            .O(N__39347),
            .I(N__39337));
    LocalMux I__8847 (
            .O(N__39344),
            .I(N__39337));
    InMux I__8846 (
            .O(N__39343),
            .I(N__39334));
    InMux I__8845 (
            .O(N__39342),
            .I(N__39331));
    Span4Mux_h I__8844 (
            .O(N__39337),
            .I(N__39326));
    LocalMux I__8843 (
            .O(N__39334),
            .I(N__39326));
    LocalMux I__8842 (
            .O(N__39331),
            .I(N__39322));
    Span4Mux_v I__8841 (
            .O(N__39326),
            .I(N__39319));
    InMux I__8840 (
            .O(N__39325),
            .I(N__39316));
    Span4Mux_v I__8839 (
            .O(N__39322),
            .I(N__39313));
    Odrv4 I__8838 (
            .O(N__39319),
            .I(rand_data_29));
    LocalMux I__8837 (
            .O(N__39316),
            .I(rand_data_29));
    Odrv4 I__8836 (
            .O(N__39313),
            .I(rand_data_29));
    CascadeMux I__8835 (
            .O(N__39306),
            .I(N__39302));
    InMux I__8834 (
            .O(N__39305),
            .I(N__39299));
    InMux I__8833 (
            .O(N__39302),
            .I(N__39296));
    LocalMux I__8832 (
            .O(N__39299),
            .I(rand_setpoint_29));
    LocalMux I__8831 (
            .O(N__39296),
            .I(rand_setpoint_29));
    InMux I__8830 (
            .O(N__39291),
            .I(n16606));
    CascadeMux I__8829 (
            .O(N__39288),
            .I(N__39284));
    InMux I__8828 (
            .O(N__39287),
            .I(N__39279));
    InMux I__8827 (
            .O(N__39284),
            .I(N__39275));
    InMux I__8826 (
            .O(N__39283),
            .I(N__39272));
    InMux I__8825 (
            .O(N__39282),
            .I(N__39269));
    LocalMux I__8824 (
            .O(N__39279),
            .I(N__39266));
    InMux I__8823 (
            .O(N__39278),
            .I(N__39262));
    LocalMux I__8822 (
            .O(N__39275),
            .I(N__39257));
    LocalMux I__8821 (
            .O(N__39272),
            .I(N__39257));
    LocalMux I__8820 (
            .O(N__39269),
            .I(N__39252));
    Span4Mux_v I__8819 (
            .O(N__39266),
            .I(N__39252));
    InMux I__8818 (
            .O(N__39265),
            .I(N__39249));
    LocalMux I__8817 (
            .O(N__39262),
            .I(N__39244));
    Sp12to4 I__8816 (
            .O(N__39257),
            .I(N__39244));
    Odrv4 I__8815 (
            .O(N__39252),
            .I(rand_data_14));
    LocalMux I__8814 (
            .O(N__39249),
            .I(rand_data_14));
    Odrv12 I__8813 (
            .O(N__39244),
            .I(rand_data_14));
    InMux I__8812 (
            .O(N__39237),
            .I(n16591));
    InMux I__8811 (
            .O(N__39234),
            .I(N__39225));
    InMux I__8810 (
            .O(N__39233),
            .I(N__39225));
    InMux I__8809 (
            .O(N__39232),
            .I(N__39222));
    InMux I__8808 (
            .O(N__39231),
            .I(N__39219));
    CascadeMux I__8807 (
            .O(N__39230),
            .I(N__39216));
    LocalMux I__8806 (
            .O(N__39225),
            .I(N__39213));
    LocalMux I__8805 (
            .O(N__39222),
            .I(N__39208));
    LocalMux I__8804 (
            .O(N__39219),
            .I(N__39208));
    InMux I__8803 (
            .O(N__39216),
            .I(N__39204));
    Span4Mux_h I__8802 (
            .O(N__39213),
            .I(N__39201));
    Span4Mux_h I__8801 (
            .O(N__39208),
            .I(N__39198));
    InMux I__8800 (
            .O(N__39207),
            .I(N__39195));
    LocalMux I__8799 (
            .O(N__39204),
            .I(N__39192));
    Odrv4 I__8798 (
            .O(N__39201),
            .I(rand_data_15));
    Odrv4 I__8797 (
            .O(N__39198),
            .I(rand_data_15));
    LocalMux I__8796 (
            .O(N__39195),
            .I(rand_data_15));
    Odrv12 I__8795 (
            .O(N__39192),
            .I(rand_data_15));
    InMux I__8794 (
            .O(N__39183),
            .I(N__39180));
    LocalMux I__8793 (
            .O(N__39180),
            .I(N__39177));
    Span4Mux_h I__8792 (
            .O(N__39177),
            .I(N__39174));
    Span4Mux_v I__8791 (
            .O(N__39174),
            .I(N__39170));
    InMux I__8790 (
            .O(N__39173),
            .I(N__39167));
    Odrv4 I__8789 (
            .O(N__39170),
            .I(rand_setpoint_15));
    LocalMux I__8788 (
            .O(N__39167),
            .I(rand_setpoint_15));
    InMux I__8787 (
            .O(N__39162),
            .I(n16592));
    CascadeMux I__8786 (
            .O(N__39159),
            .I(N__39156));
    InMux I__8785 (
            .O(N__39156),
            .I(N__39152));
    InMux I__8784 (
            .O(N__39155),
            .I(N__39149));
    LocalMux I__8783 (
            .O(N__39152),
            .I(N__39143));
    LocalMux I__8782 (
            .O(N__39149),
            .I(N__39143));
    InMux I__8781 (
            .O(N__39148),
            .I(N__39140));
    Span4Mux_v I__8780 (
            .O(N__39143),
            .I(N__39137));
    LocalMux I__8779 (
            .O(N__39140),
            .I(N__39132));
    Span4Mux_h I__8778 (
            .O(N__39137),
            .I(N__39129));
    InMux I__8777 (
            .O(N__39136),
            .I(N__39126));
    InMux I__8776 (
            .O(N__39135),
            .I(N__39123));
    Span4Mux_v I__8775 (
            .O(N__39132),
            .I(N__39120));
    Odrv4 I__8774 (
            .O(N__39129),
            .I(rand_data_16));
    LocalMux I__8773 (
            .O(N__39126),
            .I(rand_data_16));
    LocalMux I__8772 (
            .O(N__39123),
            .I(rand_data_16));
    Odrv4 I__8771 (
            .O(N__39120),
            .I(rand_data_16));
    InMux I__8770 (
            .O(N__39111),
            .I(N__39108));
    LocalMux I__8769 (
            .O(N__39108),
            .I(N__39104));
    CascadeMux I__8768 (
            .O(N__39107),
            .I(N__39101));
    Span4Mux_v I__8767 (
            .O(N__39104),
            .I(N__39098));
    InMux I__8766 (
            .O(N__39101),
            .I(N__39095));
    Odrv4 I__8765 (
            .O(N__39098),
            .I(rand_setpoint_16));
    LocalMux I__8764 (
            .O(N__39095),
            .I(rand_setpoint_16));
    InMux I__8763 (
            .O(N__39090),
            .I(bfn_14_11_0_));
    InMux I__8762 (
            .O(N__39087),
            .I(N__39082));
    InMux I__8761 (
            .O(N__39086),
            .I(N__39079));
    InMux I__8760 (
            .O(N__39085),
            .I(N__39076));
    LocalMux I__8759 (
            .O(N__39082),
            .I(N__39071));
    LocalMux I__8758 (
            .O(N__39079),
            .I(N__39071));
    LocalMux I__8757 (
            .O(N__39076),
            .I(N__39067));
    Span4Mux_v I__8756 (
            .O(N__39071),
            .I(N__39064));
    InMux I__8755 (
            .O(N__39070),
            .I(N__39061));
    Span4Mux_v I__8754 (
            .O(N__39067),
            .I(N__39056));
    Span4Mux_s2_v I__8753 (
            .O(N__39064),
            .I(N__39056));
    LocalMux I__8752 (
            .O(N__39061),
            .I(N__39052));
    Span4Mux_h I__8751 (
            .O(N__39056),
            .I(N__39049));
    InMux I__8750 (
            .O(N__39055),
            .I(N__39046));
    Span4Mux_v I__8749 (
            .O(N__39052),
            .I(N__39043));
    Odrv4 I__8748 (
            .O(N__39049),
            .I(rand_data_17));
    LocalMux I__8747 (
            .O(N__39046),
            .I(rand_data_17));
    Odrv4 I__8746 (
            .O(N__39043),
            .I(rand_data_17));
    InMux I__8745 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__8744 (
            .O(N__39033),
            .I(N__39030));
    Span4Mux_v I__8743 (
            .O(N__39030),
            .I(N__39027));
    Span4Mux_h I__8742 (
            .O(N__39027),
            .I(N__39023));
    CascadeMux I__8741 (
            .O(N__39026),
            .I(N__39020));
    Span4Mux_h I__8740 (
            .O(N__39023),
            .I(N__39017));
    InMux I__8739 (
            .O(N__39020),
            .I(N__39014));
    Odrv4 I__8738 (
            .O(N__39017),
            .I(rand_setpoint_17));
    LocalMux I__8737 (
            .O(N__39014),
            .I(rand_setpoint_17));
    InMux I__8736 (
            .O(N__39009),
            .I(n16594));
    InMux I__8735 (
            .O(N__39006),
            .I(N__39003));
    LocalMux I__8734 (
            .O(N__39003),
            .I(N__38999));
    CascadeMux I__8733 (
            .O(N__39002),
            .I(N__38996));
    Span4Mux_h I__8732 (
            .O(N__38999),
            .I(N__38993));
    InMux I__8731 (
            .O(N__38996),
            .I(N__38990));
    Odrv4 I__8730 (
            .O(N__38993),
            .I(rand_setpoint_18));
    LocalMux I__8729 (
            .O(N__38990),
            .I(rand_setpoint_18));
    InMux I__8728 (
            .O(N__38985),
            .I(n16595));
    InMux I__8727 (
            .O(N__38982),
            .I(N__38976));
    InMux I__8726 (
            .O(N__38981),
            .I(N__38973));
    InMux I__8725 (
            .O(N__38980),
            .I(N__38970));
    InMux I__8724 (
            .O(N__38979),
            .I(N__38967));
    LocalMux I__8723 (
            .O(N__38976),
            .I(N__38964));
    LocalMux I__8722 (
            .O(N__38973),
            .I(N__38961));
    LocalMux I__8721 (
            .O(N__38970),
            .I(N__38957));
    LocalMux I__8720 (
            .O(N__38967),
            .I(N__38954));
    Span4Mux_v I__8719 (
            .O(N__38964),
            .I(N__38951));
    Span4Mux_v I__8718 (
            .O(N__38961),
            .I(N__38948));
    InMux I__8717 (
            .O(N__38960),
            .I(N__38945));
    Span4Mux_v I__8716 (
            .O(N__38957),
            .I(N__38940));
    Span4Mux_v I__8715 (
            .O(N__38954),
            .I(N__38940));
    Odrv4 I__8714 (
            .O(N__38951),
            .I(rand_data_19));
    Odrv4 I__8713 (
            .O(N__38948),
            .I(rand_data_19));
    LocalMux I__8712 (
            .O(N__38945),
            .I(rand_data_19));
    Odrv4 I__8711 (
            .O(N__38940),
            .I(rand_data_19));
    InMux I__8710 (
            .O(N__38931),
            .I(N__38928));
    LocalMux I__8709 (
            .O(N__38928),
            .I(N__38924));
    CascadeMux I__8708 (
            .O(N__38927),
            .I(N__38921));
    Span4Mux_h I__8707 (
            .O(N__38924),
            .I(N__38918));
    InMux I__8706 (
            .O(N__38921),
            .I(N__38915));
    Odrv4 I__8705 (
            .O(N__38918),
            .I(rand_setpoint_19));
    LocalMux I__8704 (
            .O(N__38915),
            .I(rand_setpoint_19));
    InMux I__8703 (
            .O(N__38910),
            .I(n16596));
    InMux I__8702 (
            .O(N__38907),
            .I(N__38901));
    InMux I__8701 (
            .O(N__38906),
            .I(N__38898));
    CascadeMux I__8700 (
            .O(N__38905),
            .I(N__38895));
    CascadeMux I__8699 (
            .O(N__38904),
            .I(N__38892));
    LocalMux I__8698 (
            .O(N__38901),
            .I(N__38888));
    LocalMux I__8697 (
            .O(N__38898),
            .I(N__38885));
    InMux I__8696 (
            .O(N__38895),
            .I(N__38880));
    InMux I__8695 (
            .O(N__38892),
            .I(N__38880));
    InMux I__8694 (
            .O(N__38891),
            .I(N__38877));
    Span4Mux_h I__8693 (
            .O(N__38888),
            .I(N__38872));
    Span4Mux_v I__8692 (
            .O(N__38885),
            .I(N__38872));
    LocalMux I__8691 (
            .O(N__38880),
            .I(rand_data_20));
    LocalMux I__8690 (
            .O(N__38877),
            .I(rand_data_20));
    Odrv4 I__8689 (
            .O(N__38872),
            .I(rand_data_20));
    CascadeMux I__8688 (
            .O(N__38865),
            .I(N__38861));
    InMux I__8687 (
            .O(N__38864),
            .I(N__38858));
    InMux I__8686 (
            .O(N__38861),
            .I(N__38855));
    LocalMux I__8685 (
            .O(N__38858),
            .I(rand_setpoint_20));
    LocalMux I__8684 (
            .O(N__38855),
            .I(rand_setpoint_20));
    InMux I__8683 (
            .O(N__38850),
            .I(n16597));
    InMux I__8682 (
            .O(N__38847),
            .I(N__38843));
    InMux I__8681 (
            .O(N__38846),
            .I(N__38840));
    LocalMux I__8680 (
            .O(N__38843),
            .I(N__38835));
    LocalMux I__8679 (
            .O(N__38840),
            .I(N__38832));
    InMux I__8678 (
            .O(N__38839),
            .I(N__38829));
    InMux I__8677 (
            .O(N__38838),
            .I(N__38826));
    Span4Mux_h I__8676 (
            .O(N__38835),
            .I(N__38823));
    Span4Mux_v I__8675 (
            .O(N__38832),
            .I(N__38820));
    LocalMux I__8674 (
            .O(N__38829),
            .I(N__38817));
    LocalMux I__8673 (
            .O(N__38826),
            .I(N__38813));
    Span4Mux_h I__8672 (
            .O(N__38823),
            .I(N__38810));
    Span4Mux_h I__8671 (
            .O(N__38820),
            .I(N__38805));
    Span4Mux_v I__8670 (
            .O(N__38817),
            .I(N__38805));
    InMux I__8669 (
            .O(N__38816),
            .I(N__38802));
    Span4Mux_v I__8668 (
            .O(N__38813),
            .I(N__38799));
    Odrv4 I__8667 (
            .O(N__38810),
            .I(rand_data_21));
    Odrv4 I__8666 (
            .O(N__38805),
            .I(rand_data_21));
    LocalMux I__8665 (
            .O(N__38802),
            .I(rand_data_21));
    Odrv4 I__8664 (
            .O(N__38799),
            .I(rand_data_21));
    CascadeMux I__8663 (
            .O(N__38790),
            .I(N__38786));
    InMux I__8662 (
            .O(N__38789),
            .I(N__38783));
    InMux I__8661 (
            .O(N__38786),
            .I(N__38780));
    LocalMux I__8660 (
            .O(N__38783),
            .I(rand_setpoint_21));
    LocalMux I__8659 (
            .O(N__38780),
            .I(rand_setpoint_21));
    InMux I__8658 (
            .O(N__38775),
            .I(n16598));
    InMux I__8657 (
            .O(N__38772),
            .I(N__38769));
    LocalMux I__8656 (
            .O(N__38769),
            .I(N__38766));
    Span4Mux_v I__8655 (
            .O(N__38766),
            .I(N__38763));
    Span4Mux_v I__8654 (
            .O(N__38763),
            .I(N__38759));
    InMux I__8653 (
            .O(N__38762),
            .I(N__38756));
    Odrv4 I__8652 (
            .O(N__38759),
            .I(rand_setpoint_6));
    LocalMux I__8651 (
            .O(N__38756),
            .I(rand_setpoint_6));
    InMux I__8650 (
            .O(N__38751),
            .I(n16583));
    InMux I__8649 (
            .O(N__38748),
            .I(N__38745));
    LocalMux I__8648 (
            .O(N__38745),
            .I(N__38742));
    Span4Mux_v I__8647 (
            .O(N__38742),
            .I(N__38739));
    Span4Mux_h I__8646 (
            .O(N__38739),
            .I(N__38735));
    InMux I__8645 (
            .O(N__38738),
            .I(N__38732));
    Odrv4 I__8644 (
            .O(N__38735),
            .I(rand_setpoint_7));
    LocalMux I__8643 (
            .O(N__38732),
            .I(rand_setpoint_7));
    InMux I__8642 (
            .O(N__38727),
            .I(n16584));
    CascadeMux I__8641 (
            .O(N__38724),
            .I(N__38721));
    InMux I__8640 (
            .O(N__38721),
            .I(N__38716));
    InMux I__8639 (
            .O(N__38720),
            .I(N__38712));
    InMux I__8638 (
            .O(N__38719),
            .I(N__38709));
    LocalMux I__8637 (
            .O(N__38716),
            .I(N__38706));
    InMux I__8636 (
            .O(N__38715),
            .I(N__38703));
    LocalMux I__8635 (
            .O(N__38712),
            .I(N__38699));
    LocalMux I__8634 (
            .O(N__38709),
            .I(N__38694));
    Span4Mux_s1_v I__8633 (
            .O(N__38706),
            .I(N__38694));
    LocalMux I__8632 (
            .O(N__38703),
            .I(N__38690));
    InMux I__8631 (
            .O(N__38702),
            .I(N__38687));
    Span4Mux_h I__8630 (
            .O(N__38699),
            .I(N__38684));
    Span4Mux_v I__8629 (
            .O(N__38694),
            .I(N__38681));
    InMux I__8628 (
            .O(N__38693),
            .I(N__38678));
    Sp12to4 I__8627 (
            .O(N__38690),
            .I(N__38673));
    LocalMux I__8626 (
            .O(N__38687),
            .I(N__38673));
    Odrv4 I__8625 (
            .O(N__38684),
            .I(rand_data_8));
    Odrv4 I__8624 (
            .O(N__38681),
            .I(rand_data_8));
    LocalMux I__8623 (
            .O(N__38678),
            .I(rand_data_8));
    Odrv12 I__8622 (
            .O(N__38673),
            .I(rand_data_8));
    InMux I__8621 (
            .O(N__38664),
            .I(bfn_14_10_0_));
    InMux I__8620 (
            .O(N__38661),
            .I(N__38657));
    InMux I__8619 (
            .O(N__38660),
            .I(N__38654));
    LocalMux I__8618 (
            .O(N__38657),
            .I(N__38651));
    LocalMux I__8617 (
            .O(N__38654),
            .I(N__38646));
    Span4Mux_s1_v I__8616 (
            .O(N__38651),
            .I(N__38643));
    InMux I__8615 (
            .O(N__38650),
            .I(N__38640));
    InMux I__8614 (
            .O(N__38649),
            .I(N__38636));
    Span4Mux_s2_v I__8613 (
            .O(N__38646),
            .I(N__38633));
    Span4Mux_h I__8612 (
            .O(N__38643),
            .I(N__38630));
    LocalMux I__8611 (
            .O(N__38640),
            .I(N__38627));
    InMux I__8610 (
            .O(N__38639),
            .I(N__38623));
    LocalMux I__8609 (
            .O(N__38636),
            .I(N__38620));
    Span4Mux_h I__8608 (
            .O(N__38633),
            .I(N__38617));
    Span4Mux_v I__8607 (
            .O(N__38630),
            .I(N__38612));
    Span4Mux_h I__8606 (
            .O(N__38627),
            .I(N__38612));
    InMux I__8605 (
            .O(N__38626),
            .I(N__38609));
    LocalMux I__8604 (
            .O(N__38623),
            .I(N__38604));
    Span4Mux_v I__8603 (
            .O(N__38620),
            .I(N__38604));
    Odrv4 I__8602 (
            .O(N__38617),
            .I(rand_data_9));
    Odrv4 I__8601 (
            .O(N__38612),
            .I(rand_data_9));
    LocalMux I__8600 (
            .O(N__38609),
            .I(rand_data_9));
    Odrv4 I__8599 (
            .O(N__38604),
            .I(rand_data_9));
    CascadeMux I__8598 (
            .O(N__38595),
            .I(N__38592));
    InMux I__8597 (
            .O(N__38592),
            .I(N__38589));
    LocalMux I__8596 (
            .O(N__38589),
            .I(N__38585));
    CascadeMux I__8595 (
            .O(N__38588),
            .I(N__38582));
    Span4Mux_v I__8594 (
            .O(N__38585),
            .I(N__38579));
    InMux I__8593 (
            .O(N__38582),
            .I(N__38576));
    Odrv4 I__8592 (
            .O(N__38579),
            .I(rand_setpoint_9));
    LocalMux I__8591 (
            .O(N__38576),
            .I(rand_setpoint_9));
    InMux I__8590 (
            .O(N__38571),
            .I(n16586));
    InMux I__8589 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__8588 (
            .O(N__38565),
            .I(N__38560));
    InMux I__8587 (
            .O(N__38564),
            .I(N__38557));
    InMux I__8586 (
            .O(N__38563),
            .I(N__38553));
    Span4Mux_v I__8585 (
            .O(N__38560),
            .I(N__38549));
    LocalMux I__8584 (
            .O(N__38557),
            .I(N__38546));
    CascadeMux I__8583 (
            .O(N__38556),
            .I(N__38543));
    LocalMux I__8582 (
            .O(N__38553),
            .I(N__38539));
    InMux I__8581 (
            .O(N__38552),
            .I(N__38536));
    Span4Mux_h I__8580 (
            .O(N__38549),
            .I(N__38533));
    Span4Mux_v I__8579 (
            .O(N__38546),
            .I(N__38530));
    InMux I__8578 (
            .O(N__38543),
            .I(N__38527));
    InMux I__8577 (
            .O(N__38542),
            .I(N__38524));
    Span12Mux_h I__8576 (
            .O(N__38539),
            .I(N__38519));
    LocalMux I__8575 (
            .O(N__38536),
            .I(N__38519));
    Odrv4 I__8574 (
            .O(N__38533),
            .I(rand_data_10));
    Odrv4 I__8573 (
            .O(N__38530),
            .I(rand_data_10));
    LocalMux I__8572 (
            .O(N__38527),
            .I(rand_data_10));
    LocalMux I__8571 (
            .O(N__38524),
            .I(rand_data_10));
    Odrv12 I__8570 (
            .O(N__38519),
            .I(rand_data_10));
    CascadeMux I__8569 (
            .O(N__38508),
            .I(N__38504));
    InMux I__8568 (
            .O(N__38507),
            .I(N__38501));
    InMux I__8567 (
            .O(N__38504),
            .I(N__38498));
    LocalMux I__8566 (
            .O(N__38501),
            .I(rand_setpoint_10));
    LocalMux I__8565 (
            .O(N__38498),
            .I(rand_setpoint_10));
    InMux I__8564 (
            .O(N__38493),
            .I(n16587));
    InMux I__8563 (
            .O(N__38490),
            .I(n16588));
    InMux I__8562 (
            .O(N__38487),
            .I(N__38484));
    LocalMux I__8561 (
            .O(N__38484),
            .I(N__38481));
    Span4Mux_h I__8560 (
            .O(N__38481),
            .I(N__38477));
    CascadeMux I__8559 (
            .O(N__38480),
            .I(N__38474));
    Span4Mux_v I__8558 (
            .O(N__38477),
            .I(N__38471));
    InMux I__8557 (
            .O(N__38474),
            .I(N__38468));
    Odrv4 I__8556 (
            .O(N__38471),
            .I(rand_setpoint_12));
    LocalMux I__8555 (
            .O(N__38468),
            .I(rand_setpoint_12));
    InMux I__8554 (
            .O(N__38463),
            .I(n16589));
    InMux I__8553 (
            .O(N__38460),
            .I(N__38454));
    InMux I__8552 (
            .O(N__38459),
            .I(N__38454));
    LocalMux I__8551 (
            .O(N__38454),
            .I(N__38451));
    Span4Mux_v I__8550 (
            .O(N__38451),
            .I(N__38446));
    InMux I__8549 (
            .O(N__38450),
            .I(N__38442));
    InMux I__8548 (
            .O(N__38449),
            .I(N__38438));
    Span4Mux_h I__8547 (
            .O(N__38446),
            .I(N__38435));
    InMux I__8546 (
            .O(N__38445),
            .I(N__38432));
    LocalMux I__8545 (
            .O(N__38442),
            .I(N__38429));
    InMux I__8544 (
            .O(N__38441),
            .I(N__38426));
    LocalMux I__8543 (
            .O(N__38438),
            .I(N__38423));
    Odrv4 I__8542 (
            .O(N__38435),
            .I(rand_data_13));
    LocalMux I__8541 (
            .O(N__38432),
            .I(rand_data_13));
    Odrv12 I__8540 (
            .O(N__38429),
            .I(rand_data_13));
    LocalMux I__8539 (
            .O(N__38426),
            .I(rand_data_13));
    Odrv12 I__8538 (
            .O(N__38423),
            .I(rand_data_13));
    InMux I__8537 (
            .O(N__38412),
            .I(n16590));
    InMux I__8536 (
            .O(N__38409),
            .I(n16575));
    InMux I__8535 (
            .O(N__38406),
            .I(n16576));
    InMux I__8534 (
            .O(N__38403),
            .I(n16577));
    InMux I__8533 (
            .O(N__38400),
            .I(N__38396));
    InMux I__8532 (
            .O(N__38399),
            .I(N__38393));
    LocalMux I__8531 (
            .O(N__38396),
            .I(N__38389));
    LocalMux I__8530 (
            .O(N__38393),
            .I(N__38385));
    InMux I__8529 (
            .O(N__38392),
            .I(N__38382));
    Span4Mux_v I__8528 (
            .O(N__38389),
            .I(N__38378));
    CascadeMux I__8527 (
            .O(N__38388),
            .I(N__38375));
    Span4Mux_v I__8526 (
            .O(N__38385),
            .I(N__38370));
    LocalMux I__8525 (
            .O(N__38382),
            .I(N__38370));
    InMux I__8524 (
            .O(N__38381),
            .I(N__38366));
    Span4Mux_h I__8523 (
            .O(N__38378),
            .I(N__38363));
    InMux I__8522 (
            .O(N__38375),
            .I(N__38360));
    Span4Mux_h I__8521 (
            .O(N__38370),
            .I(N__38357));
    InMux I__8520 (
            .O(N__38369),
            .I(N__38354));
    LocalMux I__8519 (
            .O(N__38366),
            .I(N__38351));
    Odrv4 I__8518 (
            .O(N__38363),
            .I(rand_data_0));
    LocalMux I__8517 (
            .O(N__38360),
            .I(rand_data_0));
    Odrv4 I__8516 (
            .O(N__38357),
            .I(rand_data_0));
    LocalMux I__8515 (
            .O(N__38354),
            .I(rand_data_0));
    Odrv12 I__8514 (
            .O(N__38351),
            .I(rand_data_0));
    InMux I__8513 (
            .O(N__38340),
            .I(N__38337));
    LocalMux I__8512 (
            .O(N__38337),
            .I(N__38332));
    InMux I__8511 (
            .O(N__38336),
            .I(N__38329));
    InMux I__8510 (
            .O(N__38335),
            .I(N__38326));
    Span4Mux_h I__8509 (
            .O(N__38332),
            .I(N__38321));
    LocalMux I__8508 (
            .O(N__38329),
            .I(N__38321));
    LocalMux I__8507 (
            .O(N__38326),
            .I(N__38317));
    Span4Mux_v I__8506 (
            .O(N__38321),
            .I(N__38313));
    CascadeMux I__8505 (
            .O(N__38320),
            .I(N__38310));
    Span4Mux_h I__8504 (
            .O(N__38317),
            .I(N__38306));
    InMux I__8503 (
            .O(N__38316),
            .I(N__38303));
    Sp12to4 I__8502 (
            .O(N__38313),
            .I(N__38300));
    InMux I__8501 (
            .O(N__38310),
            .I(N__38297));
    InMux I__8500 (
            .O(N__38309),
            .I(N__38294));
    Sp12to4 I__8499 (
            .O(N__38306),
            .I(N__38289));
    LocalMux I__8498 (
            .O(N__38303),
            .I(N__38289));
    Odrv12 I__8497 (
            .O(N__38300),
            .I(rand_data_1));
    LocalMux I__8496 (
            .O(N__38297),
            .I(rand_data_1));
    LocalMux I__8495 (
            .O(N__38294),
            .I(rand_data_1));
    Odrv12 I__8494 (
            .O(N__38289),
            .I(rand_data_1));
    InMux I__8493 (
            .O(N__38280),
            .I(n16578));
    InMux I__8492 (
            .O(N__38277),
            .I(N__38272));
    InMux I__8491 (
            .O(N__38276),
            .I(N__38268));
    InMux I__8490 (
            .O(N__38275),
            .I(N__38265));
    LocalMux I__8489 (
            .O(N__38272),
            .I(N__38262));
    InMux I__8488 (
            .O(N__38271),
            .I(N__38258));
    LocalMux I__8487 (
            .O(N__38268),
            .I(N__38255));
    LocalMux I__8486 (
            .O(N__38265),
            .I(N__38252));
    Sp12to4 I__8485 (
            .O(N__38262),
            .I(N__38248));
    InMux I__8484 (
            .O(N__38261),
            .I(N__38245));
    LocalMux I__8483 (
            .O(N__38258),
            .I(N__38242));
    Span4Mux_h I__8482 (
            .O(N__38255),
            .I(N__38239));
    Span4Mux_h I__8481 (
            .O(N__38252),
            .I(N__38236));
    InMux I__8480 (
            .O(N__38251),
            .I(N__38233));
    Span12Mux_h I__8479 (
            .O(N__38248),
            .I(N__38228));
    LocalMux I__8478 (
            .O(N__38245),
            .I(N__38228));
    Odrv12 I__8477 (
            .O(N__38242),
            .I(rand_data_2));
    Odrv4 I__8476 (
            .O(N__38239),
            .I(rand_data_2));
    Odrv4 I__8475 (
            .O(N__38236),
            .I(rand_data_2));
    LocalMux I__8474 (
            .O(N__38233),
            .I(rand_data_2));
    Odrv12 I__8473 (
            .O(N__38228),
            .I(rand_data_2));
    CascadeMux I__8472 (
            .O(N__38217),
            .I(N__38214));
    InMux I__8471 (
            .O(N__38214),
            .I(N__38211));
    LocalMux I__8470 (
            .O(N__38211),
            .I(N__38208));
    Span4Mux_h I__8469 (
            .O(N__38208),
            .I(N__38204));
    CascadeMux I__8468 (
            .O(N__38207),
            .I(N__38201));
    Sp12to4 I__8467 (
            .O(N__38204),
            .I(N__38198));
    InMux I__8466 (
            .O(N__38201),
            .I(N__38195));
    Odrv12 I__8465 (
            .O(N__38198),
            .I(rand_setpoint_2));
    LocalMux I__8464 (
            .O(N__38195),
            .I(rand_setpoint_2));
    InMux I__8463 (
            .O(N__38190),
            .I(n16579));
    InMux I__8462 (
            .O(N__38187),
            .I(N__38183));
    InMux I__8461 (
            .O(N__38186),
            .I(N__38179));
    LocalMux I__8460 (
            .O(N__38183),
            .I(N__38176));
    InMux I__8459 (
            .O(N__38182),
            .I(N__38171));
    LocalMux I__8458 (
            .O(N__38179),
            .I(N__38168));
    Span4Mux_v I__8457 (
            .O(N__38176),
            .I(N__38165));
    InMux I__8456 (
            .O(N__38175),
            .I(N__38161));
    InMux I__8455 (
            .O(N__38174),
            .I(N__38158));
    LocalMux I__8454 (
            .O(N__38171),
            .I(N__38155));
    Span4Mux_h I__8453 (
            .O(N__38168),
            .I(N__38150));
    Span4Mux_v I__8452 (
            .O(N__38165),
            .I(N__38150));
    InMux I__8451 (
            .O(N__38164),
            .I(N__38147));
    LocalMux I__8450 (
            .O(N__38161),
            .I(N__38144));
    LocalMux I__8449 (
            .O(N__38158),
            .I(rand_data_3));
    Odrv4 I__8448 (
            .O(N__38155),
            .I(rand_data_3));
    Odrv4 I__8447 (
            .O(N__38150),
            .I(rand_data_3));
    LocalMux I__8446 (
            .O(N__38147),
            .I(rand_data_3));
    Odrv12 I__8445 (
            .O(N__38144),
            .I(rand_data_3));
    InMux I__8444 (
            .O(N__38133),
            .I(N__38130));
    LocalMux I__8443 (
            .O(N__38130),
            .I(N__38126));
    CascadeMux I__8442 (
            .O(N__38129),
            .I(N__38123));
    Span4Mux_v I__8441 (
            .O(N__38126),
            .I(N__38120));
    InMux I__8440 (
            .O(N__38123),
            .I(N__38117));
    Odrv4 I__8439 (
            .O(N__38120),
            .I(rand_setpoint_3));
    LocalMux I__8438 (
            .O(N__38117),
            .I(rand_setpoint_3));
    InMux I__8437 (
            .O(N__38112),
            .I(n16580));
    InMux I__8436 (
            .O(N__38109),
            .I(N__38104));
    InMux I__8435 (
            .O(N__38108),
            .I(N__38101));
    InMux I__8434 (
            .O(N__38107),
            .I(N__38098));
    LocalMux I__8433 (
            .O(N__38104),
            .I(N__38091));
    LocalMux I__8432 (
            .O(N__38101),
            .I(N__38091));
    LocalMux I__8431 (
            .O(N__38098),
            .I(N__38091));
    Span4Mux_v I__8430 (
            .O(N__38091),
            .I(N__38087));
    CascadeMux I__8429 (
            .O(N__38090),
            .I(N__38084));
    Sp12to4 I__8428 (
            .O(N__38087),
            .I(N__38079));
    InMux I__8427 (
            .O(N__38084),
            .I(N__38076));
    InMux I__8426 (
            .O(N__38083),
            .I(N__38073));
    InMux I__8425 (
            .O(N__38082),
            .I(N__38070));
    Span12Mux_h I__8424 (
            .O(N__38079),
            .I(N__38065));
    LocalMux I__8423 (
            .O(N__38076),
            .I(N__38065));
    LocalMux I__8422 (
            .O(N__38073),
            .I(rand_data_4));
    LocalMux I__8421 (
            .O(N__38070),
            .I(rand_data_4));
    Odrv12 I__8420 (
            .O(N__38065),
            .I(rand_data_4));
    InMux I__8419 (
            .O(N__38058),
            .I(N__38055));
    LocalMux I__8418 (
            .O(N__38055),
            .I(N__38052));
    Span4Mux_h I__8417 (
            .O(N__38052),
            .I(N__38049));
    Span4Mux_v I__8416 (
            .O(N__38049),
            .I(N__38045));
    InMux I__8415 (
            .O(N__38048),
            .I(N__38042));
    Odrv4 I__8414 (
            .O(N__38045),
            .I(rand_setpoint_4));
    LocalMux I__8413 (
            .O(N__38042),
            .I(rand_setpoint_4));
    InMux I__8412 (
            .O(N__38037),
            .I(n16581));
    InMux I__8411 (
            .O(N__38034),
            .I(N__38031));
    LocalMux I__8410 (
            .O(N__38031),
            .I(N__38028));
    Span4Mux_v I__8409 (
            .O(N__38028),
            .I(N__38025));
    Span4Mux_h I__8408 (
            .O(N__38025),
            .I(N__38021));
    InMux I__8407 (
            .O(N__38024),
            .I(N__38018));
    Odrv4 I__8406 (
            .O(N__38021),
            .I(rand_setpoint_5));
    LocalMux I__8405 (
            .O(N__38018),
            .I(rand_setpoint_5));
    InMux I__8404 (
            .O(N__38013),
            .I(n16582));
    InMux I__8403 (
            .O(N__38010),
            .I(n16566));
    InMux I__8402 (
            .O(N__38007),
            .I(n16567));
    InMux I__8401 (
            .O(N__38004),
            .I(n16568));
    InMux I__8400 (
            .O(N__38001),
            .I(n16569));
    InMux I__8399 (
            .O(N__37998),
            .I(bfn_14_8_0_));
    InMux I__8398 (
            .O(N__37995),
            .I(n16571));
    InMux I__8397 (
            .O(N__37992),
            .I(n16572));
    InMux I__8396 (
            .O(N__37989),
            .I(n16573));
    InMux I__8395 (
            .O(N__37986),
            .I(n16574));
    InMux I__8394 (
            .O(N__37983),
            .I(n16557));
    InMux I__8393 (
            .O(N__37980),
            .I(n16558));
    InMux I__8392 (
            .O(N__37977),
            .I(n16559));
    InMux I__8391 (
            .O(N__37974),
            .I(n16560));
    InMux I__8390 (
            .O(N__37971),
            .I(n16561));
    InMux I__8389 (
            .O(N__37968),
            .I(bfn_14_7_0_));
    InMux I__8388 (
            .O(N__37965),
            .I(n16563));
    InMux I__8387 (
            .O(N__37962),
            .I(n16564));
    InMux I__8386 (
            .O(N__37959),
            .I(n16565));
    InMux I__8385 (
            .O(N__37956),
            .I(n16548));
    InMux I__8384 (
            .O(N__37953),
            .I(n16549));
    InMux I__8383 (
            .O(N__37950),
            .I(n16550));
    InMux I__8382 (
            .O(N__37947),
            .I(n16551));
    InMux I__8381 (
            .O(N__37944),
            .I(n16552));
    InMux I__8380 (
            .O(N__37941),
            .I(n16553));
    InMux I__8379 (
            .O(N__37938),
            .I(bfn_14_6_0_));
    InMux I__8378 (
            .O(N__37935),
            .I(n16555));
    InMux I__8377 (
            .O(N__37932),
            .I(n16556));
    InMux I__8376 (
            .O(N__37929),
            .I(N__37926));
    LocalMux I__8375 (
            .O(N__37926),
            .I(N__37923));
    Span4Mux_s2_v I__8374 (
            .O(N__37923),
            .I(N__37920));
    Span4Mux_h I__8373 (
            .O(N__37920),
            .I(N__37917));
    Odrv4 I__8372 (
            .O(N__37917),
            .I(\c0.n18681 ));
    InMux I__8371 (
            .O(N__37914),
            .I(bfn_14_5_0_));
    InMux I__8370 (
            .O(N__37911),
            .I(n16547));
    InMux I__8369 (
            .O(N__37908),
            .I(N__37905));
    LocalMux I__8368 (
            .O(N__37905),
            .I(\c0.n17783 ));
    CascadeMux I__8367 (
            .O(N__37902),
            .I(\c0.n15_adj_2414_cascade_ ));
    InMux I__8366 (
            .O(N__37899),
            .I(N__37896));
    LocalMux I__8365 (
            .O(N__37896),
            .I(N__37893));
    Span4Mux_s1_v I__8364 (
            .O(N__37893),
            .I(N__37890));
    Odrv4 I__8363 (
            .O(N__37890),
            .I(\c0.data_out_frame2_20_1 ));
    InMux I__8362 (
            .O(N__37887),
            .I(N__37884));
    LocalMux I__8361 (
            .O(N__37884),
            .I(N__37881));
    Span4Mux_v I__8360 (
            .O(N__37881),
            .I(N__37878));
    Odrv4 I__8359 (
            .O(N__37878),
            .I(\c0.n31 ));
    CascadeMux I__8358 (
            .O(N__37875),
            .I(\c0.n32_cascade_ ));
    InMux I__8357 (
            .O(N__37872),
            .I(N__37869));
    LocalMux I__8356 (
            .O(N__37869),
            .I(N__37866));
    Span12Mux_s2_v I__8355 (
            .O(N__37866),
            .I(N__37863));
    Odrv12 I__8354 (
            .O(N__37863),
            .I(\c0.data_out_frame2_19_7 ));
    InMux I__8353 (
            .O(N__37860),
            .I(N__37855));
    InMux I__8352 (
            .O(N__37859),
            .I(N__37850));
    InMux I__8351 (
            .O(N__37858),
            .I(N__37850));
    LocalMux I__8350 (
            .O(N__37855),
            .I(N__37847));
    LocalMux I__8349 (
            .O(N__37850),
            .I(N__37844));
    Span4Mux_s2_v I__8348 (
            .O(N__37847),
            .I(N__37839));
    Span4Mux_h I__8347 (
            .O(N__37844),
            .I(N__37836));
    InMux I__8346 (
            .O(N__37843),
            .I(N__37831));
    InMux I__8345 (
            .O(N__37842),
            .I(N__37831));
    Span4Mux_h I__8344 (
            .O(N__37839),
            .I(N__37828));
    Odrv4 I__8343 (
            .O(N__37836),
            .I(\c0.data_out_frame2_0_7 ));
    LocalMux I__8342 (
            .O(N__37831),
            .I(\c0.data_out_frame2_0_7 ));
    Odrv4 I__8341 (
            .O(N__37828),
            .I(\c0.data_out_frame2_0_7 ));
    InMux I__8340 (
            .O(N__37821),
            .I(N__37818));
    LocalMux I__8339 (
            .O(N__37818),
            .I(N__37815));
    Odrv12 I__8338 (
            .O(N__37815),
            .I(\c0.n17777 ));
    InMux I__8337 (
            .O(N__37812),
            .I(N__37809));
    LocalMux I__8336 (
            .O(N__37809),
            .I(\c0.n6_adj_2430 ));
    CascadeMux I__8335 (
            .O(N__37806),
            .I(\c0.n17777_cascade_ ));
    InMux I__8334 (
            .O(N__37803),
            .I(N__37799));
    InMux I__8333 (
            .O(N__37802),
            .I(N__37796));
    LocalMux I__8332 (
            .O(N__37799),
            .I(N__37793));
    LocalMux I__8331 (
            .O(N__37796),
            .I(N__37789));
    Span4Mux_s3_v I__8330 (
            .O(N__37793),
            .I(N__37786));
    CascadeMux I__8329 (
            .O(N__37792),
            .I(N__37782));
    Span4Mux_h I__8328 (
            .O(N__37789),
            .I(N__37779));
    Span4Mux_h I__8327 (
            .O(N__37786),
            .I(N__37776));
    InMux I__8326 (
            .O(N__37785),
            .I(N__37771));
    InMux I__8325 (
            .O(N__37782),
            .I(N__37771));
    Odrv4 I__8324 (
            .O(N__37779),
            .I(data_out_frame2_5_5));
    Odrv4 I__8323 (
            .O(N__37776),
            .I(data_out_frame2_5_5));
    LocalMux I__8322 (
            .O(N__37771),
            .I(data_out_frame2_5_5));
    CascadeMux I__8321 (
            .O(N__37764),
            .I(\c0.n10617_cascade_ ));
    InMux I__8320 (
            .O(N__37761),
            .I(N__37758));
    LocalMux I__8319 (
            .O(N__37758),
            .I(N__37755));
    Span4Mux_s2_v I__8318 (
            .O(N__37755),
            .I(N__37751));
    InMux I__8317 (
            .O(N__37754),
            .I(N__37748));
    Odrv4 I__8316 (
            .O(N__37751),
            .I(\c0.n17765 ));
    LocalMux I__8315 (
            .O(N__37748),
            .I(\c0.n17765 ));
    InMux I__8314 (
            .O(N__37743),
            .I(N__37737));
    InMux I__8313 (
            .O(N__37742),
            .I(N__37734));
    CascadeMux I__8312 (
            .O(N__37741),
            .I(N__37731));
    InMux I__8311 (
            .O(N__37740),
            .I(N__37728));
    LocalMux I__8310 (
            .O(N__37737),
            .I(N__37725));
    LocalMux I__8309 (
            .O(N__37734),
            .I(N__37722));
    InMux I__8308 (
            .O(N__37731),
            .I(N__37718));
    LocalMux I__8307 (
            .O(N__37728),
            .I(N__37715));
    Span4Mux_s2_v I__8306 (
            .O(N__37725),
            .I(N__37710));
    Span4Mux_h I__8305 (
            .O(N__37722),
            .I(N__37710));
    InMux I__8304 (
            .O(N__37721),
            .I(N__37707));
    LocalMux I__8303 (
            .O(N__37718),
            .I(N__37702));
    Span4Mux_h I__8302 (
            .O(N__37715),
            .I(N__37702));
    Span4Mux_h I__8301 (
            .O(N__37710),
            .I(N__37699));
    LocalMux I__8300 (
            .O(N__37707),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv4 I__8299 (
            .O(N__37702),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv4 I__8298 (
            .O(N__37699),
            .I(\c0.data_out_frame2_0_4 ));
    CascadeMux I__8297 (
            .O(N__37692),
            .I(\c0.n18759_cascade_ ));
    CascadeMux I__8296 (
            .O(N__37689),
            .I(N__37686));
    InMux I__8295 (
            .O(N__37686),
            .I(N__37683));
    LocalMux I__8294 (
            .O(N__37683),
            .I(N__37680));
    Span4Mux_s0_v I__8293 (
            .O(N__37680),
            .I(N__37676));
    CascadeMux I__8292 (
            .O(N__37679),
            .I(N__37672));
    Span4Mux_v I__8291 (
            .O(N__37676),
            .I(N__37668));
    InMux I__8290 (
            .O(N__37675),
            .I(N__37663));
    InMux I__8289 (
            .O(N__37672),
            .I(N__37663));
    InMux I__8288 (
            .O(N__37671),
            .I(N__37660));
    Odrv4 I__8287 (
            .O(N__37668),
            .I(data_out_frame2_6_0));
    LocalMux I__8286 (
            .O(N__37663),
            .I(data_out_frame2_6_0));
    LocalMux I__8285 (
            .O(N__37660),
            .I(data_out_frame2_6_0));
    InMux I__8284 (
            .O(N__37653),
            .I(N__37650));
    LocalMux I__8283 (
            .O(N__37650),
            .I(N__37647));
    Odrv12 I__8282 (
            .O(N__37647),
            .I(\c0.n10920 ));
    CascadeMux I__8281 (
            .O(N__37644),
            .I(\c0.n17783_cascade_ ));
    InMux I__8280 (
            .O(N__37641),
            .I(N__37638));
    LocalMux I__8279 (
            .O(N__37638),
            .I(N__37634));
    InMux I__8278 (
            .O(N__37637),
            .I(N__37631));
    Odrv4 I__8277 (
            .O(N__37634),
            .I(\c0.n10849 ));
    LocalMux I__8276 (
            .O(N__37631),
            .I(\c0.n10849 ));
    InMux I__8275 (
            .O(N__37626),
            .I(N__37623));
    LocalMux I__8274 (
            .O(N__37623),
            .I(N__37619));
    CascadeMux I__8273 (
            .O(N__37622),
            .I(N__37616));
    Span4Mux_s1_v I__8272 (
            .O(N__37619),
            .I(N__37613));
    InMux I__8271 (
            .O(N__37616),
            .I(N__37610));
    Odrv4 I__8270 (
            .O(N__37613),
            .I(\c0.n17859 ));
    LocalMux I__8269 (
            .O(N__37610),
            .I(\c0.n17859 ));
    CascadeMux I__8268 (
            .O(N__37605),
            .I(\c0.n15_cascade_ ));
    CascadeMux I__8267 (
            .O(N__37602),
            .I(N__37599));
    InMux I__8266 (
            .O(N__37599),
            .I(N__37596));
    LocalMux I__8265 (
            .O(N__37596),
            .I(N__37593));
    Span4Mux_v I__8264 (
            .O(N__37593),
            .I(N__37590));
    Odrv4 I__8263 (
            .O(N__37590),
            .I(\c0.data_out_frame2_19_0 ));
    InMux I__8262 (
            .O(N__37587),
            .I(N__37584));
    LocalMux I__8261 (
            .O(N__37584),
            .I(N__37580));
    CascadeMux I__8260 (
            .O(N__37583),
            .I(N__37577));
    Sp12to4 I__8259 (
            .O(N__37580),
            .I(N__37574));
    InMux I__8258 (
            .O(N__37577),
            .I(N__37571));
    Span12Mux_s2_v I__8257 (
            .O(N__37574),
            .I(N__37566));
    LocalMux I__8256 (
            .O(N__37571),
            .I(N__37566));
    Odrv12 I__8255 (
            .O(N__37566),
            .I(\c0.n10688 ));
    CascadeMux I__8254 (
            .O(N__37563),
            .I(\c0.n10813_cascade_ ));
    InMux I__8253 (
            .O(N__37560),
            .I(N__37556));
    InMux I__8252 (
            .O(N__37559),
            .I(N__37553));
    LocalMux I__8251 (
            .O(N__37556),
            .I(N__37550));
    LocalMux I__8250 (
            .O(N__37553),
            .I(\c0.n10577 ));
    Odrv4 I__8249 (
            .O(N__37550),
            .I(\c0.n10577 ));
    InMux I__8248 (
            .O(N__37545),
            .I(N__37541));
    InMux I__8247 (
            .O(N__37544),
            .I(N__37538));
    LocalMux I__8246 (
            .O(N__37541),
            .I(N__37529));
    LocalMux I__8245 (
            .O(N__37538),
            .I(N__37529));
    InMux I__8244 (
            .O(N__37537),
            .I(N__37526));
    InMux I__8243 (
            .O(N__37536),
            .I(N__37523));
    InMux I__8242 (
            .O(N__37535),
            .I(N__37518));
    InMux I__8241 (
            .O(N__37534),
            .I(N__37518));
    Span4Mux_v I__8240 (
            .O(N__37529),
            .I(N__37515));
    LocalMux I__8239 (
            .O(N__37526),
            .I(N__37512));
    LocalMux I__8238 (
            .O(N__37523),
            .I(data_out_6_0));
    LocalMux I__8237 (
            .O(N__37518),
            .I(data_out_6_0));
    Odrv4 I__8236 (
            .O(N__37515),
            .I(data_out_6_0));
    Odrv4 I__8235 (
            .O(N__37512),
            .I(data_out_6_0));
    CascadeMux I__8234 (
            .O(N__37503),
            .I(N__37500));
    InMux I__8233 (
            .O(N__37500),
            .I(N__37497));
    LocalMux I__8232 (
            .O(N__37497),
            .I(\c0.n10680 ));
    InMux I__8231 (
            .O(N__37494),
            .I(N__37491));
    LocalMux I__8230 (
            .O(N__37491),
            .I(\c0.n17816 ));
    CascadeMux I__8229 (
            .O(N__37488),
            .I(\c0.n10680_cascade_ ));
    InMux I__8228 (
            .O(N__37485),
            .I(N__37479));
    InMux I__8227 (
            .O(N__37484),
            .I(N__37476));
    InMux I__8226 (
            .O(N__37483),
            .I(N__37473));
    InMux I__8225 (
            .O(N__37482),
            .I(N__37470));
    LocalMux I__8224 (
            .O(N__37479),
            .I(N__37464));
    LocalMux I__8223 (
            .O(N__37476),
            .I(N__37464));
    LocalMux I__8222 (
            .O(N__37473),
            .I(N__37461));
    LocalMux I__8221 (
            .O(N__37470),
            .I(N__37458));
    InMux I__8220 (
            .O(N__37469),
            .I(N__37455));
    Span4Mux_v I__8219 (
            .O(N__37464),
            .I(N__37452));
    Odrv4 I__8218 (
            .O(N__37461),
            .I(\c0.data_out_5_5 ));
    Odrv4 I__8217 (
            .O(N__37458),
            .I(\c0.data_out_5_5 ));
    LocalMux I__8216 (
            .O(N__37455),
            .I(\c0.data_out_5_5 ));
    Odrv4 I__8215 (
            .O(N__37452),
            .I(\c0.data_out_5_5 ));
    InMux I__8214 (
            .O(N__37443),
            .I(N__37438));
    InMux I__8213 (
            .O(N__37442),
            .I(N__37435));
    InMux I__8212 (
            .O(N__37441),
            .I(N__37430));
    LocalMux I__8211 (
            .O(N__37438),
            .I(N__37427));
    LocalMux I__8210 (
            .O(N__37435),
            .I(N__37424));
    InMux I__8209 (
            .O(N__37434),
            .I(N__37419));
    InMux I__8208 (
            .O(N__37433),
            .I(N__37419));
    LocalMux I__8207 (
            .O(N__37430),
            .I(N__37412));
    Span4Mux_v I__8206 (
            .O(N__37427),
            .I(N__37412));
    Span4Mux_v I__8205 (
            .O(N__37424),
            .I(N__37412));
    LocalMux I__8204 (
            .O(N__37419),
            .I(data_out_8_6));
    Odrv4 I__8203 (
            .O(N__37412),
            .I(data_out_8_6));
    InMux I__8202 (
            .O(N__37407),
            .I(N__37404));
    LocalMux I__8201 (
            .O(N__37404),
            .I(N__37400));
    InMux I__8200 (
            .O(N__37403),
            .I(N__37397));
    Span4Mux_v I__8199 (
            .O(N__37400),
            .I(N__37394));
    LocalMux I__8198 (
            .O(N__37397),
            .I(N__37391));
    Span4Mux_h I__8197 (
            .O(N__37394),
            .I(N__37383));
    Span4Mux_v I__8196 (
            .O(N__37391),
            .I(N__37383));
    InMux I__8195 (
            .O(N__37390),
            .I(N__37378));
    InMux I__8194 (
            .O(N__37389),
            .I(N__37378));
    InMux I__8193 (
            .O(N__37388),
            .I(N__37375));
    Odrv4 I__8192 (
            .O(N__37383),
            .I(data_out_8_5));
    LocalMux I__8191 (
            .O(N__37378),
            .I(data_out_8_5));
    LocalMux I__8190 (
            .O(N__37375),
            .I(data_out_8_5));
    CascadeMux I__8189 (
            .O(N__37368),
            .I(N__37365));
    InMux I__8188 (
            .O(N__37365),
            .I(N__37362));
    LocalMux I__8187 (
            .O(N__37362),
            .I(N__37358));
    InMux I__8186 (
            .O(N__37361),
            .I(N__37355));
    Span4Mux_v I__8185 (
            .O(N__37358),
            .I(N__37352));
    LocalMux I__8184 (
            .O(N__37355),
            .I(N__37349));
    Span4Mux_v I__8183 (
            .O(N__37352),
            .I(N__37346));
    Odrv4 I__8182 (
            .O(N__37349),
            .I(\c0.n17771 ));
    Odrv4 I__8181 (
            .O(N__37346),
            .I(\c0.n17771 ));
    InMux I__8180 (
            .O(N__37341),
            .I(N__37337));
    InMux I__8179 (
            .O(N__37340),
            .I(N__37332));
    LocalMux I__8178 (
            .O(N__37337),
            .I(N__37329));
    InMux I__8177 (
            .O(N__37336),
            .I(N__37326));
    InMux I__8176 (
            .O(N__37335),
            .I(N__37323));
    LocalMux I__8175 (
            .O(N__37332),
            .I(N__37320));
    Span4Mux_v I__8174 (
            .O(N__37329),
            .I(N__37317));
    LocalMux I__8173 (
            .O(N__37326),
            .I(N__37314));
    LocalMux I__8172 (
            .O(N__37323),
            .I(N__37310));
    Span4Mux_v I__8171 (
            .O(N__37320),
            .I(N__37307));
    Span4Mux_v I__8170 (
            .O(N__37317),
            .I(N__37304));
    Span4Mux_h I__8169 (
            .O(N__37314),
            .I(N__37301));
    InMux I__8168 (
            .O(N__37313),
            .I(N__37298));
    Span4Mux_h I__8167 (
            .O(N__37310),
            .I(N__37295));
    Odrv4 I__8166 (
            .O(N__37307),
            .I(data_out_5_1));
    Odrv4 I__8165 (
            .O(N__37304),
            .I(data_out_5_1));
    Odrv4 I__8164 (
            .O(N__37301),
            .I(data_out_5_1));
    LocalMux I__8163 (
            .O(N__37298),
            .I(data_out_5_1));
    Odrv4 I__8162 (
            .O(N__37295),
            .I(data_out_5_1));
    InMux I__8161 (
            .O(N__37284),
            .I(N__37279));
    InMux I__8160 (
            .O(N__37283),
            .I(N__37272));
    InMux I__8159 (
            .O(N__37282),
            .I(N__37269));
    LocalMux I__8158 (
            .O(N__37279),
            .I(N__37266));
    InMux I__8157 (
            .O(N__37278),
            .I(N__37261));
    InMux I__8156 (
            .O(N__37277),
            .I(N__37261));
    InMux I__8155 (
            .O(N__37276),
            .I(N__37256));
    InMux I__8154 (
            .O(N__37275),
            .I(N__37256));
    LocalMux I__8153 (
            .O(N__37272),
            .I(N__37253));
    LocalMux I__8152 (
            .O(N__37269),
            .I(N__37250));
    Span4Mux_v I__8151 (
            .O(N__37266),
            .I(N__37246));
    LocalMux I__8150 (
            .O(N__37261),
            .I(N__37243));
    LocalMux I__8149 (
            .O(N__37256),
            .I(N__37240));
    Span4Mux_v I__8148 (
            .O(N__37253),
            .I(N__37235));
    Span4Mux_h I__8147 (
            .O(N__37250),
            .I(N__37235));
    InMux I__8146 (
            .O(N__37249),
            .I(N__37232));
    Odrv4 I__8145 (
            .O(N__37246),
            .I(\c0.data_out_5_4 ));
    Odrv12 I__8144 (
            .O(N__37243),
            .I(\c0.data_out_5_4 ));
    Odrv4 I__8143 (
            .O(N__37240),
            .I(\c0.data_out_5_4 ));
    Odrv4 I__8142 (
            .O(N__37235),
            .I(\c0.data_out_5_4 ));
    LocalMux I__8141 (
            .O(N__37232),
            .I(\c0.data_out_5_4 ));
    InMux I__8140 (
            .O(N__37221),
            .I(N__37217));
    InMux I__8139 (
            .O(N__37220),
            .I(N__37214));
    LocalMux I__8138 (
            .O(N__37217),
            .I(N__37209));
    LocalMux I__8137 (
            .O(N__37214),
            .I(N__37206));
    InMux I__8136 (
            .O(N__37213),
            .I(N__37203));
    InMux I__8135 (
            .O(N__37212),
            .I(N__37200));
    Span12Mux_h I__8134 (
            .O(N__37209),
            .I(N__37193));
    Span12Mux_h I__8133 (
            .O(N__37206),
            .I(N__37193));
    LocalMux I__8132 (
            .O(N__37203),
            .I(N__37193));
    LocalMux I__8131 (
            .O(N__37200),
            .I(data_out_frame2_13_2));
    Odrv12 I__8130 (
            .O(N__37193),
            .I(data_out_frame2_13_2));
    InMux I__8129 (
            .O(N__37188),
            .I(N__37184));
    InMux I__8128 (
            .O(N__37187),
            .I(N__37180));
    LocalMux I__8127 (
            .O(N__37184),
            .I(N__37175));
    InMux I__8126 (
            .O(N__37183),
            .I(N__37172));
    LocalMux I__8125 (
            .O(N__37180),
            .I(N__37169));
    InMux I__8124 (
            .O(N__37179),
            .I(N__37166));
    InMux I__8123 (
            .O(N__37178),
            .I(N__37163));
    Span4Mux_h I__8122 (
            .O(N__37175),
            .I(N__37160));
    LocalMux I__8121 (
            .O(N__37172),
            .I(N__37157));
    Span4Mux_s0_v I__8120 (
            .O(N__37169),
            .I(N__37154));
    LocalMux I__8119 (
            .O(N__37166),
            .I(N__37151));
    LocalMux I__8118 (
            .O(N__37163),
            .I(data_out_frame2_16_0));
    Odrv4 I__8117 (
            .O(N__37160),
            .I(data_out_frame2_16_0));
    Odrv4 I__8116 (
            .O(N__37157),
            .I(data_out_frame2_16_0));
    Odrv4 I__8115 (
            .O(N__37154),
            .I(data_out_frame2_16_0));
    Odrv12 I__8114 (
            .O(N__37151),
            .I(data_out_frame2_16_0));
    InMux I__8113 (
            .O(N__37140),
            .I(N__37135));
    InMux I__8112 (
            .O(N__37139),
            .I(N__37130));
    InMux I__8111 (
            .O(N__37138),
            .I(N__37130));
    LocalMux I__8110 (
            .O(N__37135),
            .I(N__37125));
    LocalMux I__8109 (
            .O(N__37130),
            .I(N__37122));
    InMux I__8108 (
            .O(N__37129),
            .I(N__37119));
    InMux I__8107 (
            .O(N__37128),
            .I(N__37116));
    Span4Mux_h I__8106 (
            .O(N__37125),
            .I(N__37113));
    Span4Mux_h I__8105 (
            .O(N__37122),
            .I(N__37110));
    LocalMux I__8104 (
            .O(N__37119),
            .I(data_out_frame2_8_6));
    LocalMux I__8103 (
            .O(N__37116),
            .I(data_out_frame2_8_6));
    Odrv4 I__8102 (
            .O(N__37113),
            .I(data_out_frame2_8_6));
    Odrv4 I__8101 (
            .O(N__37110),
            .I(data_out_frame2_8_6));
    InMux I__8100 (
            .O(N__37101),
            .I(N__37098));
    LocalMux I__8099 (
            .O(N__37098),
            .I(N__37094));
    InMux I__8098 (
            .O(N__37097),
            .I(N__37089));
    Span4Mux_h I__8097 (
            .O(N__37094),
            .I(N__37086));
    InMux I__8096 (
            .O(N__37093),
            .I(N__37083));
    InMux I__8095 (
            .O(N__37092),
            .I(N__37080));
    LocalMux I__8094 (
            .O(N__37089),
            .I(data_out_10_6));
    Odrv4 I__8093 (
            .O(N__37086),
            .I(data_out_10_6));
    LocalMux I__8092 (
            .O(N__37083),
            .I(data_out_10_6));
    LocalMux I__8091 (
            .O(N__37080),
            .I(data_out_10_6));
    InMux I__8090 (
            .O(N__37071),
            .I(N__37067));
    InMux I__8089 (
            .O(N__37070),
            .I(N__37063));
    LocalMux I__8088 (
            .O(N__37067),
            .I(N__37060));
    InMux I__8087 (
            .O(N__37066),
            .I(N__37057));
    LocalMux I__8086 (
            .O(N__37063),
            .I(N__37052));
    Span4Mux_v I__8085 (
            .O(N__37060),
            .I(N__37052));
    LocalMux I__8084 (
            .O(N__37057),
            .I(\c0.data_out_7_2 ));
    Odrv4 I__8083 (
            .O(N__37052),
            .I(\c0.data_out_7_2 ));
    CascadeMux I__8082 (
            .O(N__37047),
            .I(N__37044));
    InMux I__8081 (
            .O(N__37044),
            .I(N__37040));
    InMux I__8080 (
            .O(N__37043),
            .I(N__37037));
    LocalMux I__8079 (
            .O(N__37040),
            .I(N__37031));
    LocalMux I__8078 (
            .O(N__37037),
            .I(N__37031));
    CascadeMux I__8077 (
            .O(N__37036),
            .I(N__37028));
    Span4Mux_v I__8076 (
            .O(N__37031),
            .I(N__37025));
    InMux I__8075 (
            .O(N__37028),
            .I(N__37022));
    Odrv4 I__8074 (
            .O(N__37025),
            .I(\c0.data_out_9_1 ));
    LocalMux I__8073 (
            .O(N__37022),
            .I(\c0.data_out_9_1 ));
    InMux I__8072 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__8071 (
            .O(N__37014),
            .I(N__37011));
    Span4Mux_h I__8070 (
            .O(N__37011),
            .I(N__37008));
    Odrv4 I__8069 (
            .O(N__37008),
            .I(\c0.n17730 ));
    InMux I__8068 (
            .O(N__37005),
            .I(N__37001));
    InMux I__8067 (
            .O(N__37004),
            .I(N__36998));
    LocalMux I__8066 (
            .O(N__37001),
            .I(\c0.n17835 ));
    LocalMux I__8065 (
            .O(N__36998),
            .I(\c0.n17835 ));
    InMux I__8064 (
            .O(N__36993),
            .I(N__36990));
    LocalMux I__8063 (
            .O(N__36990),
            .I(N__36986));
    InMux I__8062 (
            .O(N__36989),
            .I(N__36983));
    Span12Mux_v I__8061 (
            .O(N__36986),
            .I(N__36980));
    LocalMux I__8060 (
            .O(N__36983),
            .I(N__36977));
    Odrv12 I__8059 (
            .O(N__36980),
            .I(\c0.n17844 ));
    Odrv4 I__8058 (
            .O(N__36977),
            .I(\c0.n17844 ));
    CascadeMux I__8057 (
            .O(N__36972),
            .I(\c0.n17730_cascade_ ));
    InMux I__8056 (
            .O(N__36969),
            .I(N__36965));
    InMux I__8055 (
            .O(N__36968),
            .I(N__36962));
    LocalMux I__8054 (
            .O(N__36965),
            .I(N__36959));
    LocalMux I__8053 (
            .O(N__36962),
            .I(n17758));
    Odrv4 I__8052 (
            .O(N__36959),
            .I(n17758));
    CascadeMux I__8051 (
            .O(N__36954),
            .I(\c0.n14_adj_2363_cascade_ ));
    InMux I__8050 (
            .O(N__36951),
            .I(N__36948));
    LocalMux I__8049 (
            .O(N__36948),
            .I(N__36945));
    Odrv4 I__8048 (
            .O(N__36945),
            .I(\c0.n13 ));
    InMux I__8047 (
            .O(N__36942),
            .I(N__36939));
    LocalMux I__8046 (
            .O(N__36939),
            .I(N__36934));
    InMux I__8045 (
            .O(N__36938),
            .I(N__36930));
    InMux I__8044 (
            .O(N__36937),
            .I(N__36927));
    Span4Mux_h I__8043 (
            .O(N__36934),
            .I(N__36924));
    InMux I__8042 (
            .O(N__36933),
            .I(N__36921));
    LocalMux I__8041 (
            .O(N__36930),
            .I(\c0.data_out_9_3 ));
    LocalMux I__8040 (
            .O(N__36927),
            .I(\c0.data_out_9_3 ));
    Odrv4 I__8039 (
            .O(N__36924),
            .I(\c0.data_out_9_3 ));
    LocalMux I__8038 (
            .O(N__36921),
            .I(\c0.data_out_9_3 ));
    CascadeMux I__8037 (
            .O(N__36912),
            .I(\c0.n17816_cascade_ ));
    InMux I__8036 (
            .O(N__36909),
            .I(N__36905));
    InMux I__8035 (
            .O(N__36908),
            .I(N__36902));
    LocalMux I__8034 (
            .O(N__36905),
            .I(\c0.n17877 ));
    LocalMux I__8033 (
            .O(N__36902),
            .I(\c0.n17877 ));
    InMux I__8032 (
            .O(N__36897),
            .I(N__36894));
    LocalMux I__8031 (
            .O(N__36894),
            .I(\c0.n12 ));
    InMux I__8030 (
            .O(N__36891),
            .I(N__36887));
    InMux I__8029 (
            .O(N__36890),
            .I(N__36884));
    LocalMux I__8028 (
            .O(N__36887),
            .I(N__36881));
    LocalMux I__8027 (
            .O(N__36884),
            .I(N__36878));
    Span4Mux_h I__8026 (
            .O(N__36881),
            .I(N__36875));
    Odrv4 I__8025 (
            .O(N__36878),
            .I(\c0.n17786 ));
    Odrv4 I__8024 (
            .O(N__36875),
            .I(\c0.n17786 ));
    InMux I__8023 (
            .O(N__36870),
            .I(N__36867));
    LocalMux I__8022 (
            .O(N__36867),
            .I(N__36864));
    Span4Mux_h I__8021 (
            .O(N__36864),
            .I(N__36861));
    Odrv4 I__8020 (
            .O(N__36861),
            .I(\c0.n18184 ));
    InMux I__8019 (
            .O(N__36858),
            .I(N__36855));
    LocalMux I__8018 (
            .O(N__36855),
            .I(N__36850));
    InMux I__8017 (
            .O(N__36854),
            .I(N__36847));
    InMux I__8016 (
            .O(N__36853),
            .I(N__36844));
    Span4Mux_h I__8015 (
            .O(N__36850),
            .I(N__36841));
    LocalMux I__8014 (
            .O(N__36847),
            .I(N__36838));
    LocalMux I__8013 (
            .O(N__36844),
            .I(\c0.data_out_7_1 ));
    Odrv4 I__8012 (
            .O(N__36841),
            .I(\c0.data_out_7_1 ));
    Odrv4 I__8011 (
            .O(N__36838),
            .I(\c0.data_out_7_1 ));
    InMux I__8010 (
            .O(N__36831),
            .I(N__36824));
    InMux I__8009 (
            .O(N__36830),
            .I(N__36824));
    InMux I__8008 (
            .O(N__36829),
            .I(N__36821));
    LocalMux I__8007 (
            .O(N__36824),
            .I(N__36818));
    LocalMux I__8006 (
            .O(N__36821),
            .I(N__36815));
    Odrv4 I__8005 (
            .O(N__36818),
            .I(\c0.n10537 ));
    Odrv4 I__8004 (
            .O(N__36815),
            .I(\c0.n10537 ));
    CascadeMux I__8003 (
            .O(N__36810),
            .I(\c0.n18238_cascade_ ));
    InMux I__8002 (
            .O(N__36807),
            .I(N__36804));
    LocalMux I__8001 (
            .O(N__36804),
            .I(N__36799));
    InMux I__8000 (
            .O(N__36803),
            .I(N__36794));
    InMux I__7999 (
            .O(N__36802),
            .I(N__36794));
    Span4Mux_v I__7998 (
            .O(N__36799),
            .I(N__36791));
    LocalMux I__7997 (
            .O(N__36794),
            .I(\c0.data_out_6_4 ));
    Odrv4 I__7996 (
            .O(N__36791),
            .I(\c0.data_out_6_4 ));
    InMux I__7995 (
            .O(N__36786),
            .I(N__36783));
    LocalMux I__7994 (
            .O(N__36783),
            .I(N__36780));
    Odrv4 I__7993 (
            .O(N__36780),
            .I(\c0.n6_adj_2276 ));
    InMux I__7992 (
            .O(N__36777),
            .I(N__36773));
    InMux I__7991 (
            .O(N__36776),
            .I(N__36770));
    LocalMux I__7990 (
            .O(N__36773),
            .I(N__36766));
    LocalMux I__7989 (
            .O(N__36770),
            .I(N__36763));
    InMux I__7988 (
            .O(N__36769),
            .I(N__36760));
    Span4Mux_h I__7987 (
            .O(N__36766),
            .I(N__36757));
    Span12Mux_v I__7986 (
            .O(N__36763),
            .I(N__36754));
    LocalMux I__7985 (
            .O(N__36760),
            .I(\c0.data_out_6_7 ));
    Odrv4 I__7984 (
            .O(N__36757),
            .I(\c0.data_out_6_7 ));
    Odrv12 I__7983 (
            .O(N__36754),
            .I(\c0.data_out_6_7 ));
    InMux I__7982 (
            .O(N__36747),
            .I(N__36742));
    InMux I__7981 (
            .O(N__36746),
            .I(N__36739));
    InMux I__7980 (
            .O(N__36745),
            .I(N__36736));
    LocalMux I__7979 (
            .O(N__36742),
            .I(N__36728));
    LocalMux I__7978 (
            .O(N__36739),
            .I(N__36728));
    LocalMux I__7977 (
            .O(N__36736),
            .I(N__36728));
    InMux I__7976 (
            .O(N__36735),
            .I(N__36725));
    Span4Mux_h I__7975 (
            .O(N__36728),
            .I(N__36722));
    LocalMux I__7974 (
            .O(N__36725),
            .I(\c0.data_out_6_5 ));
    Odrv4 I__7973 (
            .O(N__36722),
            .I(\c0.data_out_6_5 ));
    InMux I__7972 (
            .O(N__36717),
            .I(N__36713));
    InMux I__7971 (
            .O(N__36716),
            .I(N__36710));
    LocalMux I__7970 (
            .O(N__36713),
            .I(N__36705));
    LocalMux I__7969 (
            .O(N__36710),
            .I(N__36702));
    InMux I__7968 (
            .O(N__36709),
            .I(N__36699));
    InMux I__7967 (
            .O(N__36708),
            .I(N__36696));
    Span4Mux_v I__7966 (
            .O(N__36705),
            .I(N__36689));
    Span4Mux_v I__7965 (
            .O(N__36702),
            .I(N__36689));
    LocalMux I__7964 (
            .O(N__36699),
            .I(N__36689));
    LocalMux I__7963 (
            .O(N__36696),
            .I(data_out_8_4));
    Odrv4 I__7962 (
            .O(N__36689),
            .I(data_out_8_4));
    CascadeMux I__7961 (
            .O(N__36684),
            .I(N__36681));
    InMux I__7960 (
            .O(N__36681),
            .I(N__36678));
    LocalMux I__7959 (
            .O(N__36678),
            .I(\c0.n17745 ));
    InMux I__7958 (
            .O(N__36675),
            .I(N__36672));
    LocalMux I__7957 (
            .O(N__36672),
            .I(N__36669));
    Odrv4 I__7956 (
            .O(N__36669),
            .I(\c0.n10542 ));
    CascadeMux I__7955 (
            .O(N__36666),
            .I(\c0.n17745_cascade_ ));
    CascadeMux I__7954 (
            .O(N__36663),
            .I(N__36660));
    InMux I__7953 (
            .O(N__36660),
            .I(N__36656));
    CascadeMux I__7952 (
            .O(N__36659),
            .I(N__36653));
    LocalMux I__7951 (
            .O(N__36656),
            .I(N__36650));
    InMux I__7950 (
            .O(N__36653),
            .I(N__36647));
    Span4Mux_h I__7949 (
            .O(N__36650),
            .I(N__36641));
    LocalMux I__7948 (
            .O(N__36647),
            .I(N__36641));
    InMux I__7947 (
            .O(N__36646),
            .I(N__36638));
    Span4Mux_h I__7946 (
            .O(N__36641),
            .I(N__36635));
    LocalMux I__7945 (
            .O(N__36638),
            .I(\c0.data_out_10_7 ));
    Odrv4 I__7944 (
            .O(N__36635),
            .I(\c0.data_out_10_7 ));
    InMux I__7943 (
            .O(N__36630),
            .I(N__36627));
    LocalMux I__7942 (
            .O(N__36627),
            .I(N__36620));
    InMux I__7941 (
            .O(N__36626),
            .I(N__36615));
    InMux I__7940 (
            .O(N__36625),
            .I(N__36615));
    InMux I__7939 (
            .O(N__36624),
            .I(N__36610));
    InMux I__7938 (
            .O(N__36623),
            .I(N__36610));
    Odrv4 I__7937 (
            .O(N__36620),
            .I(data_out_8_3));
    LocalMux I__7936 (
            .O(N__36615),
            .I(data_out_8_3));
    LocalMux I__7935 (
            .O(N__36610),
            .I(data_out_8_3));
    CascadeMux I__7934 (
            .O(N__36603),
            .I(N__36600));
    InMux I__7933 (
            .O(N__36600),
            .I(N__36597));
    LocalMux I__7932 (
            .O(N__36597),
            .I(N__36594));
    Odrv4 I__7931 (
            .O(N__36594),
            .I(\c0.n8_adj_2219 ));
    InMux I__7930 (
            .O(N__36591),
            .I(N__36588));
    LocalMux I__7929 (
            .O(N__36588),
            .I(N__36585));
    Span4Mux_h I__7928 (
            .O(N__36585),
            .I(N__36581));
    InMux I__7927 (
            .O(N__36584),
            .I(N__36578));
    Span4Mux_h I__7926 (
            .O(N__36581),
            .I(N__36575));
    LocalMux I__7925 (
            .O(N__36578),
            .I(data_out_0_3));
    Odrv4 I__7924 (
            .O(N__36575),
            .I(data_out_0_3));
    InMux I__7923 (
            .O(N__36570),
            .I(N__36567));
    LocalMux I__7922 (
            .O(N__36567),
            .I(N__36564));
    Span4Mux_h I__7921 (
            .O(N__36564),
            .I(N__36561));
    Odrv4 I__7920 (
            .O(N__36561),
            .I(\c0.n18376 ));
    CascadeMux I__7919 (
            .O(N__36558),
            .I(N__36554));
    InMux I__7918 (
            .O(N__36557),
            .I(N__36550));
    InMux I__7917 (
            .O(N__36554),
            .I(N__36547));
    InMux I__7916 (
            .O(N__36553),
            .I(N__36544));
    LocalMux I__7915 (
            .O(N__36550),
            .I(N__36541));
    LocalMux I__7914 (
            .O(N__36547),
            .I(N__36536));
    LocalMux I__7913 (
            .O(N__36544),
            .I(N__36533));
    Span4Mux_h I__7912 (
            .O(N__36541),
            .I(N__36530));
    InMux I__7911 (
            .O(N__36540),
            .I(N__36525));
    InMux I__7910 (
            .O(N__36539),
            .I(N__36525));
    Odrv4 I__7909 (
            .O(N__36536),
            .I(data_out_8_2));
    Odrv4 I__7908 (
            .O(N__36533),
            .I(data_out_8_2));
    Odrv4 I__7907 (
            .O(N__36530),
            .I(data_out_8_2));
    LocalMux I__7906 (
            .O(N__36525),
            .I(data_out_8_2));
    CEMux I__7905 (
            .O(N__36516),
            .I(N__36513));
    LocalMux I__7904 (
            .O(N__36513),
            .I(N__36509));
    CEMux I__7903 (
            .O(N__36512),
            .I(N__36506));
    Span4Mux_v I__7902 (
            .O(N__36509),
            .I(N__36503));
    LocalMux I__7901 (
            .O(N__36506),
            .I(N__36500));
    Span4Mux_h I__7900 (
            .O(N__36503),
            .I(N__36495));
    Span4Mux_v I__7899 (
            .O(N__36500),
            .I(N__36495));
    Odrv4 I__7898 (
            .O(N__36495),
            .I(\c0.n11056 ));
    CascadeMux I__7897 (
            .O(N__36492),
            .I(\c0.n18199_cascade_ ));
    InMux I__7896 (
            .O(N__36489),
            .I(N__36486));
    LocalMux I__7895 (
            .O(N__36486),
            .I(N__36482));
    InMux I__7894 (
            .O(N__36485),
            .I(N__36479));
    Span4Mux_v I__7893 (
            .O(N__36482),
            .I(N__36476));
    LocalMux I__7892 (
            .O(N__36479),
            .I(N__36473));
    Span4Mux_h I__7891 (
            .O(N__36476),
            .I(N__36468));
    Span4Mux_v I__7890 (
            .O(N__36473),
            .I(N__36468));
    Odrv4 I__7889 (
            .O(N__36468),
            .I(\c0.n17832 ));
    CascadeMux I__7888 (
            .O(N__36465),
            .I(\c0.n18242_cascade_ ));
    InMux I__7887 (
            .O(N__36462),
            .I(N__36459));
    LocalMux I__7886 (
            .O(N__36459),
            .I(N__36455));
    InMux I__7885 (
            .O(N__36458),
            .I(N__36452));
    Span4Mux_v I__7884 (
            .O(N__36455),
            .I(N__36449));
    LocalMux I__7883 (
            .O(N__36452),
            .I(\c0.data_out_6_6 ));
    Odrv4 I__7882 (
            .O(N__36449),
            .I(\c0.data_out_6_6 ));
    CascadeMux I__7881 (
            .O(N__36444),
            .I(N__36441));
    InMux I__7880 (
            .O(N__36441),
            .I(N__36438));
    LocalMux I__7879 (
            .O(N__36438),
            .I(\c0.n5 ));
    InMux I__7878 (
            .O(N__36435),
            .I(N__36432));
    LocalMux I__7877 (
            .O(N__36432),
            .I(\c0.n18247 ));
    InMux I__7876 (
            .O(N__36429),
            .I(N__36423));
    InMux I__7875 (
            .O(N__36428),
            .I(N__36420));
    InMux I__7874 (
            .O(N__36427),
            .I(N__36417));
    InMux I__7873 (
            .O(N__36426),
            .I(N__36414));
    LocalMux I__7872 (
            .O(N__36423),
            .I(N__36407));
    LocalMux I__7871 (
            .O(N__36420),
            .I(N__36407));
    LocalMux I__7870 (
            .O(N__36417),
            .I(N__36407));
    LocalMux I__7869 (
            .O(N__36414),
            .I(data_out_frame2_15_3));
    Odrv12 I__7868 (
            .O(N__36407),
            .I(data_out_frame2_15_3));
    CascadeMux I__7867 (
            .O(N__36402),
            .I(\c0.n6_adj_2422_cascade_ ));
    InMux I__7866 (
            .O(N__36399),
            .I(N__36393));
    InMux I__7865 (
            .O(N__36398),
            .I(N__36393));
    LocalMux I__7864 (
            .O(N__36393),
            .I(data_out_frame2_18_4));
    CascadeMux I__7863 (
            .O(N__36390),
            .I(\c0.n10870_cascade_ ));
    InMux I__7862 (
            .O(N__36387),
            .I(N__36384));
    LocalMux I__7861 (
            .O(N__36384),
            .I(N__36381));
    Span4Mux_v I__7860 (
            .O(N__36381),
            .I(N__36378));
    Odrv4 I__7859 (
            .O(N__36378),
            .I(\c0.n27_adj_2428 ));
    CascadeMux I__7858 (
            .O(N__36375),
            .I(N__36372));
    InMux I__7857 (
            .O(N__36372),
            .I(N__36369));
    LocalMux I__7856 (
            .O(N__36369),
            .I(\c0.n5_adj_2274 ));
    CascadeMux I__7855 (
            .O(N__36366),
            .I(\c0.n18879_cascade_ ));
    CascadeMux I__7854 (
            .O(N__36363),
            .I(N__36360));
    InMux I__7853 (
            .O(N__36360),
            .I(N__36357));
    LocalMux I__7852 (
            .O(N__36357),
            .I(N__36354));
    Span4Mux_h I__7851 (
            .O(N__36354),
            .I(N__36351));
    Odrv4 I__7850 (
            .O(N__36351),
            .I(\c0.n10852 ));
    CascadeMux I__7849 (
            .O(N__36348),
            .I(N__36345));
    InMux I__7848 (
            .O(N__36345),
            .I(N__36342));
    LocalMux I__7847 (
            .O(N__36342),
            .I(N__36339));
    Span4Mux_v I__7846 (
            .O(N__36339),
            .I(N__36336));
    Span4Mux_h I__7845 (
            .O(N__36336),
            .I(N__36332));
    InMux I__7844 (
            .O(N__36335),
            .I(N__36329));
    IoSpan4Mux I__7843 (
            .O(N__36332),
            .I(N__36326));
    LocalMux I__7842 (
            .O(N__36329),
            .I(N__36323));
    Span4Mux_s1_v I__7841 (
            .O(N__36326),
            .I(N__36320));
    Odrv4 I__7840 (
            .O(N__36323),
            .I(\c0.n10867 ));
    Odrv4 I__7839 (
            .O(N__36320),
            .I(\c0.n10867 ));
    InMux I__7838 (
            .O(N__36315),
            .I(N__36310));
    InMux I__7837 (
            .O(N__36314),
            .I(N__36307));
    InMux I__7836 (
            .O(N__36313),
            .I(N__36303));
    LocalMux I__7835 (
            .O(N__36310),
            .I(N__36300));
    LocalMux I__7834 (
            .O(N__36307),
            .I(N__36297));
    InMux I__7833 (
            .O(N__36306),
            .I(N__36294));
    LocalMux I__7832 (
            .O(N__36303),
            .I(data_out_frame2_8_5));
    Odrv4 I__7831 (
            .O(N__36300),
            .I(data_out_frame2_8_5));
    Odrv4 I__7830 (
            .O(N__36297),
            .I(data_out_frame2_8_5));
    LocalMux I__7829 (
            .O(N__36294),
            .I(data_out_frame2_8_5));
    InMux I__7828 (
            .O(N__36285),
            .I(N__36282));
    LocalMux I__7827 (
            .O(N__36282),
            .I(\c0.n14_adj_2447 ));
    CascadeMux I__7826 (
            .O(N__36279),
            .I(N__36276));
    InMux I__7825 (
            .O(N__36276),
            .I(N__36273));
    LocalMux I__7824 (
            .O(N__36273),
            .I(N__36270));
    Span12Mux_v I__7823 (
            .O(N__36270),
            .I(N__36267));
    Odrv12 I__7822 (
            .O(N__36267),
            .I(\c0.data_out_frame2_19_4 ));
    CascadeMux I__7821 (
            .O(N__36264),
            .I(N__36261));
    InMux I__7820 (
            .O(N__36261),
            .I(N__36258));
    LocalMux I__7819 (
            .O(N__36258),
            .I(\c0.n10_adj_2440 ));
    InMux I__7818 (
            .O(N__36255),
            .I(N__36252));
    LocalMux I__7817 (
            .O(N__36252),
            .I(N__36249));
    Span4Mux_s2_v I__7816 (
            .O(N__36249),
            .I(N__36246));
    Odrv4 I__7815 (
            .O(N__36246),
            .I(\c0.n6_adj_2357 ));
    InMux I__7814 (
            .O(N__36243),
            .I(N__36240));
    LocalMux I__7813 (
            .O(N__36240),
            .I(N__36236));
    InMux I__7812 (
            .O(N__36239),
            .I(N__36233));
    Odrv12 I__7811 (
            .O(N__36236),
            .I(\c0.n10864 ));
    LocalMux I__7810 (
            .O(N__36233),
            .I(\c0.n10864 ));
    InMux I__7809 (
            .O(N__36228),
            .I(N__36224));
    InMux I__7808 (
            .O(N__36227),
            .I(N__36221));
    LocalMux I__7807 (
            .O(N__36224),
            .I(N__36217));
    LocalMux I__7806 (
            .O(N__36221),
            .I(N__36213));
    InMux I__7805 (
            .O(N__36220),
            .I(N__36210));
    Span4Mux_h I__7804 (
            .O(N__36217),
            .I(N__36207));
    InMux I__7803 (
            .O(N__36216),
            .I(N__36204));
    Span4Mux_h I__7802 (
            .O(N__36213),
            .I(N__36201));
    LocalMux I__7801 (
            .O(N__36210),
            .I(data_out_frame2_6_4));
    Odrv4 I__7800 (
            .O(N__36207),
            .I(data_out_frame2_6_4));
    LocalMux I__7799 (
            .O(N__36204),
            .I(data_out_frame2_6_4));
    Odrv4 I__7798 (
            .O(N__36201),
            .I(data_out_frame2_6_4));
    CascadeMux I__7797 (
            .O(N__36192),
            .I(\c0.n10720_cascade_ ));
    InMux I__7796 (
            .O(N__36189),
            .I(N__36186));
    LocalMux I__7795 (
            .O(N__36186),
            .I(N__36180));
    InMux I__7794 (
            .O(N__36185),
            .I(N__36177));
    InMux I__7793 (
            .O(N__36184),
            .I(N__36174));
    InMux I__7792 (
            .O(N__36183),
            .I(N__36171));
    Span4Mux_h I__7791 (
            .O(N__36180),
            .I(N__36168));
    LocalMux I__7790 (
            .O(N__36177),
            .I(N__36165));
    LocalMux I__7789 (
            .O(N__36174),
            .I(N__36162));
    LocalMux I__7788 (
            .O(N__36171),
            .I(data_out_frame2_10_2));
    Odrv4 I__7787 (
            .O(N__36168),
            .I(data_out_frame2_10_2));
    Odrv4 I__7786 (
            .O(N__36165),
            .I(data_out_frame2_10_2));
    Odrv4 I__7785 (
            .O(N__36162),
            .I(data_out_frame2_10_2));
    InMux I__7784 (
            .O(N__36153),
            .I(N__36150));
    LocalMux I__7783 (
            .O(N__36150),
            .I(N__36146));
    InMux I__7782 (
            .O(N__36149),
            .I(N__36143));
    Odrv4 I__7781 (
            .O(N__36146),
            .I(\c0.n10819 ));
    LocalMux I__7780 (
            .O(N__36143),
            .I(\c0.n10819 ));
    InMux I__7779 (
            .O(N__36138),
            .I(N__36135));
    LocalMux I__7778 (
            .O(N__36135),
            .I(N__36131));
    InMux I__7777 (
            .O(N__36134),
            .I(N__36128));
    Span12Mux_s1_v I__7776 (
            .O(N__36131),
            .I(N__36125));
    LocalMux I__7775 (
            .O(N__36128),
            .I(N__36122));
    Odrv12 I__7774 (
            .O(N__36125),
            .I(\c0.n17886 ));
    Odrv4 I__7773 (
            .O(N__36122),
            .I(\c0.n17886 ));
    InMux I__7772 (
            .O(N__36117),
            .I(N__36114));
    LocalMux I__7771 (
            .O(N__36114),
            .I(N__36111));
    Odrv12 I__7770 (
            .O(N__36111),
            .I(\c0.n20_adj_2442 ));
    CascadeMux I__7769 (
            .O(N__36108),
            .I(\c0.n16_cascade_ ));
    InMux I__7768 (
            .O(N__36105),
            .I(N__36101));
    InMux I__7767 (
            .O(N__36104),
            .I(N__36098));
    LocalMux I__7766 (
            .O(N__36101),
            .I(N__36093));
    LocalMux I__7765 (
            .O(N__36098),
            .I(N__36093));
    Span4Mux_s3_v I__7764 (
            .O(N__36093),
            .I(N__36090));
    Odrv4 I__7763 (
            .O(N__36090),
            .I(\c0.n17795 ));
    CascadeMux I__7762 (
            .O(N__36087),
            .I(N__36084));
    InMux I__7761 (
            .O(N__36084),
            .I(N__36081));
    LocalMux I__7760 (
            .O(N__36081),
            .I(N__36078));
    Span4Mux_h I__7759 (
            .O(N__36078),
            .I(N__36075));
    Odrv4 I__7758 (
            .O(N__36075),
            .I(\c0.data_out_frame2_19_5 ));
    InMux I__7757 (
            .O(N__36072),
            .I(N__36063));
    InMux I__7756 (
            .O(N__36071),
            .I(N__36063));
    InMux I__7755 (
            .O(N__36070),
            .I(N__36063));
    LocalMux I__7754 (
            .O(N__36063),
            .I(\c0.n10839 ));
    InMux I__7753 (
            .O(N__36060),
            .I(N__36057));
    LocalMux I__7752 (
            .O(N__36057),
            .I(N__36054));
    Odrv4 I__7751 (
            .O(N__36054),
            .I(\c0.n10890 ));
    InMux I__7750 (
            .O(N__36051),
            .I(N__36046));
    InMux I__7749 (
            .O(N__36050),
            .I(N__36043));
    InMux I__7748 (
            .O(N__36049),
            .I(N__36040));
    LocalMux I__7747 (
            .O(N__36046),
            .I(N__36036));
    LocalMux I__7746 (
            .O(N__36043),
            .I(N__36033));
    LocalMux I__7745 (
            .O(N__36040),
            .I(N__36030));
    InMux I__7744 (
            .O(N__36039),
            .I(N__36027));
    Span4Mux_v I__7743 (
            .O(N__36036),
            .I(N__36024));
    Span4Mux_s3_v I__7742 (
            .O(N__36033),
            .I(N__36019));
    Span4Mux_h I__7741 (
            .O(N__36030),
            .I(N__36019));
    LocalMux I__7740 (
            .O(N__36027),
            .I(data_out_frame2_10_5));
    Odrv4 I__7739 (
            .O(N__36024),
            .I(data_out_frame2_10_5));
    Odrv4 I__7738 (
            .O(N__36019),
            .I(data_out_frame2_10_5));
    CascadeMux I__7737 (
            .O(N__36012),
            .I(N__36008));
    InMux I__7736 (
            .O(N__36011),
            .I(N__36005));
    InMux I__7735 (
            .O(N__36008),
            .I(N__36002));
    LocalMux I__7734 (
            .O(N__36005),
            .I(N__35999));
    LocalMux I__7733 (
            .O(N__36002),
            .I(N__35996));
    Span4Mux_v I__7732 (
            .O(N__35999),
            .I(N__35993));
    Odrv4 I__7731 (
            .O(N__35996),
            .I(\c0.n10816 ));
    Odrv4 I__7730 (
            .O(N__35993),
            .I(\c0.n10816 ));
    CascadeMux I__7729 (
            .O(N__35988),
            .I(\c0.n12_adj_2446_cascade_ ));
    InMux I__7728 (
            .O(N__35985),
            .I(N__35981));
    InMux I__7727 (
            .O(N__35984),
            .I(N__35976));
    LocalMux I__7726 (
            .O(N__35981),
            .I(N__35973));
    InMux I__7725 (
            .O(N__35980),
            .I(N__35968));
    InMux I__7724 (
            .O(N__35979),
            .I(N__35968));
    LocalMux I__7723 (
            .O(N__35976),
            .I(data_out_frame2_15_1));
    Odrv4 I__7722 (
            .O(N__35973),
            .I(data_out_frame2_15_1));
    LocalMux I__7721 (
            .O(N__35968),
            .I(data_out_frame2_15_1));
    InMux I__7720 (
            .O(N__35961),
            .I(N__35958));
    LocalMux I__7719 (
            .O(N__35958),
            .I(N__35955));
    Span4Mux_s0_v I__7718 (
            .O(N__35955),
            .I(N__35952));
    Odrv4 I__7717 (
            .O(N__35952),
            .I(\c0.n10829 ));
    CascadeMux I__7716 (
            .O(N__35949),
            .I(\c0.n10890_cascade_ ));
    InMux I__7715 (
            .O(N__35946),
            .I(N__35943));
    LocalMux I__7714 (
            .O(N__35943),
            .I(N__35940));
    Span4Mux_h I__7713 (
            .O(N__35940),
            .I(N__35937));
    Odrv4 I__7712 (
            .O(N__35937),
            .I(\c0.n17_adj_2449 ));
    CascadeMux I__7711 (
            .O(N__35934),
            .I(\c0.n16_adj_2448_cascade_ ));
    InMux I__7710 (
            .O(N__35931),
            .I(N__35927));
    InMux I__7709 (
            .O(N__35930),
            .I(N__35924));
    LocalMux I__7708 (
            .O(N__35927),
            .I(N__35919));
    LocalMux I__7707 (
            .O(N__35924),
            .I(N__35919));
    Span4Mux_s1_v I__7706 (
            .O(N__35919),
            .I(N__35916));
    Odrv4 I__7705 (
            .O(N__35916),
            .I(\c0.n17911 ));
    InMux I__7704 (
            .O(N__35913),
            .I(N__35910));
    LocalMux I__7703 (
            .O(N__35910),
            .I(\c0.n15_adj_2445 ));
    CascadeMux I__7702 (
            .O(N__35907),
            .I(\c0.n14_adj_2444_cascade_ ));
    InMux I__7701 (
            .O(N__35904),
            .I(N__35901));
    LocalMux I__7700 (
            .O(N__35901),
            .I(N__35894));
    InMux I__7699 (
            .O(N__35900),
            .I(N__35889));
    InMux I__7698 (
            .O(N__35899),
            .I(N__35889));
    InMux I__7697 (
            .O(N__35898),
            .I(N__35884));
    InMux I__7696 (
            .O(N__35897),
            .I(N__35884));
    Odrv4 I__7695 (
            .O(N__35894),
            .I(data_out_frame2_16_1));
    LocalMux I__7694 (
            .O(N__35889),
            .I(data_out_frame2_16_1));
    LocalMux I__7693 (
            .O(N__35884),
            .I(data_out_frame2_16_1));
    InMux I__7692 (
            .O(N__35877),
            .I(N__35874));
    LocalMux I__7691 (
            .O(N__35874),
            .I(N__35871));
    Odrv12 I__7690 (
            .O(N__35871),
            .I(\c0.data_out_frame2_20_5 ));
    CascadeMux I__7689 (
            .O(N__35868),
            .I(N__35865));
    InMux I__7688 (
            .O(N__35865),
            .I(N__35862));
    LocalMux I__7687 (
            .O(N__35862),
            .I(\c0.n16_adj_2358 ));
    InMux I__7686 (
            .O(N__35859),
            .I(N__35854));
    InMux I__7685 (
            .O(N__35858),
            .I(N__35847));
    InMux I__7684 (
            .O(N__35857),
            .I(N__35847));
    LocalMux I__7683 (
            .O(N__35854),
            .I(N__35844));
    InMux I__7682 (
            .O(N__35853),
            .I(N__35841));
    InMux I__7681 (
            .O(N__35852),
            .I(N__35838));
    LocalMux I__7680 (
            .O(N__35847),
            .I(N__35835));
    Span4Mux_v I__7679 (
            .O(N__35844),
            .I(N__35830));
    LocalMux I__7678 (
            .O(N__35841),
            .I(N__35830));
    LocalMux I__7677 (
            .O(N__35838),
            .I(\c0.data_out_7_4 ));
    Odrv12 I__7676 (
            .O(N__35835),
            .I(\c0.data_out_7_4 ));
    Odrv4 I__7675 (
            .O(N__35830),
            .I(\c0.data_out_7_4 ));
    InMux I__7674 (
            .O(N__35823),
            .I(N__35817));
    InMux I__7673 (
            .O(N__35822),
            .I(N__35817));
    LocalMux I__7672 (
            .O(N__35817),
            .I(data_out_3_2));
    CascadeMux I__7671 (
            .O(N__35814),
            .I(N__35811));
    InMux I__7670 (
            .O(N__35811),
            .I(N__35805));
    InMux I__7669 (
            .O(N__35810),
            .I(N__35805));
    LocalMux I__7668 (
            .O(N__35805),
            .I(\c0.data_out_1_2 ));
    InMux I__7667 (
            .O(N__35802),
            .I(N__35799));
    LocalMux I__7666 (
            .O(N__35799),
            .I(N__35796));
    Odrv12 I__7665 (
            .O(N__35796),
            .I(\c0.n18223 ));
    InMux I__7664 (
            .O(N__35793),
            .I(N__35789));
    InMux I__7663 (
            .O(N__35792),
            .I(N__35786));
    LocalMux I__7662 (
            .O(N__35789),
            .I(N__35783));
    LocalMux I__7661 (
            .O(N__35786),
            .I(data_out_2_2));
    Odrv4 I__7660 (
            .O(N__35783),
            .I(data_out_2_2));
    IoInMux I__7659 (
            .O(N__35778),
            .I(N__35775));
    LocalMux I__7658 (
            .O(N__35775),
            .I(N__35772));
    Span4Mux_s3_v I__7657 (
            .O(N__35772),
            .I(N__35769));
    Sp12to4 I__7656 (
            .O(N__35769),
            .I(N__35766));
    Span12Mux_h I__7655 (
            .O(N__35766),
            .I(N__35763));
    Odrv12 I__7654 (
            .O(N__35763),
            .I(PIN_24_c_3));
    CEMux I__7653 (
            .O(N__35760),
            .I(N__35757));
    LocalMux I__7652 (
            .O(N__35757),
            .I(N__35754));
    Span4Mux_v I__7651 (
            .O(N__35754),
            .I(N__35751));
    Odrv4 I__7650 (
            .O(N__35751),
            .I(\control.n6 ));
    SRMux I__7649 (
            .O(N__35748),
            .I(N__35745));
    LocalMux I__7648 (
            .O(N__35745),
            .I(\control.n17251 ));
    IoInMux I__7647 (
            .O(N__35742),
            .I(N__35739));
    LocalMux I__7646 (
            .O(N__35739),
            .I(N__35736));
    Span12Mux_s10_v I__7645 (
            .O(N__35736),
            .I(N__35733));
    Span12Mux_h I__7644 (
            .O(N__35733),
            .I(N__35730));
    Odrv12 I__7643 (
            .O(N__35730),
            .I(PIN_23_c_4));
    CEMux I__7642 (
            .O(N__35727),
            .I(N__35724));
    LocalMux I__7641 (
            .O(N__35724),
            .I(N__35720));
    CEMux I__7640 (
            .O(N__35723),
            .I(N__35717));
    Span4Mux_v I__7639 (
            .O(N__35720),
            .I(N__35714));
    LocalMux I__7638 (
            .O(N__35717),
            .I(N__35711));
    Span4Mux_h I__7637 (
            .O(N__35714),
            .I(N__35708));
    Span4Mux_v I__7636 (
            .O(N__35711),
            .I(N__35705));
    Odrv4 I__7635 (
            .O(N__35708),
            .I(\control.n6_adj_2460 ));
    Odrv4 I__7634 (
            .O(N__35705),
            .I(\control.n6_adj_2460 ));
    SRMux I__7633 (
            .O(N__35700),
            .I(N__35697));
    LocalMux I__7632 (
            .O(N__35697),
            .I(N__35694));
    Odrv12 I__7631 (
            .O(N__35694),
            .I(\control.n10490 ));
    InMux I__7630 (
            .O(N__35691),
            .I(N__35686));
    InMux I__7629 (
            .O(N__35690),
            .I(N__35683));
    InMux I__7628 (
            .O(N__35689),
            .I(N__35680));
    LocalMux I__7627 (
            .O(N__35686),
            .I(N__35676));
    LocalMux I__7626 (
            .O(N__35683),
            .I(N__35672));
    LocalMux I__7625 (
            .O(N__35680),
            .I(N__35669));
    InMux I__7624 (
            .O(N__35679),
            .I(N__35666));
    Span4Mux_h I__7623 (
            .O(N__35676),
            .I(N__35660));
    InMux I__7622 (
            .O(N__35675),
            .I(N__35657));
    Span4Mux_v I__7621 (
            .O(N__35672),
            .I(N__35649));
    Span4Mux_h I__7620 (
            .O(N__35669),
            .I(N__35649));
    LocalMux I__7619 (
            .O(N__35666),
            .I(N__35649));
    InMux I__7618 (
            .O(N__35665),
            .I(N__35646));
    InMux I__7617 (
            .O(N__35664),
            .I(N__35643));
    InMux I__7616 (
            .O(N__35663),
            .I(N__35640));
    Span4Mux_h I__7615 (
            .O(N__35660),
            .I(N__35633));
    LocalMux I__7614 (
            .O(N__35657),
            .I(N__35633));
    InMux I__7613 (
            .O(N__35656),
            .I(N__35630));
    Span4Mux_v I__7612 (
            .O(N__35649),
            .I(N__35625));
    LocalMux I__7611 (
            .O(N__35646),
            .I(N__35625));
    LocalMux I__7610 (
            .O(N__35643),
            .I(N__35620));
    LocalMux I__7609 (
            .O(N__35640),
            .I(N__35620));
    InMux I__7608 (
            .O(N__35639),
            .I(N__35617));
    InMux I__7607 (
            .O(N__35638),
            .I(N__35614));
    Span4Mux_h I__7606 (
            .O(N__35633),
            .I(N__35611));
    LocalMux I__7605 (
            .O(N__35630),
            .I(N__35608));
    Span4Mux_h I__7604 (
            .O(N__35625),
            .I(N__35603));
    Span4Mux_v I__7603 (
            .O(N__35620),
            .I(N__35603));
    LocalMux I__7602 (
            .O(N__35617),
            .I(N__35600));
    LocalMux I__7601 (
            .O(N__35614),
            .I(N__35593));
    Sp12to4 I__7600 (
            .O(N__35611),
            .I(N__35593));
    Sp12to4 I__7599 (
            .O(N__35608),
            .I(N__35593));
    Span4Mux_h I__7598 (
            .O(N__35603),
            .I(N__35588));
    Span4Mux_v I__7597 (
            .O(N__35600),
            .I(N__35588));
    Span12Mux_s9_v I__7596 (
            .O(N__35593),
            .I(N__35585));
    Span4Mux_v I__7595 (
            .O(N__35588),
            .I(N__35582));
    Odrv12 I__7594 (
            .O(N__35585),
            .I(hall3));
    Odrv4 I__7593 (
            .O(N__35582),
            .I(hall3));
    InMux I__7592 (
            .O(N__35577),
            .I(N__35571));
    InMux I__7591 (
            .O(N__35576),
            .I(N__35568));
    InMux I__7590 (
            .O(N__35575),
            .I(N__35563));
    InMux I__7589 (
            .O(N__35574),
            .I(N__35560));
    LocalMux I__7588 (
            .O(N__35571),
            .I(N__35556));
    LocalMux I__7587 (
            .O(N__35568),
            .I(N__35553));
    InMux I__7586 (
            .O(N__35567),
            .I(N__35550));
    InMux I__7585 (
            .O(N__35566),
            .I(N__35547));
    LocalMux I__7584 (
            .O(N__35563),
            .I(N__35542));
    LocalMux I__7583 (
            .O(N__35560),
            .I(N__35539));
    InMux I__7582 (
            .O(N__35559),
            .I(N__35536));
    Span4Mux_v I__7581 (
            .O(N__35556),
            .I(N__35527));
    Span4Mux_v I__7580 (
            .O(N__35553),
            .I(N__35527));
    LocalMux I__7579 (
            .O(N__35550),
            .I(N__35527));
    LocalMux I__7578 (
            .O(N__35547),
            .I(N__35527));
    InMux I__7577 (
            .O(N__35546),
            .I(N__35524));
    InMux I__7576 (
            .O(N__35545),
            .I(N__35521));
    Span4Mux_v I__7575 (
            .O(N__35542),
            .I(N__35516));
    Span4Mux_v I__7574 (
            .O(N__35539),
            .I(N__35516));
    LocalMux I__7573 (
            .O(N__35536),
            .I(N__35513));
    Span4Mux_h I__7572 (
            .O(N__35527),
            .I(N__35508));
    LocalMux I__7571 (
            .O(N__35524),
            .I(N__35505));
    LocalMux I__7570 (
            .O(N__35521),
            .I(N__35502));
    Span4Mux_h I__7569 (
            .O(N__35516),
            .I(N__35497));
    Span4Mux_v I__7568 (
            .O(N__35513),
            .I(N__35497));
    InMux I__7567 (
            .O(N__35512),
            .I(N__35494));
    InMux I__7566 (
            .O(N__35511),
            .I(N__35491));
    Span4Mux_h I__7565 (
            .O(N__35508),
            .I(N__35486));
    Span4Mux_v I__7564 (
            .O(N__35505),
            .I(N__35486));
    Span12Mux_h I__7563 (
            .O(N__35502),
            .I(N__35477));
    Sp12to4 I__7562 (
            .O(N__35497),
            .I(N__35477));
    LocalMux I__7561 (
            .O(N__35494),
            .I(N__35477));
    LocalMux I__7560 (
            .O(N__35491),
            .I(N__35477));
    Odrv4 I__7559 (
            .O(N__35486),
            .I(hall2));
    Odrv12 I__7558 (
            .O(N__35477),
            .I(hall2));
    CascadeMux I__7557 (
            .O(N__35472),
            .I(N__35467));
    CascadeMux I__7556 (
            .O(N__35471),
            .I(N__35464));
    InMux I__7555 (
            .O(N__35470),
            .I(N__35458));
    InMux I__7554 (
            .O(N__35467),
            .I(N__35455));
    InMux I__7553 (
            .O(N__35464),
            .I(N__35451));
    InMux I__7552 (
            .O(N__35463),
            .I(N__35448));
    InMux I__7551 (
            .O(N__35462),
            .I(N__35445));
    InMux I__7550 (
            .O(N__35461),
            .I(N__35438));
    LocalMux I__7549 (
            .O(N__35458),
            .I(N__35433));
    LocalMux I__7548 (
            .O(N__35455),
            .I(N__35433));
    CascadeMux I__7547 (
            .O(N__35454),
            .I(N__35430));
    LocalMux I__7546 (
            .O(N__35451),
            .I(N__35423));
    LocalMux I__7545 (
            .O(N__35448),
            .I(N__35423));
    LocalMux I__7544 (
            .O(N__35445),
            .I(N__35423));
    InMux I__7543 (
            .O(N__35444),
            .I(N__35420));
    InMux I__7542 (
            .O(N__35443),
            .I(N__35415));
    InMux I__7541 (
            .O(N__35442),
            .I(N__35415));
    InMux I__7540 (
            .O(N__35441),
            .I(N__35412));
    LocalMux I__7539 (
            .O(N__35438),
            .I(N__35408));
    Span4Mux_v I__7538 (
            .O(N__35433),
            .I(N__35405));
    InMux I__7537 (
            .O(N__35430),
            .I(N__35402));
    Span4Mux_v I__7536 (
            .O(N__35423),
            .I(N__35399));
    LocalMux I__7535 (
            .O(N__35420),
            .I(N__35392));
    LocalMux I__7534 (
            .O(N__35415),
            .I(N__35392));
    LocalMux I__7533 (
            .O(N__35412),
            .I(N__35392));
    InMux I__7532 (
            .O(N__35411),
            .I(N__35389));
    Span4Mux_v I__7531 (
            .O(N__35408),
            .I(N__35386));
    Span4Mux_h I__7530 (
            .O(N__35405),
            .I(N__35383));
    LocalMux I__7529 (
            .O(N__35402),
            .I(N__35380));
    Span4Mux_h I__7528 (
            .O(N__35399),
            .I(N__35375));
    Span4Mux_v I__7527 (
            .O(N__35392),
            .I(N__35375));
    LocalMux I__7526 (
            .O(N__35389),
            .I(N__35372));
    Sp12to4 I__7525 (
            .O(N__35386),
            .I(N__35369));
    Span4Mux_h I__7524 (
            .O(N__35383),
            .I(N__35364));
    Span4Mux_v I__7523 (
            .O(N__35380),
            .I(N__35364));
    Span4Mux_h I__7522 (
            .O(N__35375),
            .I(N__35359));
    Span4Mux_v I__7521 (
            .O(N__35372),
            .I(N__35359));
    Odrv12 I__7520 (
            .O(N__35369),
            .I(hall1));
    Odrv4 I__7519 (
            .O(N__35364),
            .I(hall1));
    Odrv4 I__7518 (
            .O(N__35359),
            .I(hall1));
    SRMux I__7517 (
            .O(N__35352),
            .I(N__35348));
    InMux I__7516 (
            .O(N__35351),
            .I(N__35344));
    LocalMux I__7515 (
            .O(N__35348),
            .I(N__35341));
    SRMux I__7514 (
            .O(N__35347),
            .I(N__35338));
    LocalMux I__7513 (
            .O(N__35344),
            .I(N__35334));
    Span4Mux_v I__7512 (
            .O(N__35341),
            .I(N__35329));
    LocalMux I__7511 (
            .O(N__35338),
            .I(N__35329));
    InMux I__7510 (
            .O(N__35337),
            .I(N__35326));
    Span4Mux_v I__7509 (
            .O(N__35334),
            .I(N__35321));
    Span4Mux_h I__7508 (
            .O(N__35329),
            .I(N__35316));
    LocalMux I__7507 (
            .O(N__35326),
            .I(N__35316));
    InMux I__7506 (
            .O(N__35325),
            .I(N__35312));
    InMux I__7505 (
            .O(N__35324),
            .I(N__35309));
    Span4Mux_h I__7504 (
            .O(N__35321),
            .I(N__35304));
    Span4Mux_v I__7503 (
            .O(N__35316),
            .I(N__35304));
    InMux I__7502 (
            .O(N__35315),
            .I(N__35301));
    LocalMux I__7501 (
            .O(N__35312),
            .I(\control.PHASES_5__N_2160 ));
    LocalMux I__7500 (
            .O(N__35309),
            .I(\control.PHASES_5__N_2160 ));
    Odrv4 I__7499 (
            .O(N__35304),
            .I(\control.PHASES_5__N_2160 ));
    LocalMux I__7498 (
            .O(N__35301),
            .I(\control.PHASES_5__N_2160 ));
    IoInMux I__7497 (
            .O(N__35292),
            .I(N__35289));
    LocalMux I__7496 (
            .O(N__35289),
            .I(N__35286));
    Span12Mux_s3_v I__7495 (
            .O(N__35286),
            .I(N__35283));
    Span12Mux_h I__7494 (
            .O(N__35283),
            .I(N__35280));
    Odrv12 I__7493 (
            .O(N__35280),
            .I(\control.PHASES_5_N_2130_5 ));
    CascadeMux I__7492 (
            .O(N__35277),
            .I(N__35274));
    InMux I__7491 (
            .O(N__35274),
            .I(N__35271));
    LocalMux I__7490 (
            .O(N__35271),
            .I(N__35268));
    Span12Mux_h I__7489 (
            .O(N__35268),
            .I(N__35265));
    Odrv12 I__7488 (
            .O(N__35265),
            .I(\c0.n17748 ));
    InMux I__7487 (
            .O(N__35262),
            .I(N__35259));
    LocalMux I__7486 (
            .O(N__35259),
            .I(N__35256));
    Odrv4 I__7485 (
            .O(N__35256),
            .I(\c0.n18191 ));
    CascadeMux I__7484 (
            .O(N__35253),
            .I(\c0.n18867_cascade_ ));
    InMux I__7483 (
            .O(N__35250),
            .I(N__35240));
    InMux I__7482 (
            .O(N__35249),
            .I(N__35240));
    CascadeMux I__7481 (
            .O(N__35248),
            .I(N__35237));
    InMux I__7480 (
            .O(N__35247),
            .I(N__35227));
    InMux I__7479 (
            .O(N__35246),
            .I(N__35224));
    InMux I__7478 (
            .O(N__35245),
            .I(N__35221));
    LocalMux I__7477 (
            .O(N__35240),
            .I(N__35213));
    InMux I__7476 (
            .O(N__35237),
            .I(N__35208));
    InMux I__7475 (
            .O(N__35236),
            .I(N__35208));
    InMux I__7474 (
            .O(N__35235),
            .I(N__35203));
    InMux I__7473 (
            .O(N__35234),
            .I(N__35203));
    InMux I__7472 (
            .O(N__35233),
            .I(N__35196));
    InMux I__7471 (
            .O(N__35232),
            .I(N__35196));
    InMux I__7470 (
            .O(N__35231),
            .I(N__35196));
    InMux I__7469 (
            .O(N__35230),
            .I(N__35187));
    LocalMux I__7468 (
            .O(N__35227),
            .I(N__35180));
    LocalMux I__7467 (
            .O(N__35224),
            .I(N__35180));
    LocalMux I__7466 (
            .O(N__35221),
            .I(N__35180));
    InMux I__7465 (
            .O(N__35220),
            .I(N__35177));
    InMux I__7464 (
            .O(N__35219),
            .I(N__35168));
    InMux I__7463 (
            .O(N__35218),
            .I(N__35168));
    InMux I__7462 (
            .O(N__35217),
            .I(N__35168));
    InMux I__7461 (
            .O(N__35216),
            .I(N__35168));
    Span4Mux_h I__7460 (
            .O(N__35213),
            .I(N__35165));
    LocalMux I__7459 (
            .O(N__35208),
            .I(N__35162));
    LocalMux I__7458 (
            .O(N__35203),
            .I(N__35157));
    LocalMux I__7457 (
            .O(N__35196),
            .I(N__35157));
    InMux I__7456 (
            .O(N__35195),
            .I(N__35154));
    InMux I__7455 (
            .O(N__35194),
            .I(N__35145));
    InMux I__7454 (
            .O(N__35193),
            .I(N__35145));
    InMux I__7453 (
            .O(N__35192),
            .I(N__35145));
    InMux I__7452 (
            .O(N__35191),
            .I(N__35145));
    InMux I__7451 (
            .O(N__35190),
            .I(N__35141));
    LocalMux I__7450 (
            .O(N__35187),
            .I(N__35134));
    Span4Mux_v I__7449 (
            .O(N__35180),
            .I(N__35134));
    LocalMux I__7448 (
            .O(N__35177),
            .I(N__35134));
    LocalMux I__7447 (
            .O(N__35168),
            .I(N__35127));
    Span4Mux_v I__7446 (
            .O(N__35165),
            .I(N__35127));
    Span4Mux_h I__7445 (
            .O(N__35162),
            .I(N__35127));
    Span12Mux_h I__7444 (
            .O(N__35157),
            .I(N__35120));
    LocalMux I__7443 (
            .O(N__35154),
            .I(N__35120));
    LocalMux I__7442 (
            .O(N__35145),
            .I(N__35120));
    InMux I__7441 (
            .O(N__35144),
            .I(N__35117));
    LocalMux I__7440 (
            .O(N__35141),
            .I(byte_transmit_counter_2));
    Odrv4 I__7439 (
            .O(N__35134),
            .I(byte_transmit_counter_2));
    Odrv4 I__7438 (
            .O(N__35127),
            .I(byte_transmit_counter_2));
    Odrv12 I__7437 (
            .O(N__35120),
            .I(byte_transmit_counter_2));
    LocalMux I__7436 (
            .O(N__35117),
            .I(byte_transmit_counter_2));
    InMux I__7435 (
            .O(N__35106),
            .I(N__35103));
    LocalMux I__7434 (
            .O(N__35103),
            .I(N__35100));
    Odrv4 I__7433 (
            .O(N__35100),
            .I(n10_adj_2505));
    CascadeMux I__7432 (
            .O(N__35097),
            .I(n18870_cascade_));
    InMux I__7431 (
            .O(N__35094),
            .I(N__35089));
    InMux I__7430 (
            .O(N__35093),
            .I(N__35085));
    InMux I__7429 (
            .O(N__35092),
            .I(N__35082));
    LocalMux I__7428 (
            .O(N__35089),
            .I(N__35077));
    InMux I__7427 (
            .O(N__35088),
            .I(N__35074));
    LocalMux I__7426 (
            .O(N__35085),
            .I(N__35066));
    LocalMux I__7425 (
            .O(N__35082),
            .I(N__35066));
    InMux I__7424 (
            .O(N__35081),
            .I(N__35063));
    InMux I__7423 (
            .O(N__35080),
            .I(N__35060));
    Span4Mux_h I__7422 (
            .O(N__35077),
            .I(N__35055));
    LocalMux I__7421 (
            .O(N__35074),
            .I(N__35055));
    InMux I__7420 (
            .O(N__35073),
            .I(N__35050));
    InMux I__7419 (
            .O(N__35072),
            .I(N__35050));
    InMux I__7418 (
            .O(N__35071),
            .I(N__35046));
    Span4Mux_v I__7417 (
            .O(N__35066),
            .I(N__35041));
    LocalMux I__7416 (
            .O(N__35063),
            .I(N__35041));
    LocalMux I__7415 (
            .O(N__35060),
            .I(N__35038));
    Span4Mux_v I__7414 (
            .O(N__35055),
            .I(N__35033));
    LocalMux I__7413 (
            .O(N__35050),
            .I(N__35033));
    InMux I__7412 (
            .O(N__35049),
            .I(N__35030));
    LocalMux I__7411 (
            .O(N__35046),
            .I(byte_transmit_counter_3));
    Odrv4 I__7410 (
            .O(N__35041),
            .I(byte_transmit_counter_3));
    Odrv12 I__7409 (
            .O(N__35038),
            .I(byte_transmit_counter_3));
    Odrv4 I__7408 (
            .O(N__35033),
            .I(byte_transmit_counter_3));
    LocalMux I__7407 (
            .O(N__35030),
            .I(byte_transmit_counter_3));
    InMux I__7406 (
            .O(N__35019),
            .I(N__35016));
    LocalMux I__7405 (
            .O(N__35016),
            .I(n10_adj_2530));
    CascadeMux I__7404 (
            .O(N__35013),
            .I(N__35010));
    InMux I__7403 (
            .O(N__35010),
            .I(N__35007));
    LocalMux I__7402 (
            .O(N__35007),
            .I(\c0.n5_adj_2214 ));
    InMux I__7401 (
            .O(N__35004),
            .I(N__35000));
    InMux I__7400 (
            .O(N__35003),
            .I(N__34997));
    LocalMux I__7399 (
            .O(N__35000),
            .I(N__34994));
    LocalMux I__7398 (
            .O(N__34997),
            .I(\c0.data_out_1_4 ));
    Odrv4 I__7397 (
            .O(N__34994),
            .I(\c0.data_out_1_4 ));
    InMux I__7396 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__7395 (
            .O(N__34986),
            .I(\c0.n18190 ));
    InMux I__7394 (
            .O(N__34983),
            .I(N__34980));
    LocalMux I__7393 (
            .O(N__34980),
            .I(N__34977));
    Odrv4 I__7392 (
            .O(N__34977),
            .I(\c0.n2_adj_2348 ));
    InMux I__7391 (
            .O(N__34974),
            .I(N__34971));
    LocalMux I__7390 (
            .O(N__34971),
            .I(\c0.n18334 ));
    InMux I__7389 (
            .O(N__34968),
            .I(N__34965));
    LocalMux I__7388 (
            .O(N__34965),
            .I(\c0.n17819 ));
    InMux I__7387 (
            .O(N__34962),
            .I(N__34959));
    LocalMux I__7386 (
            .O(N__34959),
            .I(\c0.n6_adj_2277 ));
    CascadeMux I__7385 (
            .O(N__34956),
            .I(N__34952));
    CascadeMux I__7384 (
            .O(N__34955),
            .I(N__34949));
    InMux I__7383 (
            .O(N__34952),
            .I(N__34945));
    InMux I__7382 (
            .O(N__34949),
            .I(N__34942));
    InMux I__7381 (
            .O(N__34948),
            .I(N__34939));
    LocalMux I__7380 (
            .O(N__34945),
            .I(\c0.data_out_9_4 ));
    LocalMux I__7379 (
            .O(N__34942),
            .I(\c0.data_out_9_4 ));
    LocalMux I__7378 (
            .O(N__34939),
            .I(\c0.data_out_9_4 ));
    CascadeMux I__7377 (
            .O(N__34932),
            .I(\c0.n8_adj_2211_cascade_ ));
    CascadeMux I__7376 (
            .O(N__34929),
            .I(\c0.n18222_cascade_ ));
    CascadeMux I__7375 (
            .O(N__34926),
            .I(\c0.n18693_cascade_ ));
    InMux I__7374 (
            .O(N__34923),
            .I(N__34920));
    LocalMux I__7373 (
            .O(N__34920),
            .I(N__34917));
    Odrv4 I__7372 (
            .O(N__34917),
            .I(n18696));
    InMux I__7371 (
            .O(N__34914),
            .I(N__34905));
    InMux I__7370 (
            .O(N__34913),
            .I(N__34905));
    InMux I__7369 (
            .O(N__34912),
            .I(N__34900));
    InMux I__7368 (
            .O(N__34911),
            .I(N__34900));
    InMux I__7367 (
            .O(N__34910),
            .I(N__34897));
    LocalMux I__7366 (
            .O(N__34905),
            .I(N__34890));
    LocalMux I__7365 (
            .O(N__34900),
            .I(N__34890));
    LocalMux I__7364 (
            .O(N__34897),
            .I(N__34890));
    Span4Mux_v I__7363 (
            .O(N__34890),
            .I(N__34887));
    Odrv4 I__7362 (
            .O(N__34887),
            .I(\c0.data_out_6_2 ));
    InMux I__7361 (
            .O(N__34884),
            .I(N__34881));
    LocalMux I__7360 (
            .O(N__34881),
            .I(\c0.n5_adj_2347 ));
    InMux I__7359 (
            .O(N__34878),
            .I(N__34873));
    InMux I__7358 (
            .O(N__34877),
            .I(N__34862));
    InMux I__7357 (
            .O(N__34876),
            .I(N__34862));
    LocalMux I__7356 (
            .O(N__34873),
            .I(N__34859));
    InMux I__7355 (
            .O(N__34872),
            .I(N__34853));
    InMux I__7354 (
            .O(N__34871),
            .I(N__34848));
    InMux I__7353 (
            .O(N__34870),
            .I(N__34845));
    InMux I__7352 (
            .O(N__34869),
            .I(N__34839));
    InMux I__7351 (
            .O(N__34868),
            .I(N__34839));
    InMux I__7350 (
            .O(N__34867),
            .I(N__34836));
    LocalMux I__7349 (
            .O(N__34862),
            .I(N__34829));
    Span4Mux_v I__7348 (
            .O(N__34859),
            .I(N__34826));
    InMux I__7347 (
            .O(N__34858),
            .I(N__34823));
    InMux I__7346 (
            .O(N__34857),
            .I(N__34820));
    CascadeMux I__7345 (
            .O(N__34856),
            .I(N__34817));
    LocalMux I__7344 (
            .O(N__34853),
            .I(N__34814));
    InMux I__7343 (
            .O(N__34852),
            .I(N__34811));
    InMux I__7342 (
            .O(N__34851),
            .I(N__34808));
    LocalMux I__7341 (
            .O(N__34848),
            .I(N__34805));
    LocalMux I__7340 (
            .O(N__34845),
            .I(N__34802));
    InMux I__7339 (
            .O(N__34844),
            .I(N__34799));
    LocalMux I__7338 (
            .O(N__34839),
            .I(N__34796));
    LocalMux I__7337 (
            .O(N__34836),
            .I(N__34793));
    InMux I__7336 (
            .O(N__34835),
            .I(N__34784));
    InMux I__7335 (
            .O(N__34834),
            .I(N__34784));
    InMux I__7334 (
            .O(N__34833),
            .I(N__34784));
    InMux I__7333 (
            .O(N__34832),
            .I(N__34784));
    Sp12to4 I__7332 (
            .O(N__34829),
            .I(N__34775));
    Sp12to4 I__7331 (
            .O(N__34826),
            .I(N__34775));
    LocalMux I__7330 (
            .O(N__34823),
            .I(N__34775));
    LocalMux I__7329 (
            .O(N__34820),
            .I(N__34775));
    InMux I__7328 (
            .O(N__34817),
            .I(N__34771));
    Span12Mux_v I__7327 (
            .O(N__34814),
            .I(N__34768));
    LocalMux I__7326 (
            .O(N__34811),
            .I(N__34763));
    LocalMux I__7325 (
            .O(N__34808),
            .I(N__34763));
    Span4Mux_v I__7324 (
            .O(N__34805),
            .I(N__34760));
    Span4Mux_v I__7323 (
            .O(N__34802),
            .I(N__34753));
    LocalMux I__7322 (
            .O(N__34799),
            .I(N__34753));
    Span4Mux_h I__7321 (
            .O(N__34796),
            .I(N__34753));
    Span12Mux_v I__7320 (
            .O(N__34793),
            .I(N__34746));
    LocalMux I__7319 (
            .O(N__34784),
            .I(N__34746));
    Span12Mux_h I__7318 (
            .O(N__34775),
            .I(N__34746));
    InMux I__7317 (
            .O(N__34774),
            .I(N__34743));
    LocalMux I__7316 (
            .O(N__34771),
            .I(byte_transmit_counter_1));
    Odrv12 I__7315 (
            .O(N__34768),
            .I(byte_transmit_counter_1));
    Odrv4 I__7314 (
            .O(N__34763),
            .I(byte_transmit_counter_1));
    Odrv4 I__7313 (
            .O(N__34760),
            .I(byte_transmit_counter_1));
    Odrv4 I__7312 (
            .O(N__34753),
            .I(byte_transmit_counter_1));
    Odrv12 I__7311 (
            .O(N__34746),
            .I(byte_transmit_counter_1));
    LocalMux I__7310 (
            .O(N__34743),
            .I(byte_transmit_counter_1));
    InMux I__7309 (
            .O(N__34728),
            .I(N__34725));
    LocalMux I__7308 (
            .O(N__34725),
            .I(N__34720));
    InMux I__7307 (
            .O(N__34724),
            .I(N__34715));
    InMux I__7306 (
            .O(N__34723),
            .I(N__34715));
    Odrv4 I__7305 (
            .O(N__34720),
            .I(\c0.data_out_9_7 ));
    LocalMux I__7304 (
            .O(N__34715),
            .I(\c0.data_out_9_7 ));
    InMux I__7303 (
            .O(N__34710),
            .I(N__34707));
    LocalMux I__7302 (
            .O(N__34707),
            .I(\c0.n17774 ));
    CascadeMux I__7301 (
            .O(N__34704),
            .I(\c0.n17774_cascade_ ));
    InMux I__7300 (
            .O(N__34701),
            .I(N__34691));
    InMux I__7299 (
            .O(N__34700),
            .I(N__34691));
    InMux I__7298 (
            .O(N__34699),
            .I(N__34691));
    InMux I__7297 (
            .O(N__34698),
            .I(N__34688));
    LocalMux I__7296 (
            .O(N__34691),
            .I(\c0.data_out_10_3 ));
    LocalMux I__7295 (
            .O(N__34688),
            .I(\c0.data_out_10_3 ));
    InMux I__7294 (
            .O(N__34683),
            .I(N__34680));
    LocalMux I__7293 (
            .O(N__34680),
            .I(N__34674));
    InMux I__7292 (
            .O(N__34679),
            .I(N__34669));
    InMux I__7291 (
            .O(N__34678),
            .I(N__34669));
    InMux I__7290 (
            .O(N__34677),
            .I(N__34666));
    Span4Mux_h I__7289 (
            .O(N__34674),
            .I(N__34661));
    LocalMux I__7288 (
            .O(N__34669),
            .I(N__34661));
    LocalMux I__7287 (
            .O(N__34666),
            .I(\c0.data_out_10_5 ));
    Odrv4 I__7286 (
            .O(N__34661),
            .I(\c0.data_out_10_5 ));
    InMux I__7285 (
            .O(N__34656),
            .I(N__34653));
    LocalMux I__7284 (
            .O(N__34653),
            .I(N__34650));
    Odrv4 I__7283 (
            .O(N__34650),
            .I(\c0.n6_adj_2314 ));
    InMux I__7282 (
            .O(N__34647),
            .I(N__34641));
    InMux I__7281 (
            .O(N__34646),
            .I(N__34641));
    LocalMux I__7280 (
            .O(N__34641),
            .I(N__34638));
    Odrv12 I__7279 (
            .O(N__34638),
            .I(\c0.n17883 ));
    CascadeMux I__7278 (
            .O(N__34635),
            .I(\c0.n10801_cascade_ ));
    InMux I__7277 (
            .O(N__34632),
            .I(N__34627));
    InMux I__7276 (
            .O(N__34631),
            .I(N__34624));
    InMux I__7275 (
            .O(N__34630),
            .I(N__34621));
    LocalMux I__7274 (
            .O(N__34627),
            .I(N__34618));
    LocalMux I__7273 (
            .O(N__34624),
            .I(N__34613));
    LocalMux I__7272 (
            .O(N__34621),
            .I(N__34613));
    Odrv4 I__7271 (
            .O(N__34618),
            .I(\c0.data_out_10_0 ));
    Odrv12 I__7270 (
            .O(N__34613),
            .I(\c0.data_out_10_0 ));
    InMux I__7269 (
            .O(N__34608),
            .I(N__34604));
    InMux I__7268 (
            .O(N__34607),
            .I(N__34601));
    LocalMux I__7267 (
            .O(N__34604),
            .I(\c0.n17768 ));
    LocalMux I__7266 (
            .O(N__34601),
            .I(\c0.n17768 ));
    CascadeMux I__7265 (
            .O(N__34596),
            .I(\c0.n10_adj_2366_cascade_ ));
    InMux I__7264 (
            .O(N__34593),
            .I(N__34585));
    InMux I__7263 (
            .O(N__34592),
            .I(N__34585));
    InMux I__7262 (
            .O(N__34591),
            .I(N__34582));
    InMux I__7261 (
            .O(N__34590),
            .I(N__34579));
    LocalMux I__7260 (
            .O(N__34585),
            .I(N__34576));
    LocalMux I__7259 (
            .O(N__34582),
            .I(\c0.data_out_10_1 ));
    LocalMux I__7258 (
            .O(N__34579),
            .I(\c0.data_out_10_1 ));
    Odrv4 I__7257 (
            .O(N__34576),
            .I(\c0.data_out_10_1 ));
    InMux I__7256 (
            .O(N__34569),
            .I(N__34566));
    LocalMux I__7255 (
            .O(N__34566),
            .I(N__34560));
    InMux I__7254 (
            .O(N__34565),
            .I(N__34557));
    InMux I__7253 (
            .O(N__34564),
            .I(N__34554));
    InMux I__7252 (
            .O(N__34563),
            .I(N__34551));
    Span4Mux_v I__7251 (
            .O(N__34560),
            .I(N__34542));
    LocalMux I__7250 (
            .O(N__34557),
            .I(N__34542));
    LocalMux I__7249 (
            .O(N__34554),
            .I(N__34542));
    LocalMux I__7248 (
            .O(N__34551),
            .I(N__34542));
    Span4Mux_h I__7247 (
            .O(N__34542),
            .I(N__34539));
    Odrv4 I__7246 (
            .O(N__34539),
            .I(\c0.data_out_6_1 ));
    CascadeMux I__7245 (
            .O(N__34536),
            .I(\c0.n6_adj_2318_cascade_ ));
    InMux I__7244 (
            .O(N__34533),
            .I(N__34529));
    InMux I__7243 (
            .O(N__34532),
            .I(N__34526));
    LocalMux I__7242 (
            .O(N__34529),
            .I(N__34520));
    LocalMux I__7241 (
            .O(N__34526),
            .I(N__34520));
    CascadeMux I__7240 (
            .O(N__34525),
            .I(N__34516));
    Span4Mux_v I__7239 (
            .O(N__34520),
            .I(N__34513));
    InMux I__7238 (
            .O(N__34519),
            .I(N__34510));
    InMux I__7237 (
            .O(N__34516),
            .I(N__34507));
    Span4Mux_h I__7236 (
            .O(N__34513),
            .I(N__34504));
    LocalMux I__7235 (
            .O(N__34510),
            .I(N__34499));
    LocalMux I__7234 (
            .O(N__34507),
            .I(N__34499));
    Odrv4 I__7233 (
            .O(N__34504),
            .I(\c0.data_out_9_0 ));
    Odrv12 I__7232 (
            .O(N__34499),
            .I(\c0.data_out_9_0 ));
    InMux I__7231 (
            .O(N__34494),
            .I(N__34489));
    CascadeMux I__7230 (
            .O(N__34493),
            .I(N__34486));
    InMux I__7229 (
            .O(N__34492),
            .I(N__34482));
    LocalMux I__7228 (
            .O(N__34489),
            .I(N__34479));
    InMux I__7227 (
            .O(N__34486),
            .I(N__34476));
    InMux I__7226 (
            .O(N__34485),
            .I(N__34473));
    LocalMux I__7225 (
            .O(N__34482),
            .I(N__34470));
    Span4Mux_h I__7224 (
            .O(N__34479),
            .I(N__34467));
    LocalMux I__7223 (
            .O(N__34476),
            .I(\c0.data_out_9_6 ));
    LocalMux I__7222 (
            .O(N__34473),
            .I(\c0.data_out_9_6 ));
    Odrv12 I__7221 (
            .O(N__34470),
            .I(\c0.data_out_9_6 ));
    Odrv4 I__7220 (
            .O(N__34467),
            .I(\c0.data_out_9_6 ));
    InMux I__7219 (
            .O(N__34458),
            .I(N__34455));
    LocalMux I__7218 (
            .O(N__34455),
            .I(\c0.n6_adj_2367 ));
    InMux I__7217 (
            .O(N__34452),
            .I(N__34449));
    LocalMux I__7216 (
            .O(N__34449),
            .I(\c0.n17850 ));
    CascadeMux I__7215 (
            .O(N__34446),
            .I(N__34443));
    InMux I__7214 (
            .O(N__34443),
            .I(N__34440));
    LocalMux I__7213 (
            .O(N__34440),
            .I(N__34436));
    InMux I__7212 (
            .O(N__34439),
            .I(N__34433));
    Span4Mux_v I__7211 (
            .O(N__34436),
            .I(N__34428));
    LocalMux I__7210 (
            .O(N__34433),
            .I(N__34428));
    Odrv4 I__7209 (
            .O(N__34428),
            .I(\c0.n10749 ));
    CascadeMux I__7208 (
            .O(N__34425),
            .I(\c0.data_out_9__2__N_367_cascade_ ));
    CascadeMux I__7207 (
            .O(N__34422),
            .I(\c0.n15_adj_2319_cascade_ ));
    InMux I__7206 (
            .O(N__34419),
            .I(N__34416));
    LocalMux I__7205 (
            .O(N__34416),
            .I(N__34413));
    Odrv4 I__7204 (
            .O(N__34413),
            .I(\c0.n14_adj_2320 ));
    InMux I__7203 (
            .O(N__34410),
            .I(N__34405));
    InMux I__7202 (
            .O(N__34409),
            .I(N__34400));
    InMux I__7201 (
            .O(N__34408),
            .I(N__34400));
    LocalMux I__7200 (
            .O(N__34405),
            .I(\c0.data_out_10_2 ));
    LocalMux I__7199 (
            .O(N__34400),
            .I(\c0.data_out_10_2 ));
    InMux I__7198 (
            .O(N__34395),
            .I(N__34389));
    InMux I__7197 (
            .O(N__34394),
            .I(N__34389));
    LocalMux I__7196 (
            .O(N__34389),
            .I(N__34386));
    Odrv4 I__7195 (
            .O(N__34386),
            .I(\c0.n17826 ));
    CascadeMux I__7194 (
            .O(N__34383),
            .I(\c0.n17761_cascade_ ));
    InMux I__7193 (
            .O(N__34380),
            .I(N__34377));
    LocalMux I__7192 (
            .O(N__34377),
            .I(N__34373));
    InMux I__7191 (
            .O(N__34376),
            .I(N__34370));
    Odrv4 I__7190 (
            .O(N__34373),
            .I(n9_adj_2477));
    LocalMux I__7189 (
            .O(N__34370),
            .I(n9_adj_2477));
    InMux I__7188 (
            .O(N__34365),
            .I(N__34362));
    LocalMux I__7187 (
            .O(N__34362),
            .I(\c0.n17761 ));
    InMux I__7186 (
            .O(N__34359),
            .I(N__34356));
    LocalMux I__7185 (
            .O(N__34356),
            .I(N__34353));
    Odrv4 I__7184 (
            .O(N__34353),
            .I(\c0.n18747 ));
    CascadeMux I__7183 (
            .O(N__34350),
            .I(\c0.n17807_cascade_ ));
    InMux I__7182 (
            .O(N__34347),
            .I(N__34344));
    LocalMux I__7181 (
            .O(N__34344),
            .I(N__34338));
    InMux I__7180 (
            .O(N__34343),
            .I(N__34333));
    InMux I__7179 (
            .O(N__34342),
            .I(N__34328));
    InMux I__7178 (
            .O(N__34341),
            .I(N__34328));
    Span4Mux_h I__7177 (
            .O(N__34338),
            .I(N__34325));
    InMux I__7176 (
            .O(N__34337),
            .I(N__34322));
    InMux I__7175 (
            .O(N__34336),
            .I(N__34319));
    LocalMux I__7174 (
            .O(N__34333),
            .I(data_out_9_2));
    LocalMux I__7173 (
            .O(N__34328),
            .I(data_out_9_2));
    Odrv4 I__7172 (
            .O(N__34325),
            .I(data_out_9_2));
    LocalMux I__7171 (
            .O(N__34322),
            .I(data_out_9_2));
    LocalMux I__7170 (
            .O(N__34319),
            .I(data_out_9_2));
    InMux I__7169 (
            .O(N__34308),
            .I(N__34305));
    LocalMux I__7168 (
            .O(N__34305),
            .I(N__34302));
    Span4Mux_h I__7167 (
            .O(N__34302),
            .I(N__34298));
    InMux I__7166 (
            .O(N__34301),
            .I(N__34294));
    Span4Mux_h I__7165 (
            .O(N__34298),
            .I(N__34291));
    InMux I__7164 (
            .O(N__34297),
            .I(N__34288));
    LocalMux I__7163 (
            .O(N__34294),
            .I(data_in_3_1));
    Odrv4 I__7162 (
            .O(N__34291),
            .I(data_in_3_1));
    LocalMux I__7161 (
            .O(N__34288),
            .I(data_in_3_1));
    InMux I__7160 (
            .O(N__34281),
            .I(N__34277));
    InMux I__7159 (
            .O(N__34280),
            .I(N__34274));
    LocalMux I__7158 (
            .O(N__34277),
            .I(N__34268));
    LocalMux I__7157 (
            .O(N__34274),
            .I(N__34268));
    InMux I__7156 (
            .O(N__34273),
            .I(N__34265));
    Span4Mux_h I__7155 (
            .O(N__34268),
            .I(N__34262));
    LocalMux I__7154 (
            .O(N__34265),
            .I(data_in_2_1));
    Odrv4 I__7153 (
            .O(N__34262),
            .I(data_in_2_1));
    InMux I__7152 (
            .O(N__34257),
            .I(N__34254));
    LocalMux I__7151 (
            .O(N__34254),
            .I(N__34251));
    Span4Mux_h I__7150 (
            .O(N__34251),
            .I(N__34247));
    InMux I__7149 (
            .O(N__34250),
            .I(N__34243));
    Span4Mux_h I__7148 (
            .O(N__34247),
            .I(N__34240));
    InMux I__7147 (
            .O(N__34246),
            .I(N__34237));
    LocalMux I__7146 (
            .O(N__34243),
            .I(data_in_3_3));
    Odrv4 I__7145 (
            .O(N__34240),
            .I(data_in_3_3));
    LocalMux I__7144 (
            .O(N__34237),
            .I(data_in_3_3));
    InMux I__7143 (
            .O(N__34230),
            .I(N__34222));
    InMux I__7142 (
            .O(N__34229),
            .I(N__34222));
    CascadeMux I__7141 (
            .O(N__34228),
            .I(N__34213));
    InMux I__7140 (
            .O(N__34227),
            .I(N__34205));
    LocalMux I__7139 (
            .O(N__34222),
            .I(N__34202));
    CascadeMux I__7138 (
            .O(N__34221),
            .I(N__34199));
    InMux I__7137 (
            .O(N__34220),
            .I(N__34189));
    InMux I__7136 (
            .O(N__34219),
            .I(N__34172));
    InMux I__7135 (
            .O(N__34218),
            .I(N__34172));
    InMux I__7134 (
            .O(N__34217),
            .I(N__34172));
    InMux I__7133 (
            .O(N__34216),
            .I(N__34165));
    InMux I__7132 (
            .O(N__34213),
            .I(N__34165));
    InMux I__7131 (
            .O(N__34212),
            .I(N__34165));
    InMux I__7130 (
            .O(N__34211),
            .I(N__34156));
    InMux I__7129 (
            .O(N__34210),
            .I(N__34156));
    InMux I__7128 (
            .O(N__34209),
            .I(N__34156));
    InMux I__7127 (
            .O(N__34208),
            .I(N__34156));
    LocalMux I__7126 (
            .O(N__34205),
            .I(N__34153));
    Span4Mux_v I__7125 (
            .O(N__34202),
            .I(N__34150));
    InMux I__7124 (
            .O(N__34199),
            .I(N__34143));
    InMux I__7123 (
            .O(N__34198),
            .I(N__34143));
    InMux I__7122 (
            .O(N__34197),
            .I(N__34143));
    InMux I__7121 (
            .O(N__34196),
            .I(N__34132));
    InMux I__7120 (
            .O(N__34195),
            .I(N__34132));
    InMux I__7119 (
            .O(N__34194),
            .I(N__34132));
    InMux I__7118 (
            .O(N__34193),
            .I(N__34132));
    InMux I__7117 (
            .O(N__34192),
            .I(N__34132));
    LocalMux I__7116 (
            .O(N__34189),
            .I(N__34129));
    InMux I__7115 (
            .O(N__34188),
            .I(N__34123));
    InMux I__7114 (
            .O(N__34187),
            .I(N__34118));
    InMux I__7113 (
            .O(N__34186),
            .I(N__34118));
    InMux I__7112 (
            .O(N__34185),
            .I(N__34113));
    InMux I__7111 (
            .O(N__34184),
            .I(N__34113));
    InMux I__7110 (
            .O(N__34183),
            .I(N__34106));
    InMux I__7109 (
            .O(N__34182),
            .I(N__34106));
    InMux I__7108 (
            .O(N__34181),
            .I(N__34106));
    InMux I__7107 (
            .O(N__34180),
            .I(N__34101));
    InMux I__7106 (
            .O(N__34179),
            .I(N__34101));
    LocalMux I__7105 (
            .O(N__34172),
            .I(N__34098));
    LocalMux I__7104 (
            .O(N__34165),
            .I(N__34093));
    LocalMux I__7103 (
            .O(N__34156),
            .I(N__34093));
    Span4Mux_v I__7102 (
            .O(N__34153),
            .I(N__34090));
    Span4Mux_h I__7101 (
            .O(N__34150),
            .I(N__34087));
    LocalMux I__7100 (
            .O(N__34143),
            .I(N__34080));
    LocalMux I__7099 (
            .O(N__34132),
            .I(N__34080));
    Span4Mux_h I__7098 (
            .O(N__34129),
            .I(N__34080));
    InMux I__7097 (
            .O(N__34128),
            .I(N__34073));
    InMux I__7096 (
            .O(N__34127),
            .I(N__34073));
    InMux I__7095 (
            .O(N__34126),
            .I(N__34073));
    LocalMux I__7094 (
            .O(N__34123),
            .I(rx_data_ready));
    LocalMux I__7093 (
            .O(N__34118),
            .I(rx_data_ready));
    LocalMux I__7092 (
            .O(N__34113),
            .I(rx_data_ready));
    LocalMux I__7091 (
            .O(N__34106),
            .I(rx_data_ready));
    LocalMux I__7090 (
            .O(N__34101),
            .I(rx_data_ready));
    Odrv4 I__7089 (
            .O(N__34098),
            .I(rx_data_ready));
    Odrv4 I__7088 (
            .O(N__34093),
            .I(rx_data_ready));
    Odrv4 I__7087 (
            .O(N__34090),
            .I(rx_data_ready));
    Odrv4 I__7086 (
            .O(N__34087),
            .I(rx_data_ready));
    Odrv4 I__7085 (
            .O(N__34080),
            .I(rx_data_ready));
    LocalMux I__7084 (
            .O(N__34073),
            .I(rx_data_ready));
    InMux I__7083 (
            .O(N__34050),
            .I(N__34045));
    InMux I__7082 (
            .O(N__34049),
            .I(N__34042));
    InMux I__7081 (
            .O(N__34048),
            .I(N__34039));
    LocalMux I__7080 (
            .O(N__34045),
            .I(N__34036));
    LocalMux I__7079 (
            .O(N__34042),
            .I(N__34033));
    LocalMux I__7078 (
            .O(N__34039),
            .I(N__34030));
    Span4Mux_v I__7077 (
            .O(N__34036),
            .I(N__34024));
    Span4Mux_h I__7076 (
            .O(N__34033),
            .I(N__34024));
    Span4Mux_v I__7075 (
            .O(N__34030),
            .I(N__34021));
    InMux I__7074 (
            .O(N__34029),
            .I(N__34018));
    Span4Mux_h I__7073 (
            .O(N__34024),
            .I(N__34013));
    Span4Mux_h I__7072 (
            .O(N__34021),
            .I(N__34013));
    LocalMux I__7071 (
            .O(N__34018),
            .I(data_in_2_3));
    Odrv4 I__7070 (
            .O(N__34013),
            .I(data_in_2_3));
    InMux I__7069 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__7068 (
            .O(N__34005),
            .I(N__34002));
    Odrv4 I__7067 (
            .O(N__34002),
            .I(\c0.n18365 ));
    InMux I__7066 (
            .O(N__33999),
            .I(N__33996));
    LocalMux I__7065 (
            .O(N__33996),
            .I(N__33993));
    Span4Mux_s1_v I__7064 (
            .O(N__33993),
            .I(N__33990));
    Span4Mux_v I__7063 (
            .O(N__33990),
            .I(N__33986));
    InMux I__7062 (
            .O(N__33989),
            .I(N__33983));
    Span4Mux_v I__7061 (
            .O(N__33986),
            .I(N__33980));
    LocalMux I__7060 (
            .O(N__33983),
            .I(data_out_frame2_18_5));
    Odrv4 I__7059 (
            .O(N__33980),
            .I(data_out_frame2_18_5));
    InMux I__7058 (
            .O(N__33975),
            .I(N__33972));
    LocalMux I__7057 (
            .O(N__33972),
            .I(n1));
    InMux I__7056 (
            .O(N__33969),
            .I(N__33966));
    LocalMux I__7055 (
            .O(N__33966),
            .I(N__33963));
    Span4Mux_h I__7054 (
            .O(N__33963),
            .I(N__33960));
    Odrv4 I__7053 (
            .O(N__33960),
            .I(n24_adj_2523));
    InMux I__7052 (
            .O(N__33957),
            .I(N__33954));
    LocalMux I__7051 (
            .O(N__33954),
            .I(n18_adj_2526));
    InMux I__7050 (
            .O(N__33951),
            .I(N__33948));
    LocalMux I__7049 (
            .O(N__33948),
            .I(N__33945));
    Odrv4 I__7048 (
            .O(N__33945),
            .I(\c0.n5_adj_2436 ));
    InMux I__7047 (
            .O(N__33942),
            .I(N__33931));
    InMux I__7046 (
            .O(N__33941),
            .I(N__33931));
    InMux I__7045 (
            .O(N__33940),
            .I(N__33928));
    InMux I__7044 (
            .O(N__33939),
            .I(N__33925));
    InMux I__7043 (
            .O(N__33938),
            .I(N__33918));
    InMux I__7042 (
            .O(N__33937),
            .I(N__33918));
    InMux I__7041 (
            .O(N__33936),
            .I(N__33918));
    LocalMux I__7040 (
            .O(N__33931),
            .I(N__33915));
    LocalMux I__7039 (
            .O(N__33928),
            .I(N__33911));
    LocalMux I__7038 (
            .O(N__33925),
            .I(N__33906));
    LocalMux I__7037 (
            .O(N__33918),
            .I(N__33906));
    Span4Mux_h I__7036 (
            .O(N__33915),
            .I(N__33903));
    InMux I__7035 (
            .O(N__33914),
            .I(N__33900));
    Span4Mux_h I__7034 (
            .O(N__33911),
            .I(N__33895));
    Span4Mux_v I__7033 (
            .O(N__33906),
            .I(N__33895));
    Span4Mux_h I__7032 (
            .O(N__33903),
            .I(N__33892));
    LocalMux I__7031 (
            .O(N__33900),
            .I(r_Bit_Index_0_adj_2519));
    Odrv4 I__7030 (
            .O(N__33895),
            .I(r_Bit_Index_0_adj_2519));
    Odrv4 I__7029 (
            .O(N__33892),
            .I(r_Bit_Index_0_adj_2519));
    InMux I__7028 (
            .O(N__33885),
            .I(N__33877));
    InMux I__7027 (
            .O(N__33884),
            .I(N__33877));
    InMux I__7026 (
            .O(N__33883),
            .I(N__33874));
    InMux I__7025 (
            .O(N__33882),
            .I(N__33871));
    LocalMux I__7024 (
            .O(N__33877),
            .I(N__33866));
    LocalMux I__7023 (
            .O(N__33874),
            .I(N__33866));
    LocalMux I__7022 (
            .O(N__33871),
            .I(N__33861));
    Span4Mux_v I__7021 (
            .O(N__33866),
            .I(N__33861));
    Odrv4 I__7020 (
            .O(N__33861),
            .I(r_Bit_Index_1_adj_2518));
    CascadeMux I__7019 (
            .O(N__33858),
            .I(N__33854));
    InMux I__7018 (
            .O(N__33857),
            .I(N__33847));
    InMux I__7017 (
            .O(N__33854),
            .I(N__33844));
    InMux I__7016 (
            .O(N__33853),
            .I(N__33835));
    InMux I__7015 (
            .O(N__33852),
            .I(N__33835));
    InMux I__7014 (
            .O(N__33851),
            .I(N__33835));
    InMux I__7013 (
            .O(N__33850),
            .I(N__33835));
    LocalMux I__7012 (
            .O(N__33847),
            .I(N__33831));
    LocalMux I__7011 (
            .O(N__33844),
            .I(N__33826));
    LocalMux I__7010 (
            .O(N__33835),
            .I(N__33826));
    InMux I__7009 (
            .O(N__33834),
            .I(N__33823));
    Span4Mux_h I__7008 (
            .O(N__33831),
            .I(N__33818));
    Span4Mux_h I__7007 (
            .O(N__33826),
            .I(N__33818));
    LocalMux I__7006 (
            .O(N__33823),
            .I(tx_transmit_N_1947_3));
    Odrv4 I__7005 (
            .O(N__33818),
            .I(tx_transmit_N_1947_3));
    InMux I__7004 (
            .O(N__33813),
            .I(N__33810));
    LocalMux I__7003 (
            .O(N__33810),
            .I(N__33807));
    Span4Mux_h I__7002 (
            .O(N__33807),
            .I(N__33803));
    InMux I__7001 (
            .O(N__33806),
            .I(N__33800));
    Odrv4 I__7000 (
            .O(N__33803),
            .I(\c0.n85 ));
    LocalMux I__6999 (
            .O(N__33800),
            .I(\c0.n85 ));
    InMux I__6998 (
            .O(N__33795),
            .I(N__33791));
    InMux I__6997 (
            .O(N__33794),
            .I(N__33784));
    LocalMux I__6996 (
            .O(N__33791),
            .I(N__33781));
    InMux I__6995 (
            .O(N__33790),
            .I(N__33772));
    InMux I__6994 (
            .O(N__33789),
            .I(N__33772));
    InMux I__6993 (
            .O(N__33788),
            .I(N__33772));
    InMux I__6992 (
            .O(N__33787),
            .I(N__33772));
    LocalMux I__6991 (
            .O(N__33784),
            .I(\c0.n14068 ));
    Odrv4 I__6990 (
            .O(N__33781),
            .I(\c0.n14068 ));
    LocalMux I__6989 (
            .O(N__33772),
            .I(\c0.n14068 ));
    InMux I__6988 (
            .O(N__33765),
            .I(N__33762));
    LocalMux I__6987 (
            .O(N__33762),
            .I(N__33759));
    Span4Mux_v I__6986 (
            .O(N__33759),
            .I(N__33756));
    Odrv4 I__6985 (
            .O(N__33756),
            .I(\c0.n18259 ));
    CascadeMux I__6984 (
            .O(N__33753),
            .I(N__33749));
    InMux I__6983 (
            .O(N__33752),
            .I(N__33743));
    InMux I__6982 (
            .O(N__33749),
            .I(N__33743));
    InMux I__6981 (
            .O(N__33748),
            .I(N__33740));
    LocalMux I__6980 (
            .O(N__33743),
            .I(N__33737));
    LocalMux I__6979 (
            .O(N__33740),
            .I(N__33734));
    Span4Mux_v I__6978 (
            .O(N__33737),
            .I(N__33731));
    Span4Mux_v I__6977 (
            .O(N__33734),
            .I(N__33728));
    Odrv4 I__6976 (
            .O(N__33731),
            .I(n18014));
    Odrv4 I__6975 (
            .O(N__33728),
            .I(n18014));
    CascadeMux I__6974 (
            .O(N__33723),
            .I(N__33720));
    InMux I__6973 (
            .O(N__33720),
            .I(N__33717));
    LocalMux I__6972 (
            .O(N__33717),
            .I(N__33714));
    Span4Mux_h I__6971 (
            .O(N__33714),
            .I(N__33711));
    Odrv4 I__6970 (
            .O(N__33711),
            .I(n4_adj_2472));
    InMux I__6969 (
            .O(N__33708),
            .I(N__33701));
    InMux I__6968 (
            .O(N__33707),
            .I(N__33701));
    InMux I__6967 (
            .O(N__33706),
            .I(N__33698));
    LocalMux I__6966 (
            .O(N__33701),
            .I(N__33695));
    LocalMux I__6965 (
            .O(N__33698),
            .I(N__33692));
    Span4Mux_v I__6964 (
            .O(N__33695),
            .I(N__33689));
    Span4Mux_v I__6963 (
            .O(N__33692),
            .I(N__33686));
    Odrv4 I__6962 (
            .O(N__33689),
            .I(n11545));
    Odrv4 I__6961 (
            .O(N__33686),
            .I(n11545));
    CascadeMux I__6960 (
            .O(N__33681),
            .I(N__33676));
    InMux I__6959 (
            .O(N__33680),
            .I(N__33673));
    InMux I__6958 (
            .O(N__33679),
            .I(N__33668));
    InMux I__6957 (
            .O(N__33676),
            .I(N__33668));
    LocalMux I__6956 (
            .O(N__33673),
            .I(N__33664));
    LocalMux I__6955 (
            .O(N__33668),
            .I(N__33661));
    InMux I__6954 (
            .O(N__33667),
            .I(N__33658));
    Span4Mux_v I__6953 (
            .O(N__33664),
            .I(N__33655));
    Span4Mux_h I__6952 (
            .O(N__33661),
            .I(N__33652));
    LocalMux I__6951 (
            .O(N__33658),
            .I(r_Bit_Index_2_adj_2517));
    Odrv4 I__6950 (
            .O(N__33655),
            .I(r_Bit_Index_2_adj_2517));
    Odrv4 I__6949 (
            .O(N__33652),
            .I(r_Bit_Index_2_adj_2517));
    InMux I__6948 (
            .O(N__33645),
            .I(N__33641));
    InMux I__6947 (
            .O(N__33644),
            .I(N__33638));
    LocalMux I__6946 (
            .O(N__33641),
            .I(N__33635));
    LocalMux I__6945 (
            .O(N__33638),
            .I(N__33632));
    Span4Mux_s2_v I__6944 (
            .O(N__33635),
            .I(N__33629));
    Span12Mux_s8_v I__6943 (
            .O(N__33632),
            .I(N__33626));
    Span4Mux_v I__6942 (
            .O(N__33629),
            .I(N__33623));
    Odrv12 I__6941 (
            .O(N__33626),
            .I(\c0.n17715 ));
    Odrv4 I__6940 (
            .O(N__33623),
            .I(\c0.n17715 ));
    InMux I__6939 (
            .O(N__33618),
            .I(N__33614));
    InMux I__6938 (
            .O(N__33617),
            .I(N__33611));
    LocalMux I__6937 (
            .O(N__33614),
            .I(N__33608));
    LocalMux I__6936 (
            .O(N__33611),
            .I(\c0.delay_counter_3 ));
    Odrv4 I__6935 (
            .O(N__33608),
            .I(\c0.delay_counter_3 ));
    InMux I__6934 (
            .O(N__33603),
            .I(N__33599));
    InMux I__6933 (
            .O(N__33602),
            .I(N__33596));
    LocalMux I__6932 (
            .O(N__33599),
            .I(\c0.delay_counter_8 ));
    LocalMux I__6931 (
            .O(N__33596),
            .I(\c0.delay_counter_8 ));
    InMux I__6930 (
            .O(N__33591),
            .I(N__33588));
    LocalMux I__6929 (
            .O(N__33588),
            .I(\c0.n18 ));
    InMux I__6928 (
            .O(N__33585),
            .I(N__33581));
    InMux I__6927 (
            .O(N__33584),
            .I(N__33578));
    LocalMux I__6926 (
            .O(N__33581),
            .I(\c0.delay_counter_10 ));
    LocalMux I__6925 (
            .O(N__33578),
            .I(\c0.delay_counter_10 ));
    CascadeMux I__6924 (
            .O(N__33573),
            .I(N__33570));
    InMux I__6923 (
            .O(N__33570),
            .I(N__33566));
    InMux I__6922 (
            .O(N__33569),
            .I(N__33563));
    LocalMux I__6921 (
            .O(N__33566),
            .I(\c0.delay_counter_0 ));
    LocalMux I__6920 (
            .O(N__33563),
            .I(\c0.delay_counter_0 ));
    CascadeMux I__6919 (
            .O(N__33558),
            .I(N__33554));
    InMux I__6918 (
            .O(N__33557),
            .I(N__33551));
    InMux I__6917 (
            .O(N__33554),
            .I(N__33548));
    LocalMux I__6916 (
            .O(N__33551),
            .I(\c0.delay_counter_13 ));
    LocalMux I__6915 (
            .O(N__33548),
            .I(\c0.delay_counter_13 ));
    InMux I__6914 (
            .O(N__33543),
            .I(N__33539));
    InMux I__6913 (
            .O(N__33542),
            .I(N__33536));
    LocalMux I__6912 (
            .O(N__33539),
            .I(\c0.delay_counter_6 ));
    LocalMux I__6911 (
            .O(N__33536),
            .I(\c0.delay_counter_6 ));
    InMux I__6910 (
            .O(N__33531),
            .I(N__33528));
    LocalMux I__6909 (
            .O(N__33528),
            .I(N__33525));
    Span4Mux_s2_v I__6908 (
            .O(N__33525),
            .I(N__33522));
    Span4Mux_v I__6907 (
            .O(N__33522),
            .I(N__33519));
    Odrv4 I__6906 (
            .O(N__33519),
            .I(\c0.n18810 ));
    InMux I__6905 (
            .O(N__33516),
            .I(N__33511));
    InMux I__6904 (
            .O(N__33515),
            .I(N__33508));
    InMux I__6903 (
            .O(N__33514),
            .I(N__33505));
    LocalMux I__6902 (
            .O(N__33511),
            .I(N__33502));
    LocalMux I__6901 (
            .O(N__33508),
            .I(N__33497));
    LocalMux I__6900 (
            .O(N__33505),
            .I(N__33497));
    Odrv4 I__6899 (
            .O(N__33502),
            .I(\c0.tx_transmit_N_1947_0 ));
    Odrv4 I__6898 (
            .O(N__33497),
            .I(\c0.tx_transmit_N_1947_0 ));
    InMux I__6897 (
            .O(N__33492),
            .I(N__33487));
    InMux I__6896 (
            .O(N__33491),
            .I(N__33484));
    InMux I__6895 (
            .O(N__33490),
            .I(N__33481));
    LocalMux I__6894 (
            .O(N__33487),
            .I(N__33478));
    LocalMux I__6893 (
            .O(N__33484),
            .I(\c0.tx_transmit_N_1947_1 ));
    LocalMux I__6892 (
            .O(N__33481),
            .I(\c0.tx_transmit_N_1947_1 ));
    Odrv4 I__6891 (
            .O(N__33478),
            .I(\c0.tx_transmit_N_1947_1 ));
    InMux I__6890 (
            .O(N__33471),
            .I(N__33466));
    InMux I__6889 (
            .O(N__33470),
            .I(N__33463));
    InMux I__6888 (
            .O(N__33469),
            .I(N__33460));
    LocalMux I__6887 (
            .O(N__33466),
            .I(N__33457));
    LocalMux I__6886 (
            .O(N__33463),
            .I(\c0.tx_transmit_N_1947_2 ));
    LocalMux I__6885 (
            .O(N__33460),
            .I(\c0.tx_transmit_N_1947_2 ));
    Odrv4 I__6884 (
            .O(N__33457),
            .I(\c0.tx_transmit_N_1947_2 ));
    InMux I__6883 (
            .O(N__33450),
            .I(N__33447));
    LocalMux I__6882 (
            .O(N__33447),
            .I(N__33442));
    InMux I__6881 (
            .O(N__33446),
            .I(N__33437));
    InMux I__6880 (
            .O(N__33445),
            .I(N__33437));
    Odrv4 I__6879 (
            .O(N__33442),
            .I(\c0.n155 ));
    LocalMux I__6878 (
            .O(N__33437),
            .I(\c0.n155 ));
    InMux I__6877 (
            .O(N__33432),
            .I(N__33428));
    InMux I__6876 (
            .O(N__33431),
            .I(N__33425));
    LocalMux I__6875 (
            .O(N__33428),
            .I(\c0.delay_counter_9 ));
    LocalMux I__6874 (
            .O(N__33425),
            .I(\c0.delay_counter_9 ));
    InMux I__6873 (
            .O(N__33420),
            .I(N__33416));
    InMux I__6872 (
            .O(N__33419),
            .I(N__33413));
    LocalMux I__6871 (
            .O(N__33416),
            .I(\c0.delay_counter_1 ));
    LocalMux I__6870 (
            .O(N__33413),
            .I(\c0.delay_counter_1 ));
    InMux I__6869 (
            .O(N__33408),
            .I(N__33405));
    LocalMux I__6868 (
            .O(N__33405),
            .I(\c0.n22 ));
    InMux I__6867 (
            .O(N__33402),
            .I(N__33399));
    LocalMux I__6866 (
            .O(N__33399),
            .I(N__33396));
    Span4Mux_h I__6865 (
            .O(N__33396),
            .I(N__33393));
    Odrv4 I__6864 (
            .O(N__33393),
            .I(n25_adj_2468));
    InMux I__6863 (
            .O(N__33390),
            .I(N__33387));
    LocalMux I__6862 (
            .O(N__33387),
            .I(\c0.n18807 ));
    InMux I__6861 (
            .O(N__33384),
            .I(N__33379));
    InMux I__6860 (
            .O(N__33383),
            .I(N__33376));
    InMux I__6859 (
            .O(N__33382),
            .I(N__33373));
    LocalMux I__6858 (
            .O(N__33379),
            .I(N__33369));
    LocalMux I__6857 (
            .O(N__33376),
            .I(N__33366));
    LocalMux I__6856 (
            .O(N__33373),
            .I(N__33363));
    InMux I__6855 (
            .O(N__33372),
            .I(N__33360));
    Span4Mux_v I__6854 (
            .O(N__33369),
            .I(N__33357));
    Span4Mux_h I__6853 (
            .O(N__33366),
            .I(N__33354));
    Odrv4 I__6852 (
            .O(N__33363),
            .I(data_out_frame2_6_7));
    LocalMux I__6851 (
            .O(N__33360),
            .I(data_out_frame2_6_7));
    Odrv4 I__6850 (
            .O(N__33357),
            .I(data_out_frame2_6_7));
    Odrv4 I__6849 (
            .O(N__33354),
            .I(data_out_frame2_6_7));
    InMux I__6848 (
            .O(N__33345),
            .I(N__33341));
    InMux I__6847 (
            .O(N__33344),
            .I(N__33338));
    LocalMux I__6846 (
            .O(N__33341),
            .I(data_out_frame2_18_0));
    LocalMux I__6845 (
            .O(N__33338),
            .I(data_out_frame2_18_0));
    InMux I__6844 (
            .O(N__33333),
            .I(N__33329));
    InMux I__6843 (
            .O(N__33332),
            .I(N__33325));
    LocalMux I__6842 (
            .O(N__33329),
            .I(N__33321));
    InMux I__6841 (
            .O(N__33328),
            .I(N__33317));
    LocalMux I__6840 (
            .O(N__33325),
            .I(N__33314));
    InMux I__6839 (
            .O(N__33324),
            .I(N__33311));
    Span4Mux_s2_v I__6838 (
            .O(N__33321),
            .I(N__33308));
    InMux I__6837 (
            .O(N__33320),
            .I(N__33305));
    LocalMux I__6836 (
            .O(N__33317),
            .I(data_out_frame2_12_1));
    Odrv4 I__6835 (
            .O(N__33314),
            .I(data_out_frame2_12_1));
    LocalMux I__6834 (
            .O(N__33311),
            .I(data_out_frame2_12_1));
    Odrv4 I__6833 (
            .O(N__33308),
            .I(data_out_frame2_12_1));
    LocalMux I__6832 (
            .O(N__33305),
            .I(data_out_frame2_12_1));
    CascadeMux I__6831 (
            .O(N__33294),
            .I(\c0.n10829_cascade_ ));
    InMux I__6830 (
            .O(N__33291),
            .I(N__33284));
    InMux I__6829 (
            .O(N__33290),
            .I(N__33284));
    InMux I__6828 (
            .O(N__33289),
            .I(N__33278));
    LocalMux I__6827 (
            .O(N__33284),
            .I(N__33274));
    InMux I__6826 (
            .O(N__33283),
            .I(N__33271));
    CascadeMux I__6825 (
            .O(N__33282),
            .I(N__33268));
    CascadeMux I__6824 (
            .O(N__33281),
            .I(N__33265));
    LocalMux I__6823 (
            .O(N__33278),
            .I(N__33260));
    CascadeMux I__6822 (
            .O(N__33277),
            .I(N__33256));
    Span4Mux_h I__6821 (
            .O(N__33274),
            .I(N__33250));
    LocalMux I__6820 (
            .O(N__33271),
            .I(N__33250));
    InMux I__6819 (
            .O(N__33268),
            .I(N__33241));
    InMux I__6818 (
            .O(N__33265),
            .I(N__33241));
    InMux I__6817 (
            .O(N__33264),
            .I(N__33241));
    InMux I__6816 (
            .O(N__33263),
            .I(N__33241));
    Span4Mux_v I__6815 (
            .O(N__33260),
            .I(N__33238));
    InMux I__6814 (
            .O(N__33259),
            .I(N__33230));
    InMux I__6813 (
            .O(N__33256),
            .I(N__33230));
    InMux I__6812 (
            .O(N__33255),
            .I(N__33230));
    Span4Mux_h I__6811 (
            .O(N__33250),
            .I(N__33225));
    LocalMux I__6810 (
            .O(N__33241),
            .I(N__33225));
    Span4Mux_v I__6809 (
            .O(N__33238),
            .I(N__33222));
    InMux I__6808 (
            .O(N__33237),
            .I(N__33219));
    LocalMux I__6807 (
            .O(N__33230),
            .I(N__33216));
    Span4Mux_h I__6806 (
            .O(N__33225),
            .I(N__33213));
    Sp12to4 I__6805 (
            .O(N__33222),
            .I(N__33210));
    LocalMux I__6804 (
            .O(N__33219),
            .I(N__33207));
    Span4Mux_h I__6803 (
            .O(N__33216),
            .I(N__33204));
    Span4Mux_v I__6802 (
            .O(N__33213),
            .I(N__33201));
    Odrv12 I__6801 (
            .O(N__33210),
            .I(\c0.FRAME_MATCHER_state_1 ));
    Odrv4 I__6800 (
            .O(N__33207),
            .I(\c0.FRAME_MATCHER_state_1 ));
    Odrv4 I__6799 (
            .O(N__33204),
            .I(\c0.FRAME_MATCHER_state_1 ));
    Odrv4 I__6798 (
            .O(N__33201),
            .I(\c0.FRAME_MATCHER_state_1 ));
    InMux I__6797 (
            .O(N__33192),
            .I(N__33189));
    LocalMux I__6796 (
            .O(N__33189),
            .I(N__33186));
    Odrv12 I__6795 (
            .O(N__33186),
            .I(\c0.n14161 ));
    CascadeMux I__6794 (
            .O(N__33183),
            .I(N__33171));
    InMux I__6793 (
            .O(N__33182),
            .I(N__33160));
    InMux I__6792 (
            .O(N__33181),
            .I(N__33160));
    InMux I__6791 (
            .O(N__33180),
            .I(N__33160));
    InMux I__6790 (
            .O(N__33179),
            .I(N__33160));
    InMux I__6789 (
            .O(N__33178),
            .I(N__33157));
    InMux I__6788 (
            .O(N__33177),
            .I(N__33154));
    InMux I__6787 (
            .O(N__33176),
            .I(N__33151));
    InMux I__6786 (
            .O(N__33175),
            .I(N__33146));
    InMux I__6785 (
            .O(N__33174),
            .I(N__33146));
    InMux I__6784 (
            .O(N__33171),
            .I(N__33143));
    InMux I__6783 (
            .O(N__33170),
            .I(N__33137));
    InMux I__6782 (
            .O(N__33169),
            .I(N__33137));
    LocalMux I__6781 (
            .O(N__33160),
            .I(N__33134));
    LocalMux I__6780 (
            .O(N__33157),
            .I(N__33131));
    LocalMux I__6779 (
            .O(N__33154),
            .I(N__33124));
    LocalMux I__6778 (
            .O(N__33151),
            .I(N__33124));
    LocalMux I__6777 (
            .O(N__33146),
            .I(N__33124));
    LocalMux I__6776 (
            .O(N__33143),
            .I(N__33121));
    InMux I__6775 (
            .O(N__33142),
            .I(N__33118));
    LocalMux I__6774 (
            .O(N__33137),
            .I(N__33113));
    Span4Mux_v I__6773 (
            .O(N__33134),
            .I(N__33113));
    Span4Mux_v I__6772 (
            .O(N__33131),
            .I(N__33108));
    Span4Mux_v I__6771 (
            .O(N__33124),
            .I(N__33108));
    Span12Mux_h I__6770 (
            .O(N__33121),
            .I(N__33103));
    LocalMux I__6769 (
            .O(N__33118),
            .I(N__33103));
    Span4Mux_h I__6768 (
            .O(N__33113),
            .I(N__33100));
    Span4Mux_h I__6767 (
            .O(N__33108),
            .I(N__33097));
    Odrv12 I__6766 (
            .O(N__33103),
            .I(\c0.FRAME_MATCHER_state_2 ));
    Odrv4 I__6765 (
            .O(N__33100),
            .I(\c0.FRAME_MATCHER_state_2 ));
    Odrv4 I__6764 (
            .O(N__33097),
            .I(\c0.FRAME_MATCHER_state_2 ));
    InMux I__6763 (
            .O(N__33090),
            .I(N__33084));
    InMux I__6762 (
            .O(N__33089),
            .I(N__33076));
    InMux I__6761 (
            .O(N__33088),
            .I(N__33076));
    InMux I__6760 (
            .O(N__33087),
            .I(N__33076));
    LocalMux I__6759 (
            .O(N__33084),
            .I(N__33073));
    InMux I__6758 (
            .O(N__33083),
            .I(N__33070));
    LocalMux I__6757 (
            .O(N__33076),
            .I(N__33067));
    Span4Mux_h I__6756 (
            .O(N__33073),
            .I(N__33062));
    LocalMux I__6755 (
            .O(N__33070),
            .I(N__33062));
    Span4Mux_s3_v I__6754 (
            .O(N__33067),
            .I(N__33052));
    Span4Mux_h I__6753 (
            .O(N__33062),
            .I(N__33052));
    InMux I__6752 (
            .O(N__33061),
            .I(N__33041));
    InMux I__6751 (
            .O(N__33060),
            .I(N__33041));
    InMux I__6750 (
            .O(N__33059),
            .I(N__33041));
    InMux I__6749 (
            .O(N__33058),
            .I(N__33041));
    InMux I__6748 (
            .O(N__33057),
            .I(N__33041));
    Span4Mux_h I__6747 (
            .O(N__33052),
            .I(N__33038));
    LocalMux I__6746 (
            .O(N__33041),
            .I(\c0.n50 ));
    Odrv4 I__6745 (
            .O(N__33038),
            .I(\c0.n50 ));
    CascadeMux I__6744 (
            .O(N__33033),
            .I(n11114_cascade_));
    InMux I__6743 (
            .O(N__33030),
            .I(N__33027));
    LocalMux I__6742 (
            .O(N__33027),
            .I(\c0.n17874 ));
    InMux I__6741 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__6740 (
            .O(N__33021),
            .I(\c0.n17908 ));
    InMux I__6739 (
            .O(N__33018),
            .I(N__33015));
    LocalMux I__6738 (
            .O(N__33015),
            .I(N__33012));
    Odrv12 I__6737 (
            .O(N__33012),
            .I(\c0.n18_adj_2423 ));
    CascadeMux I__6736 (
            .O(N__33009),
            .I(\c0.n17908_cascade_ ));
    InMux I__6735 (
            .O(N__33006),
            .I(N__33003));
    LocalMux I__6734 (
            .O(N__33003),
            .I(\c0.n28_adj_2425 ));
    CascadeMux I__6733 (
            .O(N__33000),
            .I(\c0.n30_adj_2424_cascade_ ));
    InMux I__6732 (
            .O(N__32997),
            .I(N__32994));
    LocalMux I__6731 (
            .O(N__32994),
            .I(\c0.n29_adj_2427 ));
    InMux I__6730 (
            .O(N__32991),
            .I(N__32988));
    LocalMux I__6729 (
            .O(N__32988),
            .I(N__32985));
    Span4Mux_s2_v I__6728 (
            .O(N__32985),
            .I(N__32981));
    InMux I__6727 (
            .O(N__32984),
            .I(N__32978));
    Span4Mux_h I__6726 (
            .O(N__32981),
            .I(N__32975));
    LocalMux I__6725 (
            .O(N__32978),
            .I(data_out_frame2_17_5));
    Odrv4 I__6724 (
            .O(N__32975),
            .I(data_out_frame2_17_5));
    CascadeMux I__6723 (
            .O(N__32970),
            .I(\c0.n18639_cascade_ ));
    CascadeMux I__6722 (
            .O(N__32967),
            .I(\c0.n10700_cascade_ ));
    InMux I__6721 (
            .O(N__32964),
            .I(N__32961));
    LocalMux I__6720 (
            .O(N__32961),
            .I(\c0.n21 ));
    CascadeMux I__6719 (
            .O(N__32958),
            .I(N__32955));
    InMux I__6718 (
            .O(N__32955),
            .I(N__32952));
    LocalMux I__6717 (
            .O(N__32952),
            .I(\c0.n17804 ));
    CascadeMux I__6716 (
            .O(N__32949),
            .I(n11017_cascade_));
    InMux I__6715 (
            .O(N__32946),
            .I(N__32942));
    InMux I__6714 (
            .O(N__32945),
            .I(N__32939));
    LocalMux I__6713 (
            .O(N__32942),
            .I(data_out_0_0));
    LocalMux I__6712 (
            .O(N__32939),
            .I(data_out_0_0));
    InMux I__6711 (
            .O(N__32934),
            .I(N__32928));
    InMux I__6710 (
            .O(N__32933),
            .I(N__32928));
    LocalMux I__6709 (
            .O(N__32928),
            .I(data_out_3_4));
    InMux I__6708 (
            .O(N__32925),
            .I(N__32922));
    LocalMux I__6707 (
            .O(N__32922),
            .I(N__32918));
    InMux I__6706 (
            .O(N__32921),
            .I(N__32915));
    Span4Mux_v I__6705 (
            .O(N__32918),
            .I(N__32910));
    LocalMux I__6704 (
            .O(N__32915),
            .I(N__32910));
    Odrv4 I__6703 (
            .O(N__32910),
            .I(\control.PHASES_5_N_2152_1 ));
    InMux I__6702 (
            .O(N__32907),
            .I(N__32901));
    InMux I__6701 (
            .O(N__32906),
            .I(N__32897));
    InMux I__6700 (
            .O(N__32905),
            .I(N__32894));
    InMux I__6699 (
            .O(N__32904),
            .I(N__32891));
    LocalMux I__6698 (
            .O(N__32901),
            .I(N__32888));
    InMux I__6697 (
            .O(N__32900),
            .I(N__32885));
    LocalMux I__6696 (
            .O(N__32897),
            .I(N__32882));
    LocalMux I__6695 (
            .O(N__32894),
            .I(N__32877));
    LocalMux I__6694 (
            .O(N__32891),
            .I(N__32877));
    Span4Mux_v I__6693 (
            .O(N__32888),
            .I(N__32874));
    LocalMux I__6692 (
            .O(N__32885),
            .I(N__32867));
    Span4Mux_v I__6691 (
            .O(N__32882),
            .I(N__32867));
    Span4Mux_v I__6690 (
            .O(N__32877),
            .I(N__32867));
    Odrv4 I__6689 (
            .O(N__32874),
            .I(\control.pwm_delay_9 ));
    Odrv4 I__6688 (
            .O(N__32867),
            .I(\control.pwm_delay_9 ));
    InMux I__6687 (
            .O(N__32862),
            .I(N__32859));
    LocalMux I__6686 (
            .O(N__32859),
            .I(N__32853));
    InMux I__6685 (
            .O(N__32858),
            .I(N__32850));
    InMux I__6684 (
            .O(N__32857),
            .I(N__32847));
    InMux I__6683 (
            .O(N__32856),
            .I(N__32844));
    Sp12to4 I__6682 (
            .O(N__32853),
            .I(N__32839));
    LocalMux I__6681 (
            .O(N__32850),
            .I(N__32839));
    LocalMux I__6680 (
            .O(N__32847),
            .I(N__32834));
    LocalMux I__6679 (
            .O(N__32844),
            .I(N__32834));
    Span12Mux_s10_v I__6678 (
            .O(N__32839),
            .I(N__32831));
    Span12Mux_s10_v I__6677 (
            .O(N__32834),
            .I(N__32828));
    Odrv12 I__6676 (
            .O(N__32831),
            .I(\control.n18 ));
    Odrv12 I__6675 (
            .O(N__32828),
            .I(\control.n18 ));
    InMux I__6674 (
            .O(N__32823),
            .I(N__32820));
    LocalMux I__6673 (
            .O(N__32820),
            .I(\control.n17926 ));
    CascadeMux I__6672 (
            .O(N__32817),
            .I(\control.PHASES_5__N_2160_cascade_ ));
    InMux I__6671 (
            .O(N__32814),
            .I(N__32810));
    InMux I__6670 (
            .O(N__32813),
            .I(N__32807));
    LocalMux I__6669 (
            .O(N__32810),
            .I(\control.n5 ));
    LocalMux I__6668 (
            .O(N__32807),
            .I(\control.n5 ));
    CascadeMux I__6667 (
            .O(N__32802),
            .I(N__32799));
    InMux I__6666 (
            .O(N__32799),
            .I(N__32796));
    LocalMux I__6665 (
            .O(N__32796),
            .I(\control.n17950 ));
    CEMux I__6664 (
            .O(N__32793),
            .I(N__32790));
    LocalMux I__6663 (
            .O(N__32790),
            .I(N__32787));
    Span4Mux_s3_v I__6662 (
            .O(N__32787),
            .I(N__32784));
    Span4Mux_h I__6661 (
            .O(N__32784),
            .I(N__32781));
    Span4Mux_h I__6660 (
            .O(N__32781),
            .I(N__32778));
    Span4Mux_h I__6659 (
            .O(N__32778),
            .I(N__32775));
    Odrv4 I__6658 (
            .O(N__32775),
            .I(\control.n9 ));
    CascadeMux I__6657 (
            .O(N__32772),
            .I(\c0.n1_cascade_ ));
    CascadeMux I__6656 (
            .O(N__32769),
            .I(N__32766));
    InMux I__6655 (
            .O(N__32766),
            .I(N__32763));
    LocalMux I__6654 (
            .O(N__32763),
            .I(N__32760));
    Odrv12 I__6653 (
            .O(N__32760),
            .I(n22));
    InMux I__6652 (
            .O(N__32757),
            .I(N__32754));
    LocalMux I__6651 (
            .O(N__32754),
            .I(\c0.n18849 ));
    CascadeMux I__6650 (
            .O(N__32751),
            .I(n18852_cascade_));
    InMux I__6649 (
            .O(N__32748),
            .I(N__32745));
    LocalMux I__6648 (
            .O(N__32745),
            .I(n10));
    CascadeMux I__6647 (
            .O(N__32742),
            .I(N__32739));
    InMux I__6646 (
            .O(N__32739),
            .I(N__32736));
    LocalMux I__6645 (
            .O(N__32736),
            .I(\c0.n18264 ));
    CascadeMux I__6644 (
            .O(N__32733),
            .I(N__32730));
    InMux I__6643 (
            .O(N__32730),
            .I(N__32727));
    LocalMux I__6642 (
            .O(N__32727),
            .I(\c0.n8 ));
    InMux I__6641 (
            .O(N__32724),
            .I(N__32721));
    LocalMux I__6640 (
            .O(N__32721),
            .I(n10_adj_2527));
    InMux I__6639 (
            .O(N__32718),
            .I(N__32715));
    LocalMux I__6638 (
            .O(N__32715),
            .I(\c0.n18322 ));
    InMux I__6637 (
            .O(N__32712),
            .I(N__32708));
    InMux I__6636 (
            .O(N__32711),
            .I(N__32705));
    LocalMux I__6635 (
            .O(N__32708),
            .I(N__32702));
    LocalMux I__6634 (
            .O(N__32705),
            .I(data_out_0_1));
    Odrv12 I__6633 (
            .O(N__32702),
            .I(data_out_0_1));
    InMux I__6632 (
            .O(N__32697),
            .I(N__32694));
    LocalMux I__6631 (
            .O(N__32694),
            .I(\c0.n17742 ));
    CascadeMux I__6630 (
            .O(N__32691),
            .I(N__32688));
    InMux I__6629 (
            .O(N__32688),
            .I(N__32685));
    LocalMux I__6628 (
            .O(N__32685),
            .I(\c0.n10558 ));
    InMux I__6627 (
            .O(N__32682),
            .I(N__32678));
    InMux I__6626 (
            .O(N__32681),
            .I(N__32675));
    LocalMux I__6625 (
            .O(N__32678),
            .I(N__32671));
    LocalMux I__6624 (
            .O(N__32675),
            .I(N__32668));
    InMux I__6623 (
            .O(N__32674),
            .I(N__32665));
    Odrv4 I__6622 (
            .O(N__32671),
            .I(\c0.data_out_9_5 ));
    Odrv4 I__6621 (
            .O(N__32668),
            .I(\c0.data_out_9_5 ));
    LocalMux I__6620 (
            .O(N__32665),
            .I(\c0.data_out_9_5 ));
    CascadeMux I__6619 (
            .O(N__32658),
            .I(\c0.n6_adj_2365_cascade_ ));
    CascadeMux I__6618 (
            .O(N__32655),
            .I(N__32652));
    InMux I__6617 (
            .O(N__32652),
            .I(N__32649));
    LocalMux I__6616 (
            .O(N__32649),
            .I(\c0.n5_adj_2220 ));
    InMux I__6615 (
            .O(N__32646),
            .I(N__32642));
    CascadeMux I__6614 (
            .O(N__32645),
            .I(N__32639));
    LocalMux I__6613 (
            .O(N__32642),
            .I(N__32636));
    InMux I__6612 (
            .O(N__32639),
            .I(N__32633));
    Span4Mux_v I__6611 (
            .O(N__32636),
            .I(N__32630));
    LocalMux I__6610 (
            .O(N__32633),
            .I(r_Tx_Data_4));
    Odrv4 I__6609 (
            .O(N__32630),
            .I(r_Tx_Data_4));
    InMux I__6608 (
            .O(N__32625),
            .I(N__32622));
    LocalMux I__6607 (
            .O(N__32622),
            .I(\c0.n18265 ));
    CascadeMux I__6606 (
            .O(N__32619),
            .I(N__32615));
    InMux I__6605 (
            .O(N__32618),
            .I(N__32608));
    InMux I__6604 (
            .O(N__32615),
            .I(N__32608));
    InMux I__6603 (
            .O(N__32614),
            .I(N__32605));
    CascadeMux I__6602 (
            .O(N__32613),
            .I(N__32602));
    LocalMux I__6601 (
            .O(N__32608),
            .I(N__32595));
    LocalMux I__6600 (
            .O(N__32605),
            .I(N__32595));
    InMux I__6599 (
            .O(N__32602),
            .I(N__32592));
    InMux I__6598 (
            .O(N__32601),
            .I(N__32589));
    CascadeMux I__6597 (
            .O(N__32600),
            .I(N__32586));
    Span4Mux_v I__6596 (
            .O(N__32595),
            .I(N__32580));
    LocalMux I__6595 (
            .O(N__32592),
            .I(N__32580));
    LocalMux I__6594 (
            .O(N__32589),
            .I(N__32577));
    InMux I__6593 (
            .O(N__32586),
            .I(N__32574));
    InMux I__6592 (
            .O(N__32585),
            .I(N__32571));
    Span4Mux_v I__6591 (
            .O(N__32580),
            .I(N__32567));
    Span4Mux_h I__6590 (
            .O(N__32577),
            .I(N__32564));
    LocalMux I__6589 (
            .O(N__32574),
            .I(N__32561));
    LocalMux I__6588 (
            .O(N__32571),
            .I(N__32558));
    InMux I__6587 (
            .O(N__32570),
            .I(N__32555));
    Span4Mux_h I__6586 (
            .O(N__32567),
            .I(N__32552));
    Span4Mux_h I__6585 (
            .O(N__32564),
            .I(N__32549));
    Span4Mux_h I__6584 (
            .O(N__32561),
            .I(N__32542));
    Span4Mux_v I__6583 (
            .O(N__32558),
            .I(N__32542));
    LocalMux I__6582 (
            .O(N__32555),
            .I(N__32542));
    Odrv4 I__6581 (
            .O(N__32552),
            .I(n9667));
    Odrv4 I__6580 (
            .O(N__32549),
            .I(n9667));
    Odrv4 I__6579 (
            .O(N__32542),
            .I(n9667));
    InMux I__6578 (
            .O(N__32535),
            .I(N__32532));
    LocalMux I__6577 (
            .O(N__32532),
            .I(N__32526));
    InMux I__6576 (
            .O(N__32531),
            .I(N__32520));
    InMux I__6575 (
            .O(N__32530),
            .I(N__32517));
    InMux I__6574 (
            .O(N__32529),
            .I(N__32514));
    Span4Mux_v I__6573 (
            .O(N__32526),
            .I(N__32510));
    InMux I__6572 (
            .O(N__32525),
            .I(N__32507));
    InMux I__6571 (
            .O(N__32524),
            .I(N__32503));
    InMux I__6570 (
            .O(N__32523),
            .I(N__32500));
    LocalMux I__6569 (
            .O(N__32520),
            .I(N__32493));
    LocalMux I__6568 (
            .O(N__32517),
            .I(N__32493));
    LocalMux I__6567 (
            .O(N__32514),
            .I(N__32493));
    InMux I__6566 (
            .O(N__32513),
            .I(N__32490));
    Span4Mux_v I__6565 (
            .O(N__32510),
            .I(N__32485));
    LocalMux I__6564 (
            .O(N__32507),
            .I(N__32485));
    InMux I__6563 (
            .O(N__32506),
            .I(N__32481));
    LocalMux I__6562 (
            .O(N__32503),
            .I(N__32474));
    LocalMux I__6561 (
            .O(N__32500),
            .I(N__32474));
    Span4Mux_v I__6560 (
            .O(N__32493),
            .I(N__32474));
    LocalMux I__6559 (
            .O(N__32490),
            .I(N__32469));
    Span4Mux_v I__6558 (
            .O(N__32485),
            .I(N__32469));
    InMux I__6557 (
            .O(N__32484),
            .I(N__32466));
    LocalMux I__6556 (
            .O(N__32481),
            .I(byte_transmit_counter_4));
    Odrv4 I__6555 (
            .O(N__32474),
            .I(byte_transmit_counter_4));
    Odrv4 I__6554 (
            .O(N__32469),
            .I(byte_transmit_counter_4));
    LocalMux I__6553 (
            .O(N__32466),
            .I(byte_transmit_counter_4));
    InMux I__6552 (
            .O(N__32457),
            .I(N__32454));
    LocalMux I__6551 (
            .O(N__32454),
            .I(N__32450));
    InMux I__6550 (
            .O(N__32453),
            .I(N__32447));
    Span4Mux_v I__6549 (
            .O(N__32450),
            .I(N__32444));
    LocalMux I__6548 (
            .O(N__32447),
            .I(r_Tx_Data_0));
    Odrv4 I__6547 (
            .O(N__32444),
            .I(r_Tx_Data_0));
    InMux I__6546 (
            .O(N__32439),
            .I(N__32435));
    InMux I__6545 (
            .O(N__32438),
            .I(N__32432));
    LocalMux I__6544 (
            .O(N__32435),
            .I(N__32429));
    LocalMux I__6543 (
            .O(N__32432),
            .I(\c0.n10524 ));
    Odrv4 I__6542 (
            .O(N__32429),
            .I(\c0.n10524 ));
    InMux I__6541 (
            .O(N__32424),
            .I(N__32420));
    InMux I__6540 (
            .O(N__32423),
            .I(N__32417));
    LocalMux I__6539 (
            .O(N__32420),
            .I(\c0.n10550 ));
    LocalMux I__6538 (
            .O(N__32417),
            .I(\c0.n10550 ));
    InMux I__6537 (
            .O(N__32412),
            .I(N__32409));
    LocalMux I__6536 (
            .O(N__32409),
            .I(N__32406));
    Span4Mux_h I__6535 (
            .O(N__32406),
            .I(N__32403));
    Span4Mux_h I__6534 (
            .O(N__32403),
            .I(N__32400));
    Odrv4 I__6533 (
            .O(N__32400),
            .I(\c0.n10746 ));
    InMux I__6532 (
            .O(N__32397),
            .I(N__32394));
    LocalMux I__6531 (
            .O(N__32394),
            .I(\c0.n6_adj_2361 ));
    CascadeMux I__6530 (
            .O(N__32391),
            .I(\c0.n10746_cascade_ ));
    CascadeMux I__6529 (
            .O(N__32388),
            .I(n17758_cascade_));
    InMux I__6528 (
            .O(N__32385),
            .I(N__32382));
    LocalMux I__6527 (
            .O(N__32382),
            .I(\c0.n10734 ));
    CascadeMux I__6526 (
            .O(N__32379),
            .I(N__32376));
    InMux I__6525 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__6524 (
            .O(N__32373),
            .I(\c0.n8_adj_2232 ));
    CascadeMux I__6523 (
            .O(N__32370),
            .I(N__32367));
    InMux I__6522 (
            .O(N__32367),
            .I(N__32364));
    LocalMux I__6521 (
            .O(N__32364),
            .I(N__32361));
    Odrv4 I__6520 (
            .O(N__32361),
            .I(n10_adj_2461));
    InMux I__6519 (
            .O(N__32358),
            .I(N__32354));
    InMux I__6518 (
            .O(N__32357),
            .I(N__32349));
    LocalMux I__6517 (
            .O(N__32354),
            .I(N__32346));
    InMux I__6516 (
            .O(N__32353),
            .I(N__32343));
    InMux I__6515 (
            .O(N__32352),
            .I(N__32340));
    LocalMux I__6514 (
            .O(N__32349),
            .I(data_out_8_7));
    Odrv4 I__6513 (
            .O(N__32346),
            .I(data_out_8_7));
    LocalMux I__6512 (
            .O(N__32343),
            .I(data_out_8_7));
    LocalMux I__6511 (
            .O(N__32340),
            .I(data_out_8_7));
    CascadeMux I__6510 (
            .O(N__32331),
            .I(\c0.n17742_cascade_ ));
    CascadeMux I__6509 (
            .O(N__32328),
            .I(n18864_cascade_));
    CascadeMux I__6508 (
            .O(N__32325),
            .I(n10_adj_2529_cascade_));
    InMux I__6507 (
            .O(N__32322),
            .I(N__32318));
    InMux I__6506 (
            .O(N__32321),
            .I(N__32315));
    LocalMux I__6505 (
            .O(N__32318),
            .I(N__32312));
    LocalMux I__6504 (
            .O(N__32315),
            .I(r_Tx_Data_3));
    Odrv4 I__6503 (
            .O(N__32312),
            .I(r_Tx_Data_3));
    InMux I__6502 (
            .O(N__32307),
            .I(N__32304));
    LocalMux I__6501 (
            .O(N__32304),
            .I(n10_adj_2499));
    CascadeMux I__6500 (
            .O(N__32301),
            .I(\c0.n10550_cascade_ ));
    CascadeMux I__6499 (
            .O(N__32298),
            .I(n17978_cascade_));
    InMux I__6498 (
            .O(N__32295),
            .I(N__32288));
    InMux I__6497 (
            .O(N__32294),
            .I(N__32288));
    InMux I__6496 (
            .O(N__32293),
            .I(N__32285));
    LocalMux I__6495 (
            .O(N__32288),
            .I(UART_TRANSMITTER_state_7_N_1223_1));
    LocalMux I__6494 (
            .O(N__32285),
            .I(UART_TRANSMITTER_state_7_N_1223_1));
    InMux I__6493 (
            .O(N__32280),
            .I(N__32277));
    LocalMux I__6492 (
            .O(N__32277),
            .I(n18202));
    CascadeMux I__6491 (
            .O(N__32274),
            .I(N__32271));
    InMux I__6490 (
            .O(N__32271),
            .I(N__32265));
    InMux I__6489 (
            .O(N__32270),
            .I(N__32265));
    LocalMux I__6488 (
            .O(N__32265),
            .I(n574));
    InMux I__6487 (
            .O(N__32262),
            .I(N__32259));
    LocalMux I__6486 (
            .O(N__32259),
            .I(N__32253));
    InMux I__6485 (
            .O(N__32258),
            .I(N__32246));
    InMux I__6484 (
            .O(N__32257),
            .I(N__32246));
    InMux I__6483 (
            .O(N__32256),
            .I(N__32246));
    Odrv4 I__6482 (
            .O(N__32253),
            .I(n4));
    LocalMux I__6481 (
            .O(N__32246),
            .I(n4));
    InMux I__6480 (
            .O(N__32241),
            .I(N__32238));
    LocalMux I__6479 (
            .O(N__32238),
            .I(n22_adj_2522));
    CascadeMux I__6478 (
            .O(N__32235),
            .I(N__32232));
    InMux I__6477 (
            .O(N__32232),
            .I(N__32229));
    LocalMux I__6476 (
            .O(N__32229),
            .I(\c0.n18226 ));
    InMux I__6475 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__6474 (
            .O(N__32223),
            .I(n21_adj_2524));
    InMux I__6473 (
            .O(N__32220),
            .I(N__32217));
    LocalMux I__6472 (
            .O(N__32217),
            .I(n6_adj_2470));
    InMux I__6471 (
            .O(N__32214),
            .I(N__32211));
    LocalMux I__6470 (
            .O(N__32211),
            .I(n18368));
    CascadeMux I__6469 (
            .O(N__32208),
            .I(\c0.n18861_cascade_ ));
    InMux I__6468 (
            .O(N__32205),
            .I(N__32202));
    LocalMux I__6467 (
            .O(N__32202),
            .I(N__32199));
    Span4Mux_v I__6466 (
            .O(N__32199),
            .I(N__32196));
    Odrv4 I__6465 (
            .O(N__32196),
            .I(\c0.n18377 ));
    InMux I__6464 (
            .O(N__32193),
            .I(N__32190));
    LocalMux I__6463 (
            .O(N__32190),
            .I(\c0.n18019 ));
    InMux I__6462 (
            .O(N__32187),
            .I(N__32184));
    LocalMux I__6461 (
            .O(N__32184),
            .I(n129));
    InMux I__6460 (
            .O(N__32181),
            .I(N__32175));
    InMux I__6459 (
            .O(N__32180),
            .I(N__32172));
    InMux I__6458 (
            .O(N__32179),
            .I(N__32169));
    CascadeMux I__6457 (
            .O(N__32178),
            .I(N__32165));
    LocalMux I__6456 (
            .O(N__32175),
            .I(N__32161));
    LocalMux I__6455 (
            .O(N__32172),
            .I(N__32156));
    LocalMux I__6454 (
            .O(N__32169),
            .I(N__32156));
    InMux I__6453 (
            .O(N__32168),
            .I(N__32153));
    InMux I__6452 (
            .O(N__32165),
            .I(N__32148));
    InMux I__6451 (
            .O(N__32164),
            .I(N__32148));
    Odrv12 I__6450 (
            .O(N__32161),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    Odrv4 I__6449 (
            .O(N__32156),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    LocalMux I__6448 (
            .O(N__32153),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    LocalMux I__6447 (
            .O(N__32148),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    CascadeMux I__6446 (
            .O(N__32139),
            .I(n129_cascade_));
    InMux I__6445 (
            .O(N__32136),
            .I(N__32133));
    LocalMux I__6444 (
            .O(N__32133),
            .I(N__32126));
    InMux I__6443 (
            .O(N__32132),
            .I(N__32121));
    InMux I__6442 (
            .O(N__32131),
            .I(N__32121));
    InMux I__6441 (
            .O(N__32130),
            .I(N__32115));
    InMux I__6440 (
            .O(N__32129),
            .I(N__32115));
    Span4Mux_h I__6439 (
            .O(N__32126),
            .I(N__32112));
    LocalMux I__6438 (
            .O(N__32121),
            .I(N__32109));
    InMux I__6437 (
            .O(N__32120),
            .I(N__32106));
    LocalMux I__6436 (
            .O(N__32115),
            .I(\c0.tx_active ));
    Odrv4 I__6435 (
            .O(N__32112),
            .I(\c0.tx_active ));
    Odrv4 I__6434 (
            .O(N__32109),
            .I(\c0.tx_active ));
    LocalMux I__6433 (
            .O(N__32106),
            .I(\c0.tx_active ));
    InMux I__6432 (
            .O(N__32097),
            .I(N__32094));
    LocalMux I__6431 (
            .O(N__32094),
            .I(N__32091));
    Odrv4 I__6430 (
            .O(N__32091),
            .I(\c0.n1707 ));
    InMux I__6429 (
            .O(N__32088),
            .I(N__32084));
    InMux I__6428 (
            .O(N__32087),
            .I(N__32081));
    LocalMux I__6427 (
            .O(N__32084),
            .I(\c0.delay_counter_11 ));
    LocalMux I__6426 (
            .O(N__32081),
            .I(\c0.delay_counter_11 ));
    InMux I__6425 (
            .O(N__32076),
            .I(N__32072));
    InMux I__6424 (
            .O(N__32075),
            .I(N__32069));
    LocalMux I__6423 (
            .O(N__32072),
            .I(\c0.delay_counter_12 ));
    LocalMux I__6422 (
            .O(N__32069),
            .I(\c0.delay_counter_12 ));
    CascadeMux I__6421 (
            .O(N__32064),
            .I(N__32061));
    InMux I__6420 (
            .O(N__32061),
            .I(N__32057));
    InMux I__6419 (
            .O(N__32060),
            .I(N__32054));
    LocalMux I__6418 (
            .O(N__32057),
            .I(N__32051));
    LocalMux I__6417 (
            .O(N__32054),
            .I(\c0.delay_counter_4 ));
    Odrv12 I__6416 (
            .O(N__32051),
            .I(\c0.delay_counter_4 ));
    InMux I__6415 (
            .O(N__32046),
            .I(N__32042));
    InMux I__6414 (
            .O(N__32045),
            .I(N__32039));
    LocalMux I__6413 (
            .O(N__32042),
            .I(N__32036));
    LocalMux I__6412 (
            .O(N__32039),
            .I(\c0.delay_counter_7 ));
    Odrv4 I__6411 (
            .O(N__32036),
            .I(\c0.delay_counter_7 ));
    InMux I__6410 (
            .O(N__32031),
            .I(N__32028));
    LocalMux I__6409 (
            .O(N__32028),
            .I(\c0.n24 ));
    CascadeMux I__6408 (
            .O(N__32025),
            .I(N__32020));
    InMux I__6407 (
            .O(N__32024),
            .I(N__32016));
    InMux I__6406 (
            .O(N__32023),
            .I(N__32011));
    InMux I__6405 (
            .O(N__32020),
            .I(N__32011));
    InMux I__6404 (
            .O(N__32019),
            .I(N__32008));
    LocalMux I__6403 (
            .O(N__32016),
            .I(N__32003));
    LocalMux I__6402 (
            .O(N__32011),
            .I(N__32003));
    LocalMux I__6401 (
            .O(N__32008),
            .I(n12227));
    Odrv4 I__6400 (
            .O(N__32003),
            .I(n12227));
    CascadeMux I__6399 (
            .O(N__31998),
            .I(n574_cascade_));
    InMux I__6398 (
            .O(N__31995),
            .I(N__31992));
    LocalMux I__6397 (
            .O(N__31992),
            .I(\c0.n98 ));
    CascadeMux I__6396 (
            .O(N__31989),
            .I(N__31986));
    InMux I__6395 (
            .O(N__31986),
            .I(N__31983));
    LocalMux I__6394 (
            .O(N__31983),
            .I(N__31980));
    Span4Mux_v I__6393 (
            .O(N__31980),
            .I(N__31977));
    Odrv4 I__6392 (
            .O(N__31977),
            .I(\c0.n18230 ));
    InMux I__6391 (
            .O(N__31974),
            .I(\c0.n16640 ));
    InMux I__6390 (
            .O(N__31971),
            .I(bfn_11_8_0_));
    InMux I__6389 (
            .O(N__31968),
            .I(\c0.n16642 ));
    InMux I__6388 (
            .O(N__31965),
            .I(\c0.n16643 ));
    InMux I__6387 (
            .O(N__31962),
            .I(\c0.n16644 ));
    InMux I__6386 (
            .O(N__31959),
            .I(\c0.n16645 ));
    InMux I__6385 (
            .O(N__31956),
            .I(\c0.n16646 ));
    InMux I__6384 (
            .O(N__31953),
            .I(N__31949));
    InMux I__6383 (
            .O(N__31952),
            .I(N__31946));
    LocalMux I__6382 (
            .O(N__31949),
            .I(N__31943));
    LocalMux I__6381 (
            .O(N__31946),
            .I(\c0.delay_counter_2 ));
    Odrv12 I__6380 (
            .O(N__31943),
            .I(\c0.delay_counter_2 ));
    CascadeMux I__6379 (
            .O(N__31938),
            .I(N__31935));
    InMux I__6378 (
            .O(N__31935),
            .I(N__31931));
    InMux I__6377 (
            .O(N__31934),
            .I(N__31928));
    LocalMux I__6376 (
            .O(N__31931),
            .I(N__31925));
    LocalMux I__6375 (
            .O(N__31928),
            .I(\c0.delay_counter_5 ));
    Odrv4 I__6374 (
            .O(N__31925),
            .I(\c0.delay_counter_5 ));
    CascadeMux I__6373 (
            .O(N__31920),
            .I(N__31917));
    InMux I__6372 (
            .O(N__31917),
            .I(N__31914));
    LocalMux I__6371 (
            .O(N__31914),
            .I(n26_adj_2466));
    InMux I__6370 (
            .O(N__31911),
            .I(N__31907));
    InMux I__6369 (
            .O(N__31910),
            .I(N__31904));
    LocalMux I__6368 (
            .O(N__31907),
            .I(N__31900));
    LocalMux I__6367 (
            .O(N__31904),
            .I(N__31897));
    InMux I__6366 (
            .O(N__31903),
            .I(N__31894));
    Span4Mux_v I__6365 (
            .O(N__31900),
            .I(N__31889));
    Span4Mux_h I__6364 (
            .O(N__31897),
            .I(N__31889));
    LocalMux I__6363 (
            .O(N__31894),
            .I(data_out_frame2_7_1));
    Odrv4 I__6362 (
            .O(N__31889),
            .I(data_out_frame2_7_1));
    InMux I__6361 (
            .O(N__31884),
            .I(\c0.n16634 ));
    InMux I__6360 (
            .O(N__31881),
            .I(\c0.n16635 ));
    InMux I__6359 (
            .O(N__31878),
            .I(\c0.n16636 ));
    InMux I__6358 (
            .O(N__31875),
            .I(\c0.n16637 ));
    InMux I__6357 (
            .O(N__31872),
            .I(\c0.n16638 ));
    InMux I__6356 (
            .O(N__31869),
            .I(\c0.n16639 ));
    InMux I__6355 (
            .O(N__31866),
            .I(N__31863));
    LocalMux I__6354 (
            .O(N__31863),
            .I(N__31860));
    Odrv4 I__6353 (
            .O(N__31860),
            .I(\c0.n17727 ));
    InMux I__6352 (
            .O(N__31857),
            .I(N__31849));
    InMux I__6351 (
            .O(N__31856),
            .I(N__31849));
    InMux I__6350 (
            .O(N__31855),
            .I(N__31846));
    InMux I__6349 (
            .O(N__31854),
            .I(N__31843));
    LocalMux I__6348 (
            .O(N__31849),
            .I(N__31840));
    LocalMux I__6347 (
            .O(N__31846),
            .I(data_out_frame2_5_1));
    LocalMux I__6346 (
            .O(N__31843),
            .I(data_out_frame2_5_1));
    Odrv4 I__6345 (
            .O(N__31840),
            .I(data_out_frame2_5_1));
    InMux I__6344 (
            .O(N__31833),
            .I(N__31830));
    LocalMux I__6343 (
            .O(N__31830),
            .I(\c0.n18837 ));
    InMux I__6342 (
            .O(N__31827),
            .I(N__31824));
    LocalMux I__6341 (
            .O(N__31824),
            .I(N__31820));
    InMux I__6340 (
            .O(N__31823),
            .I(N__31817));
    Span4Mux_s0_v I__6339 (
            .O(N__31820),
            .I(N__31814));
    LocalMux I__6338 (
            .O(N__31817),
            .I(data_out_frame2_18_1));
    Odrv4 I__6337 (
            .O(N__31814),
            .I(data_out_frame2_18_1));
    InMux I__6336 (
            .O(N__31809),
            .I(N__31806));
    LocalMux I__6335 (
            .O(N__31806),
            .I(N__31802));
    InMux I__6334 (
            .O(N__31805),
            .I(N__31799));
    Span4Mux_h I__6333 (
            .O(N__31802),
            .I(N__31796));
    LocalMux I__6332 (
            .O(N__31799),
            .I(data_out_frame2_17_7));
    Odrv4 I__6331 (
            .O(N__31796),
            .I(data_out_frame2_17_7));
    CascadeMux I__6330 (
            .O(N__31791),
            .I(\c0.n10867_cascade_ ));
    CascadeMux I__6329 (
            .O(N__31788),
            .I(\c0.n17739_cascade_ ));
    CascadeMux I__6328 (
            .O(N__31785),
            .I(N__31781));
    InMux I__6327 (
            .O(N__31784),
            .I(N__31776));
    InMux I__6326 (
            .O(N__31781),
            .I(N__31776));
    LocalMux I__6325 (
            .O(N__31776),
            .I(data_out_frame2_17_0));
    InMux I__6324 (
            .O(N__31773),
            .I(N__31770));
    LocalMux I__6323 (
            .O(N__31770),
            .I(\c0.n18840 ));
    InMux I__6322 (
            .O(N__31767),
            .I(N__31764));
    LocalMux I__6321 (
            .O(N__31764),
            .I(\c0.n18795 ));
    InMux I__6320 (
            .O(N__31761),
            .I(N__31758));
    LocalMux I__6319 (
            .O(N__31758),
            .I(N__31754));
    InMux I__6318 (
            .O(N__31757),
            .I(N__31751));
    Span4Mux_h I__6317 (
            .O(N__31754),
            .I(N__31748));
    LocalMux I__6316 (
            .O(N__31751),
            .I(data_out_frame2_18_7));
    Odrv4 I__6315 (
            .O(N__31748),
            .I(data_out_frame2_18_7));
    InMux I__6314 (
            .O(N__31743),
            .I(N__31740));
    LocalMux I__6313 (
            .O(N__31740),
            .I(N__31737));
    Span4Mux_h I__6312 (
            .O(N__31737),
            .I(N__31734));
    Odrv4 I__6311 (
            .O(N__31734),
            .I(\c0.n18360 ));
    CascadeMux I__6310 (
            .O(N__31731),
            .I(N__31728));
    InMux I__6309 (
            .O(N__31728),
            .I(N__31725));
    LocalMux I__6308 (
            .O(N__31725),
            .I(N__31722));
    Odrv4 I__6307 (
            .O(N__31722),
            .I(\c0.n18256 ));
    CascadeMux I__6306 (
            .O(N__31719),
            .I(\c0.n14_adj_2359_cascade_ ));
    InMux I__6305 (
            .O(N__31716),
            .I(N__31713));
    LocalMux I__6304 (
            .O(N__31713),
            .I(\c0.data_out_frame2_20_0 ));
    InMux I__6303 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__6302 (
            .O(N__31707),
            .I(\c0.n15_adj_2429 ));
    InMux I__6301 (
            .O(N__31704),
            .I(N__31701));
    LocalMux I__6300 (
            .O(N__31701),
            .I(\c0.n17847 ));
    InMux I__6299 (
            .O(N__31698),
            .I(N__31694));
    InMux I__6298 (
            .O(N__31697),
            .I(N__31691));
    LocalMux I__6297 (
            .O(N__31694),
            .I(N__31688));
    LocalMux I__6296 (
            .O(N__31691),
            .I(data_out_2_5));
    Odrv4 I__6295 (
            .O(N__31688),
            .I(data_out_2_5));
    InMux I__6294 (
            .O(N__31683),
            .I(N__31680));
    LocalMux I__6293 (
            .O(N__31680),
            .I(N__31677));
    Odrv4 I__6292 (
            .O(N__31677),
            .I(\c0.n18335 ));
    InMux I__6291 (
            .O(N__31674),
            .I(N__31670));
    InMux I__6290 (
            .O(N__31673),
            .I(N__31667));
    LocalMux I__6289 (
            .O(N__31670),
            .I(\c0.data_out_2_3 ));
    LocalMux I__6288 (
            .O(N__31667),
            .I(\c0.data_out_2_3 ));
    CascadeMux I__6287 (
            .O(N__31662),
            .I(\c0.n19_cascade_ ));
    CascadeMux I__6286 (
            .O(N__31659),
            .I(N__31656));
    InMux I__6285 (
            .O(N__31656),
            .I(N__31653));
    LocalMux I__6284 (
            .O(N__31653),
            .I(\c0.data_out_frame2_19_1 ));
    InMux I__6283 (
            .O(N__31650),
            .I(N__31647));
    LocalMux I__6282 (
            .O(N__31647),
            .I(\c0.n20 ));
    InMux I__6281 (
            .O(N__31644),
            .I(N__31641));
    LocalMux I__6280 (
            .O(N__31641),
            .I(N__31638));
    Odrv4 I__6279 (
            .O(N__31638),
            .I(\c0.n18266 ));
    CascadeMux I__6278 (
            .O(N__31635),
            .I(n10_adj_2528_cascade_));
    InMux I__6277 (
            .O(N__31632),
            .I(N__31629));
    LocalMux I__6276 (
            .O(N__31629),
            .I(N__31625));
    InMux I__6275 (
            .O(N__31628),
            .I(N__31622));
    Span4Mux_h I__6274 (
            .O(N__31625),
            .I(N__31619));
    LocalMux I__6273 (
            .O(N__31622),
            .I(r_Tx_Data_2));
    Odrv4 I__6272 (
            .O(N__31619),
            .I(r_Tx_Data_2));
    CascadeMux I__6271 (
            .O(N__31614),
            .I(N__31611));
    InMux I__6270 (
            .O(N__31611),
            .I(N__31607));
    InMux I__6269 (
            .O(N__31610),
            .I(N__31604));
    LocalMux I__6268 (
            .O(N__31607),
            .I(data_out_3_5));
    LocalMux I__6267 (
            .O(N__31604),
            .I(data_out_3_5));
    InMux I__6266 (
            .O(N__31599),
            .I(N__31595));
    InMux I__6265 (
            .O(N__31598),
            .I(N__31592));
    LocalMux I__6264 (
            .O(N__31595),
            .I(data_out_1_6));
    LocalMux I__6263 (
            .O(N__31592),
            .I(data_out_1_6));
    InMux I__6262 (
            .O(N__31587),
            .I(N__31581));
    InMux I__6261 (
            .O(N__31586),
            .I(N__31581));
    LocalMux I__6260 (
            .O(N__31581),
            .I(\c0.data_out_0_6 ));
    CascadeMux I__6259 (
            .O(N__31578),
            .I(N__31575));
    InMux I__6258 (
            .O(N__31575),
            .I(N__31572));
    LocalMux I__6257 (
            .O(N__31572),
            .I(N__31569));
    Span4Mux_v I__6256 (
            .O(N__31569),
            .I(N__31566));
    Odrv4 I__6255 (
            .O(N__31566),
            .I(\c0.n1_adj_2272 ));
    CascadeMux I__6254 (
            .O(N__31563),
            .I(N__31560));
    InMux I__6253 (
            .O(N__31560),
            .I(N__31557));
    LocalMux I__6252 (
            .O(N__31557),
            .I(\c0.n5_adj_2241 ));
    InMux I__6251 (
            .O(N__31554),
            .I(N__31551));
    LocalMux I__6250 (
            .O(N__31551),
            .I(\c0.n18753 ));
    InMux I__6249 (
            .O(N__31548),
            .I(N__31545));
    LocalMux I__6248 (
            .O(N__31545),
            .I(N__31542));
    Odrv4 I__6247 (
            .O(N__31542),
            .I(\c0.n2 ));
    CascadeMux I__6246 (
            .O(N__31539),
            .I(N__31536));
    InMux I__6245 (
            .O(N__31536),
            .I(N__31533));
    LocalMux I__6244 (
            .O(N__31533),
            .I(N__31530));
    Span4Mux_h I__6243 (
            .O(N__31530),
            .I(N__31527));
    Odrv4 I__6242 (
            .O(N__31527),
            .I(\c0.n18189 ));
    CascadeMux I__6241 (
            .O(N__31524),
            .I(n18876_cascade_));
    InMux I__6240 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__6239 (
            .O(N__31518),
            .I(n10_adj_2531));
    CascadeMux I__6238 (
            .O(N__31515),
            .I(\c0.n5_adj_2196_cascade_ ));
    InMux I__6237 (
            .O(N__31512),
            .I(N__31509));
    LocalMux I__6236 (
            .O(N__31509),
            .I(\c0.n18873 ));
    CascadeMux I__6235 (
            .O(N__31506),
            .I(n5_cascade_));
    CascadeMux I__6234 (
            .O(N__31503),
            .I(N__31500));
    InMux I__6233 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__6232 (
            .O(N__31497),
            .I(\c0.n8_adj_2209 ));
    InMux I__6231 (
            .O(N__31494),
            .I(N__31491));
    LocalMux I__6230 (
            .O(N__31491),
            .I(n10_adj_2533));
    InMux I__6229 (
            .O(N__31488),
            .I(N__31482));
    InMux I__6228 (
            .O(N__31487),
            .I(N__31479));
    InMux I__6227 (
            .O(N__31486),
            .I(N__31474));
    InMux I__6226 (
            .O(N__31485),
            .I(N__31474));
    LocalMux I__6225 (
            .O(N__31482),
            .I(r_Bit_Index_1));
    LocalMux I__6224 (
            .O(N__31479),
            .I(r_Bit_Index_1));
    LocalMux I__6223 (
            .O(N__31474),
            .I(r_Bit_Index_1));
    InMux I__6222 (
            .O(N__31467),
            .I(N__31464));
    LocalMux I__6221 (
            .O(N__31464),
            .I(\c0.tx.n18167 ));
    CascadeMux I__6220 (
            .O(N__31461),
            .I(N__31456));
    CascadeMux I__6219 (
            .O(N__31460),
            .I(N__31452));
    InMux I__6218 (
            .O(N__31459),
            .I(N__31449));
    InMux I__6217 (
            .O(N__31456),
            .I(N__31446));
    InMux I__6216 (
            .O(N__31455),
            .I(N__31441));
    InMux I__6215 (
            .O(N__31452),
            .I(N__31441));
    LocalMux I__6214 (
            .O(N__31449),
            .I(r_Bit_Index_2));
    LocalMux I__6213 (
            .O(N__31446),
            .I(r_Bit_Index_2));
    LocalMux I__6212 (
            .O(N__31441),
            .I(r_Bit_Index_2));
    InMux I__6211 (
            .O(N__31434),
            .I(N__31431));
    LocalMux I__6210 (
            .O(N__31431),
            .I(\c0.tx.n18711 ));
    InMux I__6209 (
            .O(N__31428),
            .I(N__31424));
    InMux I__6208 (
            .O(N__31427),
            .I(N__31421));
    LocalMux I__6207 (
            .O(N__31424),
            .I(N__31418));
    LocalMux I__6206 (
            .O(N__31421),
            .I(r_Tx_Data_1));
    Odrv4 I__6205 (
            .O(N__31418),
            .I(r_Tx_Data_1));
    InMux I__6204 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__6203 (
            .O(N__31410),
            .I(\c0.tx.n18040 ));
    InMux I__6202 (
            .O(N__31407),
            .I(N__31404));
    LocalMux I__6201 (
            .O(N__31404),
            .I(\c0.n8_adj_2205 ));
    InMux I__6200 (
            .O(N__31401),
            .I(N__31392));
    InMux I__6199 (
            .O(N__31400),
            .I(N__31387));
    InMux I__6198 (
            .O(N__31399),
            .I(N__31387));
    InMux I__6197 (
            .O(N__31398),
            .I(N__31384));
    InMux I__6196 (
            .O(N__31397),
            .I(N__31381));
    InMux I__6195 (
            .O(N__31396),
            .I(N__31374));
    InMux I__6194 (
            .O(N__31395),
            .I(N__31374));
    LocalMux I__6193 (
            .O(N__31392),
            .I(N__31365));
    LocalMux I__6192 (
            .O(N__31387),
            .I(N__31365));
    LocalMux I__6191 (
            .O(N__31384),
            .I(N__31365));
    LocalMux I__6190 (
            .O(N__31381),
            .I(N__31365));
    InMux I__6189 (
            .O(N__31380),
            .I(N__31362));
    InMux I__6188 (
            .O(N__31379),
            .I(N__31359));
    LocalMux I__6187 (
            .O(N__31374),
            .I(\c0.tx.r_SM_Main_2 ));
    Odrv4 I__6186 (
            .O(N__31365),
            .I(\c0.tx.r_SM_Main_2 ));
    LocalMux I__6185 (
            .O(N__31362),
            .I(\c0.tx.r_SM_Main_2 ));
    LocalMux I__6184 (
            .O(N__31359),
            .I(\c0.tx.r_SM_Main_2 ));
    InMux I__6183 (
            .O(N__31350),
            .I(N__31337));
    InMux I__6182 (
            .O(N__31349),
            .I(N__31337));
    InMux I__6181 (
            .O(N__31348),
            .I(N__31337));
    InMux I__6180 (
            .O(N__31347),
            .I(N__31334));
    InMux I__6179 (
            .O(N__31346),
            .I(N__31331));
    CascadeMux I__6178 (
            .O(N__31345),
            .I(N__31328));
    InMux I__6177 (
            .O(N__31344),
            .I(N__31322));
    LocalMux I__6176 (
            .O(N__31337),
            .I(N__31315));
    LocalMux I__6175 (
            .O(N__31334),
            .I(N__31315));
    LocalMux I__6174 (
            .O(N__31331),
            .I(N__31315));
    InMux I__6173 (
            .O(N__31328),
            .I(N__31308));
    InMux I__6172 (
            .O(N__31327),
            .I(N__31308));
    InMux I__6171 (
            .O(N__31326),
            .I(N__31308));
    InMux I__6170 (
            .O(N__31325),
            .I(N__31305));
    LocalMux I__6169 (
            .O(N__31322),
            .I(\c0.tx.r_SM_Main_0 ));
    Odrv4 I__6168 (
            .O(N__31315),
            .I(\c0.tx.r_SM_Main_0 ));
    LocalMux I__6167 (
            .O(N__31308),
            .I(\c0.tx.r_SM_Main_0 ));
    LocalMux I__6166 (
            .O(N__31305),
            .I(\c0.tx.r_SM_Main_0 ));
    CascadeMux I__6165 (
            .O(N__31296),
            .I(N__31286));
    CascadeMux I__6164 (
            .O(N__31295),
            .I(N__31282));
    CascadeMux I__6163 (
            .O(N__31294),
            .I(N__31279));
    CascadeMux I__6162 (
            .O(N__31293),
            .I(N__31276));
    InMux I__6161 (
            .O(N__31292),
            .I(N__31272));
    InMux I__6160 (
            .O(N__31291),
            .I(N__31269));
    CascadeMux I__6159 (
            .O(N__31290),
            .I(N__31266));
    InMux I__6158 (
            .O(N__31289),
            .I(N__31261));
    InMux I__6157 (
            .O(N__31286),
            .I(N__31261));
    InMux I__6156 (
            .O(N__31285),
            .I(N__31258));
    InMux I__6155 (
            .O(N__31282),
            .I(N__31253));
    InMux I__6154 (
            .O(N__31279),
            .I(N__31253));
    InMux I__6153 (
            .O(N__31276),
            .I(N__31247));
    InMux I__6152 (
            .O(N__31275),
            .I(N__31247));
    LocalMux I__6151 (
            .O(N__31272),
            .I(N__31242));
    LocalMux I__6150 (
            .O(N__31269),
            .I(N__31242));
    InMux I__6149 (
            .O(N__31266),
            .I(N__31239));
    LocalMux I__6148 (
            .O(N__31261),
            .I(N__31232));
    LocalMux I__6147 (
            .O(N__31258),
            .I(N__31232));
    LocalMux I__6146 (
            .O(N__31253),
            .I(N__31232));
    InMux I__6145 (
            .O(N__31252),
            .I(N__31229));
    LocalMux I__6144 (
            .O(N__31247),
            .I(\c0.tx.r_SM_Main_1 ));
    Odrv4 I__6143 (
            .O(N__31242),
            .I(\c0.tx.r_SM_Main_1 ));
    LocalMux I__6142 (
            .O(N__31239),
            .I(\c0.tx.r_SM_Main_1 ));
    Odrv4 I__6141 (
            .O(N__31232),
            .I(\c0.tx.r_SM_Main_1 ));
    LocalMux I__6140 (
            .O(N__31229),
            .I(\c0.tx.r_SM_Main_1 ));
    InMux I__6139 (
            .O(N__31218),
            .I(N__31208));
    InMux I__6138 (
            .O(N__31217),
            .I(N__31208));
    InMux I__6137 (
            .O(N__31216),
            .I(N__31202));
    InMux I__6136 (
            .O(N__31215),
            .I(N__31202));
    InMux I__6135 (
            .O(N__31214),
            .I(N__31197));
    InMux I__6134 (
            .O(N__31213),
            .I(N__31197));
    LocalMux I__6133 (
            .O(N__31208),
            .I(N__31194));
    InMux I__6132 (
            .O(N__31207),
            .I(N__31191));
    LocalMux I__6131 (
            .O(N__31202),
            .I(N__31188));
    LocalMux I__6130 (
            .O(N__31197),
            .I(N__31181));
    Span4Mux_v I__6129 (
            .O(N__31194),
            .I(N__31181));
    LocalMux I__6128 (
            .O(N__31191),
            .I(N__31181));
    Span4Mux_v I__6127 (
            .O(N__31188),
            .I(N__31178));
    Span4Mux_h I__6126 (
            .O(N__31181),
            .I(N__31175));
    Odrv4 I__6125 (
            .O(N__31178),
            .I(\c0.tx.r_SM_Main_2_N_2031_1 ));
    Odrv4 I__6124 (
            .O(N__31175),
            .I(\c0.tx.r_SM_Main_2_N_2031_1 ));
    InMux I__6123 (
            .O(N__31170),
            .I(N__31161));
    InMux I__6122 (
            .O(N__31169),
            .I(N__31161));
    InMux I__6121 (
            .O(N__31168),
            .I(N__31161));
    LocalMux I__6120 (
            .O(N__31161),
            .I(N__31158));
    Odrv4 I__6119 (
            .O(N__31158),
            .I(n18012));
    InMux I__6118 (
            .O(N__31155),
            .I(N__31145));
    InMux I__6117 (
            .O(N__31154),
            .I(N__31142));
    InMux I__6116 (
            .O(N__31153),
            .I(N__31137));
    InMux I__6115 (
            .O(N__31152),
            .I(N__31137));
    InMux I__6114 (
            .O(N__31151),
            .I(N__31134));
    InMux I__6113 (
            .O(N__31150),
            .I(N__31129));
    InMux I__6112 (
            .O(N__31149),
            .I(N__31129));
    InMux I__6111 (
            .O(N__31148),
            .I(N__31126));
    LocalMux I__6110 (
            .O(N__31145),
            .I(N__31121));
    LocalMux I__6109 (
            .O(N__31142),
            .I(N__31121));
    LocalMux I__6108 (
            .O(N__31137),
            .I(r_Bit_Index_0));
    LocalMux I__6107 (
            .O(N__31134),
            .I(r_Bit_Index_0));
    LocalMux I__6106 (
            .O(N__31129),
            .I(r_Bit_Index_0));
    LocalMux I__6105 (
            .O(N__31126),
            .I(r_Bit_Index_0));
    Odrv4 I__6104 (
            .O(N__31121),
            .I(r_Bit_Index_0));
    InMux I__6103 (
            .O(N__31110),
            .I(N__31104));
    InMux I__6102 (
            .O(N__31109),
            .I(N__31104));
    LocalMux I__6101 (
            .O(N__31104),
            .I(r_Tx_Data_5));
    InMux I__6100 (
            .O(N__31101),
            .I(N__31098));
    LocalMux I__6099 (
            .O(N__31098),
            .I(\c0.tx.n18166 ));
    CascadeMux I__6098 (
            .O(N__31095),
            .I(n5440_cascade_));
    InMux I__6097 (
            .O(N__31092),
            .I(N__31089));
    LocalMux I__6096 (
            .O(N__31089),
            .I(n18016));
    CascadeMux I__6095 (
            .O(N__31086),
            .I(n18016_cascade_));
    CascadeMux I__6094 (
            .O(N__31083),
            .I(N__31080));
    InMux I__6093 (
            .O(N__31080),
            .I(N__31077));
    LocalMux I__6092 (
            .O(N__31077),
            .I(\c0.n8_adj_2207 ));
    InMux I__6091 (
            .O(N__31074),
            .I(N__31070));
    InMux I__6090 (
            .O(N__31073),
            .I(N__31067));
    LocalMux I__6089 (
            .O(N__31070),
            .I(\c0.tx.n13802 ));
    LocalMux I__6088 (
            .O(N__31067),
            .I(\c0.tx.n13802 ));
    CascadeMux I__6087 (
            .O(N__31062),
            .I(\c0.tx.n13802_cascade_ ));
    CascadeMux I__6086 (
            .O(N__31059),
            .I(\c0.tx.n6796_cascade_ ));
    CascadeMux I__6085 (
            .O(N__31056),
            .I(\c0.n4_cascade_ ));
    CascadeMux I__6084 (
            .O(N__31053),
            .I(n5341_cascade_));
    InMux I__6083 (
            .O(N__31050),
            .I(N__31047));
    LocalMux I__6082 (
            .O(N__31047),
            .I(N__31043));
    InMux I__6081 (
            .O(N__31046),
            .I(N__31040));
    Odrv4 I__6080 (
            .O(N__31043),
            .I(tx_transmit_N_1947_7));
    LocalMux I__6079 (
            .O(N__31040),
            .I(tx_transmit_N_1947_7));
    InMux I__6078 (
            .O(N__31035),
            .I(N__31031));
    InMux I__6077 (
            .O(N__31034),
            .I(N__31028));
    LocalMux I__6076 (
            .O(N__31031),
            .I(N__31025));
    LocalMux I__6075 (
            .O(N__31028),
            .I(byte_transmit_counter_7));
    Odrv4 I__6074 (
            .O(N__31025),
            .I(byte_transmit_counter_7));
    InMux I__6073 (
            .O(N__31020),
            .I(N__31017));
    LocalMux I__6072 (
            .O(N__31017),
            .I(N__31013));
    InMux I__6071 (
            .O(N__31016),
            .I(N__31010));
    Odrv4 I__6070 (
            .O(N__31013),
            .I(\c0.tx_transmit_N_1947_5 ));
    LocalMux I__6069 (
            .O(N__31010),
            .I(\c0.tx_transmit_N_1947_5 ));
    CascadeMux I__6068 (
            .O(N__31005),
            .I(N__30997));
    CascadeMux I__6067 (
            .O(N__31004),
            .I(N__30994));
    CascadeMux I__6066 (
            .O(N__31003),
            .I(N__30990));
    CascadeMux I__6065 (
            .O(N__31002),
            .I(N__30986));
    CascadeMux I__6064 (
            .O(N__31001),
            .I(N__30983));
    InMux I__6063 (
            .O(N__31000),
            .I(N__30979));
    InMux I__6062 (
            .O(N__30997),
            .I(N__30968));
    InMux I__6061 (
            .O(N__30994),
            .I(N__30968));
    InMux I__6060 (
            .O(N__30993),
            .I(N__30968));
    InMux I__6059 (
            .O(N__30990),
            .I(N__30968));
    InMux I__6058 (
            .O(N__30989),
            .I(N__30968));
    InMux I__6057 (
            .O(N__30986),
            .I(N__30961));
    InMux I__6056 (
            .O(N__30983),
            .I(N__30961));
    InMux I__6055 (
            .O(N__30982),
            .I(N__30961));
    LocalMux I__6054 (
            .O(N__30979),
            .I(n10973));
    LocalMux I__6053 (
            .O(N__30968),
            .I(n10973));
    LocalMux I__6052 (
            .O(N__30961),
            .I(n10973));
    InMux I__6051 (
            .O(N__30954),
            .I(N__30943));
    InMux I__6050 (
            .O(N__30953),
            .I(N__30943));
    InMux I__6049 (
            .O(N__30952),
            .I(N__30932));
    InMux I__6048 (
            .O(N__30951),
            .I(N__30932));
    InMux I__6047 (
            .O(N__30950),
            .I(N__30932));
    InMux I__6046 (
            .O(N__30949),
            .I(N__30932));
    InMux I__6045 (
            .O(N__30948),
            .I(N__30932));
    LocalMux I__6044 (
            .O(N__30943),
            .I(n5341));
    LocalMux I__6043 (
            .O(N__30932),
            .I(n5341));
    InMux I__6042 (
            .O(N__30927),
            .I(N__30923));
    InMux I__6041 (
            .O(N__30926),
            .I(N__30920));
    LocalMux I__6040 (
            .O(N__30923),
            .I(N__30917));
    LocalMux I__6039 (
            .O(N__30920),
            .I(\c0.byte_transmit_counter_5 ));
    Odrv4 I__6038 (
            .O(N__30917),
            .I(\c0.byte_transmit_counter_5 ));
    InMux I__6037 (
            .O(N__30912),
            .I(N__30909));
    LocalMux I__6036 (
            .O(N__30909),
            .I(\c0.n17998 ));
    InMux I__6035 (
            .O(N__30906),
            .I(N__30903));
    LocalMux I__6034 (
            .O(N__30903),
            .I(N__30900));
    Odrv4 I__6033 (
            .O(N__30900),
            .I(\c0.tx.n17938 ));
    CascadeMux I__6032 (
            .O(N__30897),
            .I(N__30894));
    InMux I__6031 (
            .O(N__30894),
            .I(N__30891));
    LocalMux I__6030 (
            .O(N__30891),
            .I(n10_adj_2536));
    InMux I__6029 (
            .O(N__30888),
            .I(N__30884));
    InMux I__6028 (
            .O(N__30887),
            .I(N__30881));
    LocalMux I__6027 (
            .O(N__30884),
            .I(byte_transmit_counter_6));
    LocalMux I__6026 (
            .O(N__30881),
            .I(byte_transmit_counter_6));
    InMux I__6025 (
            .O(N__30876),
            .I(N__30870));
    InMux I__6024 (
            .O(N__30875),
            .I(N__30870));
    LocalMux I__6023 (
            .O(N__30870),
            .I(tx_transmit_N_1947_6));
    CascadeMux I__6022 (
            .O(N__30867),
            .I(N__30863));
    InMux I__6021 (
            .O(N__30866),
            .I(N__30858));
    InMux I__6020 (
            .O(N__30863),
            .I(N__30858));
    LocalMux I__6019 (
            .O(N__30858),
            .I(tx_transmit_N_1947_4));
    InMux I__6018 (
            .O(N__30855),
            .I(N__30850));
    InMux I__6017 (
            .O(N__30854),
            .I(N__30847));
    InMux I__6016 (
            .O(N__30853),
            .I(N__30844));
    LocalMux I__6015 (
            .O(N__30850),
            .I(N__30841));
    LocalMux I__6014 (
            .O(N__30847),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__6013 (
            .O(N__30844),
            .I(\c0.tx2.r_Clock_Count_5 ));
    Odrv4 I__6012 (
            .O(N__30841),
            .I(\c0.tx2.r_Clock_Count_5 ));
    CascadeMux I__6011 (
            .O(N__30834),
            .I(\c0.tx2.n10_cascade_ ));
    CascadeMux I__6010 (
            .O(N__30831),
            .I(N__30826));
    InMux I__6009 (
            .O(N__30830),
            .I(N__30823));
    InMux I__6008 (
            .O(N__30829),
            .I(N__30820));
    InMux I__6007 (
            .O(N__30826),
            .I(N__30817));
    LocalMux I__6006 (
            .O(N__30823),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__6005 (
            .O(N__30820),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__6004 (
            .O(N__30817),
            .I(\c0.tx2.r_Clock_Count_3 ));
    InMux I__6003 (
            .O(N__30810),
            .I(N__30807));
    LocalMux I__6002 (
            .O(N__30807),
            .I(N__30804));
    Sp12to4 I__6001 (
            .O(N__30804),
            .I(N__30801));
    Odrv12 I__6000 (
            .O(N__30801),
            .I(\c0.tx2.n12775 ));
    InMux I__5999 (
            .O(N__30798),
            .I(N__30795));
    LocalMux I__5998 (
            .O(N__30795),
            .I(N__30792));
    Odrv12 I__5997 (
            .O(N__30792),
            .I(\c0.tx2.r_Tx_Data_1 ));
    InMux I__5996 (
            .O(N__30789),
            .I(N__30786));
    LocalMux I__5995 (
            .O(N__30786),
            .I(\c0.tx2.n18061 ));
    InMux I__5994 (
            .O(N__30783),
            .I(N__30778));
    InMux I__5993 (
            .O(N__30782),
            .I(N__30775));
    InMux I__5992 (
            .O(N__30781),
            .I(N__30770));
    LocalMux I__5991 (
            .O(N__30778),
            .I(N__30766));
    LocalMux I__5990 (
            .O(N__30775),
            .I(N__30763));
    InMux I__5989 (
            .O(N__30774),
            .I(N__30758));
    InMux I__5988 (
            .O(N__30773),
            .I(N__30755));
    LocalMux I__5987 (
            .O(N__30770),
            .I(N__30752));
    InMux I__5986 (
            .O(N__30769),
            .I(N__30749));
    Span4Mux_h I__5985 (
            .O(N__30766),
            .I(N__30744));
    Span4Mux_v I__5984 (
            .O(N__30763),
            .I(N__30744));
    InMux I__5983 (
            .O(N__30762),
            .I(N__30739));
    InMux I__5982 (
            .O(N__30761),
            .I(N__30739));
    LocalMux I__5981 (
            .O(N__30758),
            .I(r_SM_Main_2));
    LocalMux I__5980 (
            .O(N__30755),
            .I(r_SM_Main_2));
    Odrv4 I__5979 (
            .O(N__30752),
            .I(r_SM_Main_2));
    LocalMux I__5978 (
            .O(N__30749),
            .I(r_SM_Main_2));
    Odrv4 I__5977 (
            .O(N__30744),
            .I(r_SM_Main_2));
    LocalMux I__5976 (
            .O(N__30739),
            .I(r_SM_Main_2));
    CEMux I__5975 (
            .O(N__30726),
            .I(N__30721));
    CEMux I__5974 (
            .O(N__30725),
            .I(N__30718));
    InMux I__5973 (
            .O(N__30724),
            .I(N__30715));
    LocalMux I__5972 (
            .O(N__30721),
            .I(N__30712));
    LocalMux I__5971 (
            .O(N__30718),
            .I(N__30709));
    LocalMux I__5970 (
            .O(N__30715),
            .I(N__30706));
    Odrv4 I__5969 (
            .O(N__30712),
            .I(n11096));
    Odrv4 I__5968 (
            .O(N__30709),
            .I(n11096));
    Odrv12 I__5967 (
            .O(N__30706),
            .I(n11096));
    CascadeMux I__5966 (
            .O(N__30699),
            .I(\c0.n18260_cascade_ ));
    InMux I__5965 (
            .O(N__30696),
            .I(N__30693));
    LocalMux I__5964 (
            .O(N__30693),
            .I(\c0.n130 ));
    InMux I__5963 (
            .O(N__30690),
            .I(N__30687));
    LocalMux I__5962 (
            .O(N__30687),
            .I(\c0.n3465 ));
    SRMux I__5961 (
            .O(N__30684),
            .I(N__30681));
    LocalMux I__5960 (
            .O(N__30681),
            .I(N__30678));
    Odrv4 I__5959 (
            .O(N__30678),
            .I(\c0.n4806 ));
    InMux I__5958 (
            .O(N__30675),
            .I(N__30672));
    LocalMux I__5957 (
            .O(N__30672),
            .I(N__30669));
    Span4Mux_h I__5956 (
            .O(N__30669),
            .I(N__30666));
    Odrv4 I__5955 (
            .O(N__30666),
            .I(\c0.n18362 ));
    CascadeMux I__5954 (
            .O(N__30663),
            .I(N__30660));
    InMux I__5953 (
            .O(N__30660),
            .I(N__30654));
    CascadeMux I__5952 (
            .O(N__30659),
            .I(N__30651));
    CascadeMux I__5951 (
            .O(N__30658),
            .I(N__30647));
    CascadeMux I__5950 (
            .O(N__30657),
            .I(N__30644));
    LocalMux I__5949 (
            .O(N__30654),
            .I(N__30639));
    InMux I__5948 (
            .O(N__30651),
            .I(N__30636));
    CascadeMux I__5947 (
            .O(N__30650),
            .I(N__30633));
    InMux I__5946 (
            .O(N__30647),
            .I(N__30630));
    InMux I__5945 (
            .O(N__30644),
            .I(N__30627));
    CascadeMux I__5944 (
            .O(N__30643),
            .I(N__30624));
    CascadeMux I__5943 (
            .O(N__30642),
            .I(N__30621));
    Span4Mux_v I__5942 (
            .O(N__30639),
            .I(N__30618));
    LocalMux I__5941 (
            .O(N__30636),
            .I(N__30615));
    InMux I__5940 (
            .O(N__30633),
            .I(N__30612));
    LocalMux I__5939 (
            .O(N__30630),
            .I(N__30607));
    LocalMux I__5938 (
            .O(N__30627),
            .I(N__30607));
    InMux I__5937 (
            .O(N__30624),
            .I(N__30604));
    InMux I__5936 (
            .O(N__30621),
            .I(N__30601));
    Span4Mux_h I__5935 (
            .O(N__30618),
            .I(N__30592));
    Span4Mux_s0_v I__5934 (
            .O(N__30615),
            .I(N__30592));
    LocalMux I__5933 (
            .O(N__30612),
            .I(N__30592));
    Span4Mux_s2_v I__5932 (
            .O(N__30607),
            .I(N__30587));
    LocalMux I__5931 (
            .O(N__30604),
            .I(N__30587));
    LocalMux I__5930 (
            .O(N__30601),
            .I(N__30584));
    CascadeMux I__5929 (
            .O(N__30600),
            .I(N__30581));
    CascadeMux I__5928 (
            .O(N__30599),
            .I(N__30578));
    Span4Mux_v I__5927 (
            .O(N__30592),
            .I(N__30575));
    Span4Mux_h I__5926 (
            .O(N__30587),
            .I(N__30570));
    Span4Mux_v I__5925 (
            .O(N__30584),
            .I(N__30570));
    InMux I__5924 (
            .O(N__30581),
            .I(N__30567));
    InMux I__5923 (
            .O(N__30578),
            .I(N__30564));
    Odrv4 I__5922 (
            .O(N__30575),
            .I(\c0.n12359 ));
    Odrv4 I__5921 (
            .O(N__30570),
            .I(\c0.n12359 ));
    LocalMux I__5920 (
            .O(N__30567),
            .I(\c0.n12359 ));
    LocalMux I__5919 (
            .O(N__30564),
            .I(\c0.n12359 ));
    InMux I__5918 (
            .O(N__30555),
            .I(N__30548));
    InMux I__5917 (
            .O(N__30554),
            .I(N__30543));
    InMux I__5916 (
            .O(N__30553),
            .I(N__30540));
    InMux I__5915 (
            .O(N__30552),
            .I(N__30537));
    InMux I__5914 (
            .O(N__30551),
            .I(N__30534));
    LocalMux I__5913 (
            .O(N__30548),
            .I(N__30531));
    InMux I__5912 (
            .O(N__30547),
            .I(N__30528));
    InMux I__5911 (
            .O(N__30546),
            .I(N__30525));
    LocalMux I__5910 (
            .O(N__30543),
            .I(N__30520));
    LocalMux I__5909 (
            .O(N__30540),
            .I(N__30520));
    LocalMux I__5908 (
            .O(N__30537),
            .I(N__30512));
    LocalMux I__5907 (
            .O(N__30534),
            .I(N__30512));
    Span4Mux_s0_v I__5906 (
            .O(N__30531),
            .I(N__30505));
    LocalMux I__5905 (
            .O(N__30528),
            .I(N__30505));
    LocalMux I__5904 (
            .O(N__30525),
            .I(N__30505));
    Span4Mux_v I__5903 (
            .O(N__30520),
            .I(N__30502));
    InMux I__5902 (
            .O(N__30519),
            .I(N__30499));
    InMux I__5901 (
            .O(N__30518),
            .I(N__30496));
    InMux I__5900 (
            .O(N__30517),
            .I(N__30493));
    Span12Mux_s4_v I__5899 (
            .O(N__30512),
            .I(N__30489));
    Span4Mux_v I__5898 (
            .O(N__30505),
            .I(N__30484));
    Span4Mux_h I__5897 (
            .O(N__30502),
            .I(N__30484));
    LocalMux I__5896 (
            .O(N__30499),
            .I(N__30481));
    LocalMux I__5895 (
            .O(N__30496),
            .I(N__30478));
    LocalMux I__5894 (
            .O(N__30493),
            .I(N__30475));
    InMux I__5893 (
            .O(N__30492),
            .I(N__30472));
    Odrv12 I__5892 (
            .O(N__30489),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__5891 (
            .O(N__30484),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__5890 (
            .O(N__30481),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__5889 (
            .O(N__30478),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__5888 (
            .O(N__30475),
            .I(FRAME_MATCHER_i_31__N_1272));
    LocalMux I__5887 (
            .O(N__30472),
            .I(FRAME_MATCHER_i_31__N_1272));
    SRMux I__5886 (
            .O(N__30459),
            .I(N__30456));
    LocalMux I__5885 (
            .O(N__30456),
            .I(N__30453));
    Odrv12 I__5884 (
            .O(N__30453),
            .I(\c0.n4_adj_2204 ));
    InMux I__5883 (
            .O(N__30450),
            .I(N__30444));
    InMux I__5882 (
            .O(N__30449),
            .I(N__30444));
    LocalMux I__5881 (
            .O(N__30444),
            .I(\c0.tx2.n13800 ));
    CascadeMux I__5880 (
            .O(N__30441),
            .I(N__30431));
    InMux I__5879 (
            .O(N__30440),
            .I(N__30427));
    InMux I__5878 (
            .O(N__30439),
            .I(N__30424));
    InMux I__5877 (
            .O(N__30438),
            .I(N__30417));
    InMux I__5876 (
            .O(N__30437),
            .I(N__30417));
    InMux I__5875 (
            .O(N__30436),
            .I(N__30417));
    InMux I__5874 (
            .O(N__30435),
            .I(N__30407));
    InMux I__5873 (
            .O(N__30434),
            .I(N__30407));
    InMux I__5872 (
            .O(N__30431),
            .I(N__30407));
    InMux I__5871 (
            .O(N__30430),
            .I(N__30407));
    LocalMux I__5870 (
            .O(N__30427),
            .I(N__30404));
    LocalMux I__5869 (
            .O(N__30424),
            .I(N__30399));
    LocalMux I__5868 (
            .O(N__30417),
            .I(N__30399));
    CascadeMux I__5867 (
            .O(N__30416),
            .I(N__30396));
    LocalMux I__5866 (
            .O(N__30407),
            .I(N__30393));
    Span4Mux_v I__5865 (
            .O(N__30404),
            .I(N__30388));
    Span4Mux_v I__5864 (
            .O(N__30399),
            .I(N__30388));
    InMux I__5863 (
            .O(N__30396),
            .I(N__30385));
    Span4Mux_h I__5862 (
            .O(N__30393),
            .I(N__30382));
    Span4Mux_h I__5861 (
            .O(N__30388),
            .I(N__30379));
    LocalMux I__5860 (
            .O(N__30385),
            .I(r_SM_Main_1));
    Odrv4 I__5859 (
            .O(N__30382),
            .I(r_SM_Main_1));
    Odrv4 I__5858 (
            .O(N__30379),
            .I(r_SM_Main_1));
    InMux I__5857 (
            .O(N__30372),
            .I(N__30369));
    LocalMux I__5856 (
            .O(N__30369),
            .I(N__30363));
    InMux I__5855 (
            .O(N__30368),
            .I(N__30360));
    InMux I__5854 (
            .O(N__30367),
            .I(N__30357));
    CascadeMux I__5853 (
            .O(N__30366),
            .I(N__30352));
    Span4Mux_v I__5852 (
            .O(N__30363),
            .I(N__30349));
    LocalMux I__5851 (
            .O(N__30360),
            .I(N__30344));
    LocalMux I__5850 (
            .O(N__30357),
            .I(N__30344));
    InMux I__5849 (
            .O(N__30356),
            .I(N__30341));
    CascadeMux I__5848 (
            .O(N__30355),
            .I(N__30336));
    InMux I__5847 (
            .O(N__30352),
            .I(N__30333));
    Span4Mux_s2_v I__5846 (
            .O(N__30349),
            .I(N__30330));
    Span4Mux_v I__5845 (
            .O(N__30344),
            .I(N__30327));
    LocalMux I__5844 (
            .O(N__30341),
            .I(N__30324));
    InMux I__5843 (
            .O(N__30340),
            .I(N__30317));
    InMux I__5842 (
            .O(N__30339),
            .I(N__30317));
    InMux I__5841 (
            .O(N__30336),
            .I(N__30317));
    LocalMux I__5840 (
            .O(N__30333),
            .I(r_SM_Main_0));
    Odrv4 I__5839 (
            .O(N__30330),
            .I(r_SM_Main_0));
    Odrv4 I__5838 (
            .O(N__30327),
            .I(r_SM_Main_0));
    Odrv4 I__5837 (
            .O(N__30324),
            .I(r_SM_Main_0));
    LocalMux I__5836 (
            .O(N__30317),
            .I(r_SM_Main_0));
    InMux I__5835 (
            .O(N__30306),
            .I(N__30303));
    LocalMux I__5834 (
            .O(N__30303),
            .I(N__30300));
    Span4Mux_h I__5833 (
            .O(N__30300),
            .I(N__30297));
    Odrv4 I__5832 (
            .O(N__30297),
            .I(n3));
    InMux I__5831 (
            .O(N__30294),
            .I(N__30291));
    LocalMux I__5830 (
            .O(N__30291),
            .I(N__30288));
    Span12Mux_s7_v I__5829 (
            .O(N__30288),
            .I(N__30285));
    Odrv12 I__5828 (
            .O(N__30285),
            .I(\c0.tx2.n18164 ));
    InMux I__5827 (
            .O(N__30282),
            .I(N__30279));
    LocalMux I__5826 (
            .O(N__30279),
            .I(N__30276));
    Span4Mux_v I__5825 (
            .O(N__30276),
            .I(N__30273));
    Span4Mux_h I__5824 (
            .O(N__30273),
            .I(N__30270));
    Odrv4 I__5823 (
            .O(N__30270),
            .I(\c0.tx2.n18163 ));
    InMux I__5822 (
            .O(N__30267),
            .I(N__30264));
    LocalMux I__5821 (
            .O(N__30264),
            .I(\c0.tx2.n18062 ));
    CascadeMux I__5820 (
            .O(N__30261),
            .I(\c0.tx2.n18717_cascade_ ));
    InMux I__5819 (
            .O(N__30258),
            .I(N__30255));
    LocalMux I__5818 (
            .O(N__30255),
            .I(\c0.tx2.o_Tx_Serial_N_2062 ));
    InMux I__5817 (
            .O(N__30252),
            .I(N__30248));
    InMux I__5816 (
            .O(N__30251),
            .I(N__30245));
    LocalMux I__5815 (
            .O(N__30248),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__5814 (
            .O(N__30245),
            .I(\c0.tx2.r_Clock_Count_4 ));
    InMux I__5813 (
            .O(N__30240),
            .I(N__30236));
    InMux I__5812 (
            .O(N__30239),
            .I(N__30233));
    LocalMux I__5811 (
            .O(N__30236),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__5810 (
            .O(N__30233),
            .I(\c0.tx2.r_Clock_Count_2 ));
    CascadeMux I__5809 (
            .O(N__30228),
            .I(N__30224));
    InMux I__5808 (
            .O(N__30227),
            .I(N__30221));
    InMux I__5807 (
            .O(N__30224),
            .I(N__30218));
    LocalMux I__5806 (
            .O(N__30221),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__5805 (
            .O(N__30218),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__5804 (
            .O(N__30213),
            .I(N__30209));
    InMux I__5803 (
            .O(N__30212),
            .I(N__30206));
    LocalMux I__5802 (
            .O(N__30209),
            .I(\c0.tx2.r_Clock_Count_0 ));
    LocalMux I__5801 (
            .O(N__30206),
            .I(\c0.tx2.r_Clock_Count_0 ));
    InMux I__5800 (
            .O(N__30201),
            .I(N__30198));
    LocalMux I__5799 (
            .O(N__30198),
            .I(N__30195));
    Odrv4 I__5798 (
            .O(N__30195),
            .I(\c0.tx2.n10 ));
    InMux I__5797 (
            .O(N__30192),
            .I(N__30188));
    InMux I__5796 (
            .O(N__30191),
            .I(N__30185));
    LocalMux I__5795 (
            .O(N__30188),
            .I(N__30181));
    LocalMux I__5794 (
            .O(N__30185),
            .I(N__30178));
    InMux I__5793 (
            .O(N__30184),
            .I(N__30175));
    Span4Mux_v I__5792 (
            .O(N__30181),
            .I(N__30172));
    Span4Mux_h I__5791 (
            .O(N__30178),
            .I(N__30169));
    LocalMux I__5790 (
            .O(N__30175),
            .I(tx2_active));
    Odrv4 I__5789 (
            .O(N__30172),
            .I(tx2_active));
    Odrv4 I__5788 (
            .O(N__30169),
            .I(tx2_active));
    InMux I__5787 (
            .O(N__30162),
            .I(N__30158));
    InMux I__5786 (
            .O(N__30161),
            .I(N__30155));
    LocalMux I__5785 (
            .O(N__30158),
            .I(N__30150));
    LocalMux I__5784 (
            .O(N__30155),
            .I(N__30150));
    Span4Mux_h I__5783 (
            .O(N__30150),
            .I(N__30146));
    InMux I__5782 (
            .O(N__30149),
            .I(N__30143));
    Odrv4 I__5781 (
            .O(N__30146),
            .I(\c0.n14064 ));
    LocalMux I__5780 (
            .O(N__30143),
            .I(\c0.n14064 ));
    CascadeMux I__5779 (
            .O(N__30138),
            .I(\c0.n12359_cascade_ ));
    CascadeMux I__5778 (
            .O(N__30135),
            .I(\c0.n6_adj_2443_cascade_ ));
    InMux I__5777 (
            .O(N__30132),
            .I(N__30128));
    SRMux I__5776 (
            .O(N__30131),
            .I(N__30125));
    LocalMux I__5775 (
            .O(N__30128),
            .I(N__30121));
    LocalMux I__5774 (
            .O(N__30125),
            .I(N__30118));
    InMux I__5773 (
            .O(N__30124),
            .I(N__30115));
    Span4Mux_v I__5772 (
            .O(N__30121),
            .I(N__30105));
    Sp12to4 I__5771 (
            .O(N__30118),
            .I(N__30100));
    LocalMux I__5770 (
            .O(N__30115),
            .I(N__30100));
    InMux I__5769 (
            .O(N__30114),
            .I(N__30097));
    InMux I__5768 (
            .O(N__30113),
            .I(N__30090));
    InMux I__5767 (
            .O(N__30112),
            .I(N__30090));
    InMux I__5766 (
            .O(N__30111),
            .I(N__30090));
    InMux I__5765 (
            .O(N__30110),
            .I(N__30083));
    InMux I__5764 (
            .O(N__30109),
            .I(N__30083));
    InMux I__5763 (
            .O(N__30108),
            .I(N__30083));
    Odrv4 I__5762 (
            .O(N__30105),
            .I(\c0.n10513 ));
    Odrv12 I__5761 (
            .O(N__30100),
            .I(\c0.n10513 ));
    LocalMux I__5760 (
            .O(N__30097),
            .I(\c0.n10513 ));
    LocalMux I__5759 (
            .O(N__30090),
            .I(\c0.n10513 ));
    LocalMux I__5758 (
            .O(N__30083),
            .I(\c0.n10513 ));
    InMux I__5757 (
            .O(N__30072),
            .I(N__30061));
    InMux I__5756 (
            .O(N__30071),
            .I(N__30061));
    InMux I__5755 (
            .O(N__30070),
            .I(N__30058));
    InMux I__5754 (
            .O(N__30069),
            .I(N__30051));
    InMux I__5753 (
            .O(N__30068),
            .I(N__30051));
    InMux I__5752 (
            .O(N__30067),
            .I(N__30051));
    CascadeMux I__5751 (
            .O(N__30066),
            .I(N__30046));
    LocalMux I__5750 (
            .O(N__30061),
            .I(N__30036));
    LocalMux I__5749 (
            .O(N__30058),
            .I(N__30036));
    LocalMux I__5748 (
            .O(N__30051),
            .I(N__30036));
    InMux I__5747 (
            .O(N__30050),
            .I(N__30031));
    InMux I__5746 (
            .O(N__30049),
            .I(N__30026));
    InMux I__5745 (
            .O(N__30046),
            .I(N__30026));
    InMux I__5744 (
            .O(N__30045),
            .I(N__30023));
    CascadeMux I__5743 (
            .O(N__30044),
            .I(N__30018));
    CascadeMux I__5742 (
            .O(N__30043),
            .I(N__30015));
    Span4Mux_h I__5741 (
            .O(N__30036),
            .I(N__30012));
    CascadeMux I__5740 (
            .O(N__30035),
            .I(N__30008));
    InMux I__5739 (
            .O(N__30034),
            .I(N__30004));
    LocalMux I__5738 (
            .O(N__30031),
            .I(N__29997));
    LocalMux I__5737 (
            .O(N__30026),
            .I(N__29997));
    LocalMux I__5736 (
            .O(N__30023),
            .I(N__29997));
    InMux I__5735 (
            .O(N__30022),
            .I(N__29990));
    InMux I__5734 (
            .O(N__30021),
            .I(N__29990));
    InMux I__5733 (
            .O(N__30018),
            .I(N__29990));
    InMux I__5732 (
            .O(N__30015),
            .I(N__29987));
    Span4Mux_v I__5731 (
            .O(N__30012),
            .I(N__29984));
    InMux I__5730 (
            .O(N__30011),
            .I(N__29979));
    InMux I__5729 (
            .O(N__30008),
            .I(N__29974));
    InMux I__5728 (
            .O(N__30007),
            .I(N__29974));
    LocalMux I__5727 (
            .O(N__30004),
            .I(N__29967));
    Span4Mux_h I__5726 (
            .O(N__29997),
            .I(N__29967));
    LocalMux I__5725 (
            .O(N__29990),
            .I(N__29967));
    LocalMux I__5724 (
            .O(N__29987),
            .I(N__29962));
    Span4Mux_h I__5723 (
            .O(N__29984),
            .I(N__29962));
    InMux I__5722 (
            .O(N__29983),
            .I(N__29957));
    InMux I__5721 (
            .O(N__29982),
            .I(N__29957));
    LocalMux I__5720 (
            .O(N__29979),
            .I(N__29950));
    LocalMux I__5719 (
            .O(N__29974),
            .I(N__29950));
    Span4Mux_h I__5718 (
            .O(N__29967),
            .I(N__29950));
    Odrv4 I__5717 (
            .O(N__29962),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__5716 (
            .O(N__29957),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__5715 (
            .O(N__29950),
            .I(\c0.FRAME_MATCHER_state_0 ));
    CascadeMux I__5714 (
            .O(N__29943),
            .I(N__29940));
    InMux I__5713 (
            .O(N__29940),
            .I(N__29937));
    LocalMux I__5712 (
            .O(N__29937),
            .I(N__29934));
    Span12Mux_v I__5711 (
            .O(N__29934),
            .I(N__29931));
    Odrv12 I__5710 (
            .O(N__29931),
            .I(\c0.n10958 ));
    InMux I__5709 (
            .O(N__29928),
            .I(N__29922));
    CascadeMux I__5708 (
            .O(N__29927),
            .I(N__29919));
    InMux I__5707 (
            .O(N__29926),
            .I(N__29913));
    InMux I__5706 (
            .O(N__29925),
            .I(N__29913));
    LocalMux I__5705 (
            .O(N__29922),
            .I(N__29910));
    InMux I__5704 (
            .O(N__29919),
            .I(N__29907));
    InMux I__5703 (
            .O(N__29918),
            .I(N__29904));
    LocalMux I__5702 (
            .O(N__29913),
            .I(N__29901));
    Span4Mux_h I__5701 (
            .O(N__29910),
            .I(N__29898));
    LocalMux I__5700 (
            .O(N__29907),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2213 ));
    LocalMux I__5699 (
            .O(N__29904),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2213 ));
    Odrv4 I__5698 (
            .O(N__29901),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2213 ));
    Odrv4 I__5697 (
            .O(N__29898),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2213 ));
    InMux I__5696 (
            .O(N__29889),
            .I(N__29886));
    LocalMux I__5695 (
            .O(N__29886),
            .I(N__29883));
    Span4Mux_s3_v I__5694 (
            .O(N__29883),
            .I(N__29880));
    Odrv4 I__5693 (
            .O(N__29880),
            .I(n6707));
    InMux I__5692 (
            .O(N__29877),
            .I(N__29873));
    InMux I__5691 (
            .O(N__29876),
            .I(N__29870));
    LocalMux I__5690 (
            .O(N__29873),
            .I(N__29867));
    LocalMux I__5689 (
            .O(N__29870),
            .I(N__29864));
    Span4Mux_v I__5688 (
            .O(N__29867),
            .I(N__29861));
    Span12Mux_s7_v I__5687 (
            .O(N__29864),
            .I(N__29858));
    Span4Mux_h I__5686 (
            .O(N__29861),
            .I(N__29855));
    Odrv12 I__5685 (
            .O(N__29858),
            .I(\c0.tx2.n12769 ));
    Odrv4 I__5684 (
            .O(N__29855),
            .I(\c0.tx2.n12769 ));
    InMux I__5683 (
            .O(N__29850),
            .I(N__29846));
    CascadeMux I__5682 (
            .O(N__29849),
            .I(N__29843));
    LocalMux I__5681 (
            .O(N__29846),
            .I(N__29838));
    InMux I__5680 (
            .O(N__29843),
            .I(N__29835));
    InMux I__5679 (
            .O(N__29842),
            .I(N__29832));
    InMux I__5678 (
            .O(N__29841),
            .I(N__29829));
    Span4Mux_v I__5677 (
            .O(N__29838),
            .I(N__29825));
    LocalMux I__5676 (
            .O(N__29835),
            .I(N__29818));
    LocalMux I__5675 (
            .O(N__29832),
            .I(N__29818));
    LocalMux I__5674 (
            .O(N__29829),
            .I(N__29818));
    InMux I__5673 (
            .O(N__29828),
            .I(N__29815));
    Odrv4 I__5672 (
            .O(N__29825),
            .I(r_SM_Main_2_N_2031_1));
    Odrv4 I__5671 (
            .O(N__29818),
            .I(r_SM_Main_2_N_2031_1));
    LocalMux I__5670 (
            .O(N__29815),
            .I(r_SM_Main_2_N_2031_1));
    CascadeMux I__5669 (
            .O(N__29808),
            .I(r_SM_Main_2_N_2031_1_cascade_));
    CascadeMux I__5668 (
            .O(N__29805),
            .I(n18014_cascade_));
    CascadeMux I__5667 (
            .O(N__29802),
            .I(\c0.n5_adj_2435_cascade_ ));
    CascadeMux I__5666 (
            .O(N__29799),
            .I(N__29796));
    InMux I__5665 (
            .O(N__29796),
            .I(N__29793));
    LocalMux I__5664 (
            .O(N__29793),
            .I(N__29790));
    Odrv4 I__5663 (
            .O(N__29790),
            .I(\c0.n6_adj_2223 ));
    CascadeMux I__5662 (
            .O(N__29787),
            .I(\c0.n18687_cascade_ ));
    CascadeMux I__5661 (
            .O(N__29784),
            .I(N__29781));
    InMux I__5660 (
            .O(N__29781),
            .I(N__29778));
    LocalMux I__5659 (
            .O(N__29778),
            .I(N__29775));
    Odrv4 I__5658 (
            .O(N__29775),
            .I(\c0.n18690 ));
    CascadeMux I__5657 (
            .O(N__29772),
            .I(N__29769));
    InMux I__5656 (
            .O(N__29769),
            .I(N__29766));
    LocalMux I__5655 (
            .O(N__29766),
            .I(N__29763));
    Span4Mux_v I__5654 (
            .O(N__29763),
            .I(N__29760));
    Span4Mux_h I__5653 (
            .O(N__29760),
            .I(N__29757));
    Odrv4 I__5652 (
            .O(N__29757),
            .I(\c0.n5_adj_2197 ));
    InMux I__5651 (
            .O(N__29754),
            .I(N__29751));
    LocalMux I__5650 (
            .O(N__29751),
            .I(N__29748));
    Span12Mux_s3_v I__5649 (
            .O(N__29748),
            .I(N__29745));
    Odrv12 I__5648 (
            .O(N__29745),
            .I(\c0.n6 ));
    InMux I__5647 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__5646 (
            .O(N__29739),
            .I(N__29736));
    Odrv4 I__5645 (
            .O(N__29736),
            .I(\c0.n6_adj_2354 ));
    InMux I__5644 (
            .O(N__29733),
            .I(N__29730));
    LocalMux I__5643 (
            .O(N__29730),
            .I(\c0.n18855 ));
    CascadeMux I__5642 (
            .O(N__29727),
            .I(\c0.n10893_cascade_ ));
    InMux I__5641 (
            .O(N__29724),
            .I(N__29720));
    InMux I__5640 (
            .O(N__29723),
            .I(N__29717));
    LocalMux I__5639 (
            .O(N__29720),
            .I(N__29714));
    LocalMux I__5638 (
            .O(N__29717),
            .I(data_out_frame2_17_1));
    Odrv4 I__5637 (
            .O(N__29714),
            .I(data_out_frame2_17_1));
    CascadeMux I__5636 (
            .O(N__29709),
            .I(\c0.n18888_cascade_ ));
    CascadeMux I__5635 (
            .O(N__29706),
            .I(\c0.n18789_cascade_ ));
    CascadeMux I__5634 (
            .O(N__29703),
            .I(\c0.n18792_cascade_ ));
    InMux I__5633 (
            .O(N__29700),
            .I(N__29697));
    LocalMux I__5632 (
            .O(N__29697),
            .I(\c0.n22_adj_2270 ));
    InMux I__5631 (
            .O(N__29694),
            .I(N__29691));
    LocalMux I__5630 (
            .O(N__29691),
            .I(\c0.n18885 ));
    CascadeMux I__5629 (
            .O(N__29688),
            .I(\c0.n10861_cascade_ ));
    CascadeMux I__5628 (
            .O(N__29685),
            .I(N__29682));
    InMux I__5627 (
            .O(N__29682),
            .I(N__29679));
    LocalMux I__5626 (
            .O(N__29679),
            .I(\c0.n18798 ));
    InMux I__5625 (
            .O(N__29676),
            .I(N__29672));
    InMux I__5624 (
            .O(N__29675),
            .I(N__29669));
    LocalMux I__5623 (
            .O(N__29672),
            .I(\control.pwm_delay_2 ));
    LocalMux I__5622 (
            .O(N__29669),
            .I(\control.pwm_delay_2 ));
    InMux I__5621 (
            .O(N__29664),
            .I(\control.n16648 ));
    CascadeMux I__5620 (
            .O(N__29661),
            .I(N__29657));
    InMux I__5619 (
            .O(N__29660),
            .I(N__29654));
    InMux I__5618 (
            .O(N__29657),
            .I(N__29651));
    LocalMux I__5617 (
            .O(N__29654),
            .I(\control.pwm_delay_3 ));
    LocalMux I__5616 (
            .O(N__29651),
            .I(\control.pwm_delay_3 ));
    InMux I__5615 (
            .O(N__29646),
            .I(\control.n16649 ));
    InMux I__5614 (
            .O(N__29643),
            .I(N__29639));
    InMux I__5613 (
            .O(N__29642),
            .I(N__29636));
    LocalMux I__5612 (
            .O(N__29639),
            .I(\control.pwm_delay_4 ));
    LocalMux I__5611 (
            .O(N__29636),
            .I(\control.pwm_delay_4 ));
    InMux I__5610 (
            .O(N__29631),
            .I(\control.n16650 ));
    InMux I__5609 (
            .O(N__29628),
            .I(N__29624));
    InMux I__5608 (
            .O(N__29627),
            .I(N__29621));
    LocalMux I__5607 (
            .O(N__29624),
            .I(\control.pwm_delay_5 ));
    LocalMux I__5606 (
            .O(N__29621),
            .I(\control.pwm_delay_5 ));
    InMux I__5605 (
            .O(N__29616),
            .I(\control.n16651 ));
    InMux I__5604 (
            .O(N__29613),
            .I(N__29609));
    InMux I__5603 (
            .O(N__29612),
            .I(N__29606));
    LocalMux I__5602 (
            .O(N__29609),
            .I(\control.pwm_delay_6 ));
    LocalMux I__5601 (
            .O(N__29606),
            .I(\control.pwm_delay_6 ));
    InMux I__5600 (
            .O(N__29601),
            .I(\control.n16652 ));
    InMux I__5599 (
            .O(N__29598),
            .I(N__29594));
    InMux I__5598 (
            .O(N__29597),
            .I(N__29591));
    LocalMux I__5597 (
            .O(N__29594),
            .I(\control.pwm_delay_7 ));
    LocalMux I__5596 (
            .O(N__29591),
            .I(\control.pwm_delay_7 ));
    InMux I__5595 (
            .O(N__29586),
            .I(\control.n16653 ));
    InMux I__5594 (
            .O(N__29583),
            .I(N__29579));
    InMux I__5593 (
            .O(N__29582),
            .I(N__29576));
    LocalMux I__5592 (
            .O(N__29579),
            .I(N__29573));
    LocalMux I__5591 (
            .O(N__29576),
            .I(\control.pwm_delay_8 ));
    Odrv4 I__5590 (
            .O(N__29573),
            .I(\control.pwm_delay_8 ));
    InMux I__5589 (
            .O(N__29568),
            .I(bfn_9_24_0_));
    InMux I__5588 (
            .O(N__29565),
            .I(\control.n16655 ));
    CascadeMux I__5587 (
            .O(N__29562),
            .I(N__29559));
    InMux I__5586 (
            .O(N__29559),
            .I(N__29553));
    InMux I__5585 (
            .O(N__29558),
            .I(N__29553));
    LocalMux I__5584 (
            .O(N__29553),
            .I(data_out_3_7));
    CascadeMux I__5583 (
            .O(N__29550),
            .I(N__29547));
    InMux I__5582 (
            .O(N__29547),
            .I(N__29541));
    InMux I__5581 (
            .O(N__29546),
            .I(N__29541));
    LocalMux I__5580 (
            .O(N__29541),
            .I(data_out_2_7));
    InMux I__5579 (
            .O(N__29538),
            .I(N__29535));
    LocalMux I__5578 (
            .O(N__29535),
            .I(N__29532));
    Odrv4 I__5577 (
            .O(N__29532),
            .I(\c0.n2_adj_2229 ));
    CascadeMux I__5576 (
            .O(N__29529),
            .I(n2837_cascade_));
    InMux I__5575 (
            .O(N__29526),
            .I(N__29522));
    InMux I__5574 (
            .O(N__29525),
            .I(N__29519));
    LocalMux I__5573 (
            .O(N__29522),
            .I(data_out_0_5));
    LocalMux I__5572 (
            .O(N__29519),
            .I(data_out_0_5));
    CascadeMux I__5571 (
            .O(N__29514),
            .I(\control.n12_cascade_ ));
    InMux I__5570 (
            .O(N__29511),
            .I(N__29508));
    LocalMux I__5569 (
            .O(N__29508),
            .I(\control.n10 ));
    InMux I__5568 (
            .O(N__29505),
            .I(bfn_9_23_0_));
    InMux I__5567 (
            .O(N__29502),
            .I(N__29499));
    LocalMux I__5566 (
            .O(N__29499),
            .I(\control.n9_adj_2459 ));
    InMux I__5565 (
            .O(N__29496),
            .I(\control.n16647 ));
    InMux I__5564 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__5563 (
            .O(N__29490),
            .I(N__29487));
    Odrv4 I__5562 (
            .O(N__29487),
            .I(\c0.n18188 ));
    CEMux I__5561 (
            .O(N__29484),
            .I(N__29480));
    CEMux I__5560 (
            .O(N__29483),
            .I(N__29476));
    LocalMux I__5559 (
            .O(N__29480),
            .I(N__29473));
    InMux I__5558 (
            .O(N__29479),
            .I(N__29469));
    LocalMux I__5557 (
            .O(N__29476),
            .I(N__29466));
    Span4Mux_v I__5556 (
            .O(N__29473),
            .I(N__29463));
    InMux I__5555 (
            .O(N__29472),
            .I(N__29460));
    LocalMux I__5554 (
            .O(N__29469),
            .I(N__29457));
    Span4Mux_v I__5553 (
            .O(N__29466),
            .I(N__29450));
    Span4Mux_h I__5552 (
            .O(N__29463),
            .I(N__29450));
    LocalMux I__5551 (
            .O(N__29460),
            .I(N__29450));
    Odrv12 I__5550 (
            .O(N__29457),
            .I(n5155));
    Odrv4 I__5549 (
            .O(N__29450),
            .I(n5155));
    CascadeMux I__5548 (
            .O(N__29445),
            .I(N__29442));
    InMux I__5547 (
            .O(N__29442),
            .I(N__29439));
    LocalMux I__5546 (
            .O(N__29439),
            .I(N__29436));
    Odrv4 I__5545 (
            .O(N__29436),
            .I(\c0.n18354 ));
    InMux I__5544 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__5543 (
            .O(N__29430),
            .I(n18756));
    InMux I__5542 (
            .O(N__29427),
            .I(N__29423));
    InMux I__5541 (
            .O(N__29426),
            .I(N__29420));
    LocalMux I__5540 (
            .O(N__29423),
            .I(N__29417));
    LocalMux I__5539 (
            .O(N__29420),
            .I(\c0.data_out_3_6 ));
    Odrv4 I__5538 (
            .O(N__29417),
            .I(\c0.data_out_3_6 ));
    CascadeMux I__5537 (
            .O(N__29412),
            .I(n10_adj_2532_cascade_));
    InMux I__5536 (
            .O(N__29409),
            .I(N__29403));
    InMux I__5535 (
            .O(N__29408),
            .I(N__29403));
    LocalMux I__5534 (
            .O(N__29403),
            .I(r_Tx_Data_6));
    InMux I__5533 (
            .O(N__29400),
            .I(N__29397));
    LocalMux I__5532 (
            .O(N__29397),
            .I(N__29394));
    Span4Mux_h I__5531 (
            .O(N__29394),
            .I(N__29391));
    Odrv4 I__5530 (
            .O(N__29391),
            .I(\c0.tx.n17984 ));
    CascadeMux I__5529 (
            .O(N__29388),
            .I(n10_adj_2537_cascade_));
    CascadeMux I__5528 (
            .O(N__29385),
            .I(n10_adj_2535_cascade_));
    InMux I__5527 (
            .O(N__29382),
            .I(N__29378));
    InMux I__5526 (
            .O(N__29381),
            .I(N__29375));
    LocalMux I__5525 (
            .O(N__29378),
            .I(r_Tx_Data_7));
    LocalMux I__5524 (
            .O(N__29375),
            .I(r_Tx_Data_7));
    CascadeMux I__5523 (
            .O(N__29370),
            .I(n3_adj_2525_cascade_));
    IoInMux I__5522 (
            .O(N__29367),
            .I(N__29364));
    LocalMux I__5521 (
            .O(N__29364),
            .I(N__29361));
    Span4Mux_s3_h I__5520 (
            .O(N__29361),
            .I(N__29358));
    Span4Mux_v I__5519 (
            .O(N__29358),
            .I(N__29355));
    Span4Mux_v I__5518 (
            .O(N__29355),
            .I(N__29350));
    InMux I__5517 (
            .O(N__29354),
            .I(N__29347));
    InMux I__5516 (
            .O(N__29353),
            .I(N__29344));
    Span4Mux_h I__5515 (
            .O(N__29350),
            .I(N__29341));
    LocalMux I__5514 (
            .O(N__29347),
            .I(N__29338));
    LocalMux I__5513 (
            .O(N__29344),
            .I(N__29335));
    Odrv4 I__5512 (
            .O(N__29341),
            .I(tx_o));
    Odrv4 I__5511 (
            .O(N__29338),
            .I(tx_o));
    Odrv4 I__5510 (
            .O(N__29335),
            .I(tx_o));
    InMux I__5509 (
            .O(N__29328),
            .I(N__29325));
    LocalMux I__5508 (
            .O(N__29325),
            .I(\c0.tx.n17697 ));
    InMux I__5507 (
            .O(N__29322),
            .I(N__29318));
    InMux I__5506 (
            .O(N__29321),
            .I(N__29315));
    LocalMux I__5505 (
            .O(N__29318),
            .I(data_out_1_7));
    LocalMux I__5504 (
            .O(N__29315),
            .I(data_out_1_7));
    CascadeMux I__5503 (
            .O(N__29310),
            .I(\c0.tx.n11030_cascade_ ));
    InMux I__5502 (
            .O(N__29307),
            .I(N__29304));
    LocalMux I__5501 (
            .O(N__29304),
            .I(\c0.tx.n18041 ));
    InMux I__5500 (
            .O(N__29301),
            .I(N__29298));
    LocalMux I__5499 (
            .O(N__29298),
            .I(\c0.tx.o_Tx_Serial_N_2062 ));
    InMux I__5498 (
            .O(N__29295),
            .I(N__29292));
    LocalMux I__5497 (
            .O(N__29292),
            .I(n18750));
    InMux I__5496 (
            .O(N__29289),
            .I(N__29286));
    LocalMux I__5495 (
            .O(N__29286),
            .I(\c0.tx_active_prev ));
    InMux I__5494 (
            .O(N__29283),
            .I(N__29280));
    LocalMux I__5493 (
            .O(N__29280),
            .I(N__29275));
    InMux I__5492 (
            .O(N__29279),
            .I(N__29271));
    InMux I__5491 (
            .O(N__29278),
            .I(N__29268));
    Span4Mux_v I__5490 (
            .O(N__29275),
            .I(N__29265));
    InMux I__5489 (
            .O(N__29274),
            .I(N__29262));
    LocalMux I__5488 (
            .O(N__29271),
            .I(N__29257));
    LocalMux I__5487 (
            .O(N__29268),
            .I(N__29257));
    Odrv4 I__5486 (
            .O(N__29265),
            .I(data_in_1_1));
    LocalMux I__5485 (
            .O(N__29262),
            .I(data_in_1_1));
    Odrv4 I__5484 (
            .O(N__29257),
            .I(data_in_1_1));
    InMux I__5483 (
            .O(N__29250),
            .I(\c0.n16520 ));
    InMux I__5482 (
            .O(N__29247),
            .I(\c0.n16521 ));
    InMux I__5481 (
            .O(N__29244),
            .I(\c0.n16522 ));
    InMux I__5480 (
            .O(N__29241),
            .I(\c0.n16523 ));
    InMux I__5479 (
            .O(N__29238),
            .I(N__29235));
    LocalMux I__5478 (
            .O(N__29235),
            .I(N__29232));
    Span4Mux_h I__5477 (
            .O(N__29232),
            .I(N__29229));
    Span4Mux_v I__5476 (
            .O(N__29229),
            .I(N__29226));
    Odrv4 I__5475 (
            .O(N__29226),
            .I(\c0.n18254 ));
    SRMux I__5474 (
            .O(N__29223),
            .I(N__29220));
    LocalMux I__5473 (
            .O(N__29220),
            .I(N__29217));
    Sp12to4 I__5472 (
            .O(N__29217),
            .I(N__29214));
    Span12Mux_v I__5471 (
            .O(N__29214),
            .I(N__29211));
    Odrv12 I__5470 (
            .O(N__29211),
            .I(\c0.n4_adj_2231 ));
    InMux I__5469 (
            .O(N__29208),
            .I(N__29205));
    LocalMux I__5468 (
            .O(N__29205),
            .I(N__29201));
    InMux I__5467 (
            .O(N__29204),
            .I(N__29197));
    Span4Mux_h I__5466 (
            .O(N__29201),
            .I(N__29194));
    InMux I__5465 (
            .O(N__29200),
            .I(N__29191));
    LocalMux I__5464 (
            .O(N__29197),
            .I(N__29186));
    Span4Mux_v I__5463 (
            .O(N__29194),
            .I(N__29186));
    LocalMux I__5462 (
            .O(N__29191),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__5461 (
            .O(N__29186),
            .I(\c0.rx.r_Clock_Count_7 ));
    InMux I__5460 (
            .O(N__29181),
            .I(N__29178));
    LocalMux I__5459 (
            .O(N__29178),
            .I(N__29174));
    InMux I__5458 (
            .O(N__29177),
            .I(N__29170));
    Span4Mux_h I__5457 (
            .O(N__29174),
            .I(N__29167));
    InMux I__5456 (
            .O(N__29173),
            .I(N__29164));
    LocalMux I__5455 (
            .O(N__29170),
            .I(N__29159));
    Span4Mux_v I__5454 (
            .O(N__29167),
            .I(N__29159));
    LocalMux I__5453 (
            .O(N__29164),
            .I(\c0.rx.r_Clock_Count_6 ));
    Odrv4 I__5452 (
            .O(N__29159),
            .I(\c0.rx.r_Clock_Count_6 ));
    InMux I__5451 (
            .O(N__29154),
            .I(N__29151));
    LocalMux I__5450 (
            .O(N__29151),
            .I(N__29147));
    InMux I__5449 (
            .O(N__29150),
            .I(N__29144));
    Span4Mux_v I__5448 (
            .O(N__29147),
            .I(N__29138));
    LocalMux I__5447 (
            .O(N__29144),
            .I(N__29138));
    InMux I__5446 (
            .O(N__29143),
            .I(N__29135));
    Span4Mux_v I__5445 (
            .O(N__29138),
            .I(N__29130));
    LocalMux I__5444 (
            .O(N__29135),
            .I(N__29130));
    Odrv4 I__5443 (
            .O(N__29130),
            .I(\c0.rx.n73 ));
    InMux I__5442 (
            .O(N__29127),
            .I(N__29124));
    LocalMux I__5441 (
            .O(N__29124),
            .I(\c0.n44 ));
    IoInMux I__5440 (
            .O(N__29121),
            .I(N__29118));
    LocalMux I__5439 (
            .O(N__29118),
            .I(N__29115));
    IoSpan4Mux I__5438 (
            .O(N__29115),
            .I(N__29112));
    IoSpan4Mux I__5437 (
            .O(N__29112),
            .I(N__29109));
    Span4Mux_s3_h I__5436 (
            .O(N__29109),
            .I(N__29106));
    Span4Mux_h I__5435 (
            .O(N__29106),
            .I(N__29103));
    Odrv4 I__5434 (
            .O(N__29103),
            .I(tx_enable));
    InMux I__5433 (
            .O(N__29100),
            .I(\c0.tx2.n16542 ));
    InMux I__5432 (
            .O(N__29097),
            .I(\c0.tx2.n16543 ));
    InMux I__5431 (
            .O(N__29094),
            .I(N__29091));
    LocalMux I__5430 (
            .O(N__29091),
            .I(N__29088));
    Span4Mux_h I__5429 (
            .O(N__29088),
            .I(N__29084));
    InMux I__5428 (
            .O(N__29087),
            .I(N__29081));
    Span4Mux_h I__5427 (
            .O(N__29084),
            .I(N__29078));
    LocalMux I__5426 (
            .O(N__29081),
            .I(\c0.tx2.r_Clock_Count_6 ));
    Odrv4 I__5425 (
            .O(N__29078),
            .I(\c0.tx2.r_Clock_Count_6 ));
    InMux I__5424 (
            .O(N__29073),
            .I(\c0.tx2.n16544 ));
    InMux I__5423 (
            .O(N__29070),
            .I(N__29067));
    LocalMux I__5422 (
            .O(N__29067),
            .I(N__29064));
    Span4Mux_h I__5421 (
            .O(N__29064),
            .I(N__29060));
    InMux I__5420 (
            .O(N__29063),
            .I(N__29057));
    Span4Mux_h I__5419 (
            .O(N__29060),
            .I(N__29054));
    LocalMux I__5418 (
            .O(N__29057),
            .I(\c0.tx2.r_Clock_Count_7 ));
    Odrv4 I__5417 (
            .O(N__29054),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__5416 (
            .O(N__29049),
            .I(\c0.tx2.n16545 ));
    InMux I__5415 (
            .O(N__29046),
            .I(bfn_9_7_0_));
    InMux I__5414 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__5413 (
            .O(N__29040),
            .I(N__29037));
    Span4Mux_h I__5412 (
            .O(N__29037),
            .I(N__29033));
    InMux I__5411 (
            .O(N__29036),
            .I(N__29030));
    Span4Mux_h I__5410 (
            .O(N__29033),
            .I(N__29027));
    LocalMux I__5409 (
            .O(N__29030),
            .I(\c0.tx2.r_Clock_Count_8 ));
    Odrv4 I__5408 (
            .O(N__29027),
            .I(\c0.tx2.r_Clock_Count_8 ));
    SRMux I__5407 (
            .O(N__29022),
            .I(N__29018));
    SRMux I__5406 (
            .O(N__29021),
            .I(N__29015));
    LocalMux I__5405 (
            .O(N__29018),
            .I(N__29012));
    LocalMux I__5404 (
            .O(N__29015),
            .I(N__29009));
    Span4Mux_v I__5403 (
            .O(N__29012),
            .I(N__29006));
    Span4Mux_v I__5402 (
            .O(N__29009),
            .I(N__29003));
    Odrv4 I__5401 (
            .O(N__29006),
            .I(\c0.tx2.n11312 ));
    Odrv4 I__5400 (
            .O(N__29003),
            .I(\c0.tx2.n11312 ));
    InMux I__5399 (
            .O(N__28998),
            .I(\c0.n16517 ));
    InMux I__5398 (
            .O(N__28995),
            .I(\c0.n16518 ));
    InMux I__5397 (
            .O(N__28992),
            .I(\c0.n16519 ));
    InMux I__5396 (
            .O(N__28989),
            .I(N__28977));
    InMux I__5395 (
            .O(N__28988),
            .I(N__28977));
    InMux I__5394 (
            .O(N__28987),
            .I(N__28974));
    InMux I__5393 (
            .O(N__28986),
            .I(N__28971));
    InMux I__5392 (
            .O(N__28985),
            .I(N__28968));
    InMux I__5391 (
            .O(N__28984),
            .I(N__28961));
    InMux I__5390 (
            .O(N__28983),
            .I(N__28961));
    InMux I__5389 (
            .O(N__28982),
            .I(N__28961));
    LocalMux I__5388 (
            .O(N__28977),
            .I(N__28958));
    LocalMux I__5387 (
            .O(N__28974),
            .I(N__28949));
    LocalMux I__5386 (
            .O(N__28971),
            .I(N__28949));
    LocalMux I__5385 (
            .O(N__28968),
            .I(N__28949));
    LocalMux I__5384 (
            .O(N__28961),
            .I(N__28949));
    Span4Mux_h I__5383 (
            .O(N__28958),
            .I(N__28946));
    Span12Mux_s4_v I__5382 (
            .O(N__28949),
            .I(N__28943));
    Odrv4 I__5381 (
            .O(N__28946),
            .I(\c0.n6033 ));
    Odrv12 I__5380 (
            .O(N__28943),
            .I(\c0.n6033 ));
    CascadeMux I__5379 (
            .O(N__28938),
            .I(\c0.n18085_cascade_ ));
    InMux I__5378 (
            .O(N__28935),
            .I(N__28930));
    InMux I__5377 (
            .O(N__28934),
            .I(N__28925));
    InMux I__5376 (
            .O(N__28933),
            .I(N__28925));
    LocalMux I__5375 (
            .O(N__28930),
            .I(N__28921));
    LocalMux I__5374 (
            .O(N__28925),
            .I(N__28916));
    InMux I__5373 (
            .O(N__28924),
            .I(N__28913));
    Span4Mux_h I__5372 (
            .O(N__28921),
            .I(N__28910));
    InMux I__5371 (
            .O(N__28920),
            .I(N__28905));
    InMux I__5370 (
            .O(N__28919),
            .I(N__28905));
    Span4Mux_v I__5369 (
            .O(N__28916),
            .I(N__28900));
    LocalMux I__5368 (
            .O(N__28913),
            .I(N__28900));
    Odrv4 I__5367 (
            .O(N__28910),
            .I(\c0.n4494 ));
    LocalMux I__5366 (
            .O(N__28905),
            .I(\c0.n4494 ));
    Odrv4 I__5365 (
            .O(N__28900),
            .I(\c0.n4494 ));
    InMux I__5364 (
            .O(N__28893),
            .I(N__28887));
    InMux I__5363 (
            .O(N__28892),
            .I(N__28887));
    LocalMux I__5362 (
            .O(N__28887),
            .I(N__28884));
    Span4Mux_h I__5361 (
            .O(N__28884),
            .I(N__28879));
    InMux I__5360 (
            .O(N__28883),
            .I(N__28874));
    InMux I__5359 (
            .O(N__28882),
            .I(N__28874));
    Odrv4 I__5358 (
            .O(N__28879),
            .I(\c0.n28 ));
    LocalMux I__5357 (
            .O(N__28874),
            .I(\c0.n28 ));
    InMux I__5356 (
            .O(N__28869),
            .I(N__28863));
    InMux I__5355 (
            .O(N__28868),
            .I(N__28863));
    LocalMux I__5354 (
            .O(N__28863),
            .I(N__28855));
    InMux I__5353 (
            .O(N__28862),
            .I(N__28850));
    InMux I__5352 (
            .O(N__28861),
            .I(N__28850));
    InMux I__5351 (
            .O(N__28860),
            .I(N__28843));
    InMux I__5350 (
            .O(N__28859),
            .I(N__28843));
    InMux I__5349 (
            .O(N__28858),
            .I(N__28843));
    Odrv4 I__5348 (
            .O(N__28855),
            .I(\c0.n12704 ));
    LocalMux I__5347 (
            .O(N__28850),
            .I(\c0.n12704 ));
    LocalMux I__5346 (
            .O(N__28843),
            .I(\c0.n12704 ));
    InMux I__5345 (
            .O(N__28836),
            .I(N__28833));
    LocalMux I__5344 (
            .O(N__28833),
            .I(N__28830));
    Span4Mux_h I__5343 (
            .O(N__28830),
            .I(N__28827));
    Odrv4 I__5342 (
            .O(N__28827),
            .I(\c0.n18082 ));
    InMux I__5341 (
            .O(N__28824),
            .I(N__28821));
    LocalMux I__5340 (
            .O(N__28821),
            .I(\c0.n18270 ));
    InMux I__5339 (
            .O(N__28818),
            .I(N__28805));
    InMux I__5338 (
            .O(N__28817),
            .I(N__28805));
    InMux I__5337 (
            .O(N__28816),
            .I(N__28805));
    InMux I__5336 (
            .O(N__28815),
            .I(N__28805));
    InMux I__5335 (
            .O(N__28814),
            .I(N__28800));
    LocalMux I__5334 (
            .O(N__28805),
            .I(N__28797));
    CascadeMux I__5333 (
            .O(N__28804),
            .I(N__28794));
    CascadeMux I__5332 (
            .O(N__28803),
            .I(N__28788));
    LocalMux I__5331 (
            .O(N__28800),
            .I(N__28784));
    Span4Mux_h I__5330 (
            .O(N__28797),
            .I(N__28781));
    InMux I__5329 (
            .O(N__28794),
            .I(N__28778));
    InMux I__5328 (
            .O(N__28793),
            .I(N__28767));
    InMux I__5327 (
            .O(N__28792),
            .I(N__28767));
    InMux I__5326 (
            .O(N__28791),
            .I(N__28767));
    InMux I__5325 (
            .O(N__28788),
            .I(N__28767));
    InMux I__5324 (
            .O(N__28787),
            .I(N__28767));
    Odrv12 I__5323 (
            .O(N__28784),
            .I(\c0.n6035 ));
    Odrv4 I__5322 (
            .O(N__28781),
            .I(\c0.n6035 ));
    LocalMux I__5321 (
            .O(N__28778),
            .I(\c0.n6035 ));
    LocalMux I__5320 (
            .O(N__28767),
            .I(\c0.n6035 ));
    InMux I__5319 (
            .O(N__28758),
            .I(bfn_9_6_0_));
    InMux I__5318 (
            .O(N__28755),
            .I(\c0.tx2.n16539 ));
    InMux I__5317 (
            .O(N__28752),
            .I(\c0.tx2.n16540 ));
    InMux I__5316 (
            .O(N__28749),
            .I(\c0.tx2.n16541 ));
    CascadeMux I__5315 (
            .O(N__28746),
            .I(\c0.n18284_cascade_ ));
    InMux I__5314 (
            .O(N__28743),
            .I(N__28740));
    LocalMux I__5313 (
            .O(N__28740),
            .I(N__28737));
    Odrv4 I__5312 (
            .O(N__28737),
            .I(\c0.n27_adj_2405 ));
    InMux I__5311 (
            .O(N__28734),
            .I(N__28731));
    LocalMux I__5310 (
            .O(N__28731),
            .I(N__28728));
    Span4Mux_h I__5309 (
            .O(N__28728),
            .I(N__28725));
    Odrv4 I__5308 (
            .O(N__28725),
            .I(\c0.n29_adj_2408 ));
    CascadeMux I__5307 (
            .O(N__28722),
            .I(\c0.n12704_cascade_ ));
    InMux I__5306 (
            .O(N__28719),
            .I(N__28716));
    LocalMux I__5305 (
            .O(N__28716),
            .I(\c0.n18287 ));
    CascadeMux I__5304 (
            .O(N__28713),
            .I(N__28709));
    CascadeMux I__5303 (
            .O(N__28712),
            .I(N__28706));
    InMux I__5302 (
            .O(N__28709),
            .I(N__28703));
    InMux I__5301 (
            .O(N__28706),
            .I(N__28700));
    LocalMux I__5300 (
            .O(N__28703),
            .I(N__28693));
    LocalMux I__5299 (
            .O(N__28700),
            .I(N__28690));
    InMux I__5298 (
            .O(N__28699),
            .I(N__28681));
    InMux I__5297 (
            .O(N__28698),
            .I(N__28681));
    InMux I__5296 (
            .O(N__28697),
            .I(N__28681));
    InMux I__5295 (
            .O(N__28696),
            .I(N__28681));
    Span4Mux_h I__5294 (
            .O(N__28693),
            .I(N__28678));
    Span4Mux_v I__5293 (
            .O(N__28690),
            .I(N__28675));
    LocalMux I__5292 (
            .O(N__28681),
            .I(N__28672));
    Span4Mux_v I__5291 (
            .O(N__28678),
            .I(N__28669));
    Span4Mux_h I__5290 (
            .O(N__28675),
            .I(N__28664));
    Span4Mux_v I__5289 (
            .O(N__28672),
            .I(N__28664));
    Odrv4 I__5288 (
            .O(N__28669),
            .I(n612));
    Odrv4 I__5287 (
            .O(N__28664),
            .I(n612));
    CascadeMux I__5286 (
            .O(N__28659),
            .I(\c0.n18289_cascade_ ));
    InMux I__5285 (
            .O(N__28656),
            .I(N__28651));
    InMux I__5284 (
            .O(N__28655),
            .I(N__28646));
    InMux I__5283 (
            .O(N__28654),
            .I(N__28646));
    LocalMux I__5282 (
            .O(N__28651),
            .I(\c0.n18831 ));
    LocalMux I__5281 (
            .O(N__28646),
            .I(\c0.n18831 ));
    CascadeMux I__5280 (
            .O(N__28641),
            .I(\c0.n18079_cascade_ ));
    InMux I__5279 (
            .O(N__28638),
            .I(N__28635));
    LocalMux I__5278 (
            .O(N__28635),
            .I(N__28632));
    Odrv12 I__5277 (
            .O(N__28632),
            .I(\c0.n17725 ));
    InMux I__5276 (
            .O(N__28629),
            .I(N__28626));
    LocalMux I__5275 (
            .O(N__28626),
            .I(N__28623));
    Span4Mux_v I__5274 (
            .O(N__28623),
            .I(N__28620));
    Odrv4 I__5273 (
            .O(N__28620),
            .I(\c0.n16863 ));
    CascadeMux I__5272 (
            .O(N__28617),
            .I(N__28614));
    InMux I__5271 (
            .O(N__28614),
            .I(N__28611));
    LocalMux I__5270 (
            .O(N__28611),
            .I(N__28608));
    Odrv4 I__5269 (
            .O(N__28608),
            .I(\c0.n16982 ));
    InMux I__5268 (
            .O(N__28605),
            .I(N__28602));
    LocalMux I__5267 (
            .O(N__28602),
            .I(N__28599));
    Span4Mux_h I__5266 (
            .O(N__28599),
            .I(N__28596));
    Odrv4 I__5265 (
            .O(N__28596),
            .I(\c0.n17722 ));
    CascadeMux I__5264 (
            .O(N__28593),
            .I(N__28590));
    InMux I__5263 (
            .O(N__28590),
            .I(N__28587));
    LocalMux I__5262 (
            .O(N__28587),
            .I(\c0.n28_adj_2403 ));
    CascadeMux I__5261 (
            .O(N__28584),
            .I(n17689_cascade_));
    InMux I__5260 (
            .O(N__28581),
            .I(N__28578));
    LocalMux I__5259 (
            .O(N__28578),
            .I(\c0.n18684 ));
    InMux I__5258 (
            .O(N__28575),
            .I(N__28572));
    LocalMux I__5257 (
            .O(N__28572),
            .I(N__28569));
    Odrv4 I__5256 (
            .O(N__28569),
            .I(\c0.n18072 ));
    CascadeMux I__5255 (
            .O(N__28566),
            .I(\c0.tx2.n14_cascade_ ));
    InMux I__5254 (
            .O(N__28563),
            .I(N__28560));
    LocalMux I__5253 (
            .O(N__28560),
            .I(\c0.n18843 ));
    CascadeMux I__5252 (
            .O(N__28557),
            .I(\c0.n18846_cascade_ ));
    InMux I__5251 (
            .O(N__28554),
            .I(N__28551));
    LocalMux I__5250 (
            .O(N__28551),
            .I(\c0.n22_adj_2239 ));
    InMux I__5249 (
            .O(N__28548),
            .I(N__28545));
    LocalMux I__5248 (
            .O(N__28545),
            .I(N__28542));
    Span4Mux_h I__5247 (
            .O(N__28542),
            .I(N__28539));
    Span4Mux_h I__5246 (
            .O(N__28539),
            .I(N__28536));
    Span4Mux_v I__5245 (
            .O(N__28536),
            .I(N__28533));
    Odrv4 I__5244 (
            .O(N__28533),
            .I(\c0.tx2.r_Tx_Data_7 ));
    CascadeMux I__5243 (
            .O(N__28530),
            .I(\c0.n18675_cascade_ ));
    CascadeMux I__5242 (
            .O(N__28527),
            .I(\c0.n18678_cascade_ ));
    CascadeMux I__5241 (
            .O(N__28524),
            .I(\c0.n18741_cascade_ ));
    InMux I__5240 (
            .O(N__28521),
            .I(N__28518));
    LocalMux I__5239 (
            .O(N__28518),
            .I(\c0.n22_adj_2242 ));
    CascadeMux I__5238 (
            .O(N__28515),
            .I(\c0.n18744_cascade_ ));
    InMux I__5237 (
            .O(N__28512),
            .I(N__28509));
    LocalMux I__5236 (
            .O(N__28509),
            .I(N__28506));
    Span4Mux_v I__5235 (
            .O(N__28506),
            .I(N__28503));
    Span4Mux_h I__5234 (
            .O(N__28503),
            .I(N__28500));
    Odrv4 I__5233 (
            .O(N__28500),
            .I(\c0.tx2.r_Tx_Data_5 ));
    InMux I__5232 (
            .O(N__28497),
            .I(bfn_7_16_0_));
    InMux I__5231 (
            .O(N__28494),
            .I(N__28490));
    InMux I__5230 (
            .O(N__28493),
            .I(N__28487));
    LocalMux I__5229 (
            .O(N__28490),
            .I(N__28484));
    LocalMux I__5228 (
            .O(N__28487),
            .I(\c0.tx.r_Clock_Count_8 ));
    Odrv4 I__5227 (
            .O(N__28484),
            .I(\c0.tx.r_Clock_Count_8 ));
    SRMux I__5226 (
            .O(N__28479),
            .I(N__28476));
    LocalMux I__5225 (
            .O(N__28476),
            .I(N__28472));
    SRMux I__5224 (
            .O(N__28475),
            .I(N__28469));
    Sp12to4 I__5223 (
            .O(N__28472),
            .I(N__28464));
    LocalMux I__5222 (
            .O(N__28469),
            .I(N__28464));
    Odrv12 I__5221 (
            .O(N__28464),
            .I(\c0.tx.n11297 ));
    InMux I__5220 (
            .O(N__28461),
            .I(N__28457));
    InMux I__5219 (
            .O(N__28460),
            .I(N__28454));
    LocalMux I__5218 (
            .O(N__28457),
            .I(\control.n8 ));
    LocalMux I__5217 (
            .O(N__28454),
            .I(\control.n8 ));
    CascadeMux I__5216 (
            .O(N__28449),
            .I(\control.PHASES_5_N_2152_1_cascade_ ));
    SRMux I__5215 (
            .O(N__28446),
            .I(N__28443));
    LocalMux I__5214 (
            .O(N__28443),
            .I(\control.n10356 ));
    CascadeMux I__5213 (
            .O(N__28440),
            .I(\c0.n18801_cascade_ ));
    InMux I__5212 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__5211 (
            .O(N__28434),
            .I(\c0.n18804 ));
    InMux I__5210 (
            .O(N__28431),
            .I(N__28428));
    LocalMux I__5209 (
            .O(N__28428),
            .I(\c0.tx.n54 ));
    CascadeMux I__5208 (
            .O(N__28425),
            .I(\c0.tx.n47_cascade_ ));
    CascadeMux I__5207 (
            .O(N__28422),
            .I(N__28418));
    InMux I__5206 (
            .O(N__28421),
            .I(N__28414));
    InMux I__5205 (
            .O(N__28418),
            .I(N__28409));
    InMux I__5204 (
            .O(N__28417),
            .I(N__28409));
    LocalMux I__5203 (
            .O(N__28414),
            .I(\c0.tx.r_Clock_Count_0 ));
    LocalMux I__5202 (
            .O(N__28409),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__5201 (
            .O(N__28404),
            .I(bfn_7_15_0_));
    InMux I__5200 (
            .O(N__28401),
            .I(N__28397));
    InMux I__5199 (
            .O(N__28400),
            .I(N__28394));
    LocalMux I__5198 (
            .O(N__28397),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__5197 (
            .O(N__28394),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__5196 (
            .O(N__28389),
            .I(\c0.tx.n16524 ));
    CascadeMux I__5195 (
            .O(N__28386),
            .I(N__28382));
    InMux I__5194 (
            .O(N__28385),
            .I(N__28379));
    InMux I__5193 (
            .O(N__28382),
            .I(N__28376));
    LocalMux I__5192 (
            .O(N__28379),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__5191 (
            .O(N__28376),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__5190 (
            .O(N__28371),
            .I(\c0.tx.n16525 ));
    InMux I__5189 (
            .O(N__28368),
            .I(N__28363));
    InMux I__5188 (
            .O(N__28367),
            .I(N__28358));
    InMux I__5187 (
            .O(N__28366),
            .I(N__28358));
    LocalMux I__5186 (
            .O(N__28363),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__5185 (
            .O(N__28358),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__5184 (
            .O(N__28353),
            .I(\c0.tx.n16526 ));
    InMux I__5183 (
            .O(N__28350),
            .I(N__28346));
    InMux I__5182 (
            .O(N__28349),
            .I(N__28343));
    LocalMux I__5181 (
            .O(N__28346),
            .I(\c0.tx.r_Clock_Count_4 ));
    LocalMux I__5180 (
            .O(N__28343),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__5179 (
            .O(N__28338),
            .I(\c0.tx.n16527 ));
    InMux I__5178 (
            .O(N__28335),
            .I(N__28331));
    InMux I__5177 (
            .O(N__28334),
            .I(N__28328));
    LocalMux I__5176 (
            .O(N__28331),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__5175 (
            .O(N__28328),
            .I(\c0.tx.r_Clock_Count_5 ));
    InMux I__5174 (
            .O(N__28323),
            .I(\c0.tx.n16528 ));
    InMux I__5173 (
            .O(N__28320),
            .I(N__28316));
    InMux I__5172 (
            .O(N__28319),
            .I(N__28313));
    LocalMux I__5171 (
            .O(N__28316),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__5170 (
            .O(N__28313),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__5169 (
            .O(N__28308),
            .I(\c0.tx.n16529 ));
    InMux I__5168 (
            .O(N__28305),
            .I(N__28301));
    InMux I__5167 (
            .O(N__28304),
            .I(N__28298));
    LocalMux I__5166 (
            .O(N__28301),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__5165 (
            .O(N__28298),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__5164 (
            .O(N__28293),
            .I(\c0.tx.n16530 ));
    CascadeMux I__5163 (
            .O(N__28290),
            .I(\c0.rx.n18024_cascade_ ));
    InMux I__5162 (
            .O(N__28287),
            .I(N__28283));
    InMux I__5161 (
            .O(N__28286),
            .I(N__28280));
    LocalMux I__5160 (
            .O(N__28283),
            .I(N__28277));
    LocalMux I__5159 (
            .O(N__28280),
            .I(\c0.rx.n12828 ));
    Odrv12 I__5158 (
            .O(N__28277),
            .I(\c0.rx.n12828 ));
    CascadeMux I__5157 (
            .O(N__28272),
            .I(\c0.rx.n12828_cascade_ ));
    InMux I__5156 (
            .O(N__28269),
            .I(N__28266));
    LocalMux I__5155 (
            .O(N__28266),
            .I(N__28263));
    Odrv4 I__5154 (
            .O(N__28263),
            .I(\c0.rx.n18303 ));
    CascadeMux I__5153 (
            .O(N__28260),
            .I(N__28257));
    InMux I__5152 (
            .O(N__28257),
            .I(N__28254));
    LocalMux I__5151 (
            .O(N__28254),
            .I(N__28247));
    InMux I__5150 (
            .O(N__28253),
            .I(N__28244));
    InMux I__5149 (
            .O(N__28252),
            .I(N__28239));
    InMux I__5148 (
            .O(N__28251),
            .I(N__28239));
    InMux I__5147 (
            .O(N__28250),
            .I(N__28236));
    Span4Mux_h I__5146 (
            .O(N__28247),
            .I(N__28233));
    LocalMux I__5145 (
            .O(N__28244),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__5144 (
            .O(N__28239),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__5143 (
            .O(N__28236),
            .I(\c0.rx.r_Clock_Count_5 ));
    Odrv4 I__5142 (
            .O(N__28233),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__5141 (
            .O(N__28224),
            .I(N__28219));
    InMux I__5140 (
            .O(N__28223),
            .I(N__28216));
    InMux I__5139 (
            .O(N__28222),
            .I(N__28213));
    LocalMux I__5138 (
            .O(N__28219),
            .I(N__28210));
    LocalMux I__5137 (
            .O(N__28216),
            .I(N__28207));
    LocalMux I__5136 (
            .O(N__28213),
            .I(\c0.rx.n15902 ));
    Odrv4 I__5135 (
            .O(N__28210),
            .I(\c0.rx.n15902 ));
    Odrv4 I__5134 (
            .O(N__28207),
            .I(\c0.rx.n15902 ));
    InMux I__5133 (
            .O(N__28200),
            .I(N__28193));
    InMux I__5132 (
            .O(N__28199),
            .I(N__28190));
    InMux I__5131 (
            .O(N__28198),
            .I(N__28185));
    InMux I__5130 (
            .O(N__28197),
            .I(N__28185));
    CascadeMux I__5129 (
            .O(N__28196),
            .I(N__28182));
    LocalMux I__5128 (
            .O(N__28193),
            .I(N__28179));
    LocalMux I__5127 (
            .O(N__28190),
            .I(N__28174));
    LocalMux I__5126 (
            .O(N__28185),
            .I(N__28174));
    InMux I__5125 (
            .O(N__28182),
            .I(N__28171));
    Span4Mux_h I__5124 (
            .O(N__28179),
            .I(N__28168));
    Odrv4 I__5123 (
            .O(N__28174),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__5122 (
            .O(N__28171),
            .I(\c0.rx.r_Clock_Count_0 ));
    Odrv4 I__5121 (
            .O(N__28168),
            .I(\c0.rx.r_Clock_Count_0 ));
    InMux I__5120 (
            .O(N__28161),
            .I(N__28158));
    LocalMux I__5119 (
            .O(N__28158),
            .I(\c0.rx.n18211 ));
    CascadeMux I__5118 (
            .O(N__28155),
            .I(N__28151));
    CascadeMux I__5117 (
            .O(N__28154),
            .I(N__28145));
    InMux I__5116 (
            .O(N__28151),
            .I(N__28140));
    InMux I__5115 (
            .O(N__28150),
            .I(N__28140));
    InMux I__5114 (
            .O(N__28149),
            .I(N__28132));
    InMux I__5113 (
            .O(N__28148),
            .I(N__28127));
    InMux I__5112 (
            .O(N__28145),
            .I(N__28127));
    LocalMux I__5111 (
            .O(N__28140),
            .I(N__28124));
    CascadeMux I__5110 (
            .O(N__28139),
            .I(N__28120));
    CascadeMux I__5109 (
            .O(N__28138),
            .I(N__28114));
    CascadeMux I__5108 (
            .O(N__28137),
            .I(N__28111));
    CascadeMux I__5107 (
            .O(N__28136),
            .I(N__28108));
    CascadeMux I__5106 (
            .O(N__28135),
            .I(N__28103));
    LocalMux I__5105 (
            .O(N__28132),
            .I(N__28095));
    LocalMux I__5104 (
            .O(N__28127),
            .I(N__28095));
    Span4Mux_v I__5103 (
            .O(N__28124),
            .I(N__28095));
    InMux I__5102 (
            .O(N__28123),
            .I(N__28090));
    InMux I__5101 (
            .O(N__28120),
            .I(N__28090));
    InMux I__5100 (
            .O(N__28119),
            .I(N__28087));
    CascadeMux I__5099 (
            .O(N__28118),
            .I(N__28083));
    InMux I__5098 (
            .O(N__28117),
            .I(N__28077));
    InMux I__5097 (
            .O(N__28114),
            .I(N__28077));
    InMux I__5096 (
            .O(N__28111),
            .I(N__28070));
    InMux I__5095 (
            .O(N__28108),
            .I(N__28070));
    InMux I__5094 (
            .O(N__28107),
            .I(N__28070));
    InMux I__5093 (
            .O(N__28106),
            .I(N__28063));
    InMux I__5092 (
            .O(N__28103),
            .I(N__28063));
    InMux I__5091 (
            .O(N__28102),
            .I(N__28063));
    Span4Mux_v I__5090 (
            .O(N__28095),
            .I(N__28056));
    LocalMux I__5089 (
            .O(N__28090),
            .I(N__28056));
    LocalMux I__5088 (
            .O(N__28087),
            .I(N__28056));
    InMux I__5087 (
            .O(N__28086),
            .I(N__28053));
    InMux I__5086 (
            .O(N__28083),
            .I(N__28050));
    InMux I__5085 (
            .O(N__28082),
            .I(N__28047));
    LocalMux I__5084 (
            .O(N__28077),
            .I(N__28042));
    LocalMux I__5083 (
            .O(N__28070),
            .I(N__28042));
    LocalMux I__5082 (
            .O(N__28063),
            .I(N__28037));
    Span4Mux_v I__5081 (
            .O(N__28056),
            .I(N__28037));
    LocalMux I__5080 (
            .O(N__28053),
            .I(N__28034));
    LocalMux I__5079 (
            .O(N__28050),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__5078 (
            .O(N__28047),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv12 I__5077 (
            .O(N__28042),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__5076 (
            .O(N__28037),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__5075 (
            .O(N__28034),
            .I(\c0.rx.r_SM_Main_1 ));
    InMux I__5074 (
            .O(N__28023),
            .I(N__28015));
    InMux I__5073 (
            .O(N__28022),
            .I(N__28015));
    InMux I__5072 (
            .O(N__28021),
            .I(N__28012));
    InMux I__5071 (
            .O(N__28020),
            .I(N__28007));
    LocalMux I__5070 (
            .O(N__28015),
            .I(N__28000));
    LocalMux I__5069 (
            .O(N__28012),
            .I(N__28000));
    InMux I__5068 (
            .O(N__28011),
            .I(N__27994));
    InMux I__5067 (
            .O(N__28010),
            .I(N__27994));
    LocalMux I__5066 (
            .O(N__28007),
            .I(N__27990));
    InMux I__5065 (
            .O(N__28006),
            .I(N__27985));
    InMux I__5064 (
            .O(N__28005),
            .I(N__27985));
    Span4Mux_v I__5063 (
            .O(N__28000),
            .I(N__27982));
    InMux I__5062 (
            .O(N__27999),
            .I(N__27978));
    LocalMux I__5061 (
            .O(N__27994),
            .I(N__27975));
    InMux I__5060 (
            .O(N__27993),
            .I(N__27972));
    Span4Mux_v I__5059 (
            .O(N__27990),
            .I(N__27965));
    LocalMux I__5058 (
            .O(N__27985),
            .I(N__27965));
    Span4Mux_v I__5057 (
            .O(N__27982),
            .I(N__27965));
    InMux I__5056 (
            .O(N__27981),
            .I(N__27962));
    LocalMux I__5055 (
            .O(N__27978),
            .I(N__27959));
    Odrv12 I__5054 (
            .O(N__27975),
            .I(r_Rx_Data));
    LocalMux I__5053 (
            .O(N__27972),
            .I(r_Rx_Data));
    Odrv4 I__5052 (
            .O(N__27965),
            .I(r_Rx_Data));
    LocalMux I__5051 (
            .O(N__27962),
            .I(r_Rx_Data));
    Odrv4 I__5050 (
            .O(N__27959),
            .I(r_Rx_Data));
    InMux I__5049 (
            .O(N__27948),
            .I(N__27935));
    InMux I__5048 (
            .O(N__27947),
            .I(N__27930));
    InMux I__5047 (
            .O(N__27946),
            .I(N__27930));
    InMux I__5046 (
            .O(N__27945),
            .I(N__27927));
    InMux I__5045 (
            .O(N__27944),
            .I(N__27921));
    InMux I__5044 (
            .O(N__27943),
            .I(N__27921));
    InMux I__5043 (
            .O(N__27942),
            .I(N__27911));
    InMux I__5042 (
            .O(N__27941),
            .I(N__27911));
    InMux I__5041 (
            .O(N__27940),
            .I(N__27911));
    InMux I__5040 (
            .O(N__27939),
            .I(N__27911));
    InMux I__5039 (
            .O(N__27938),
            .I(N__27908));
    LocalMux I__5038 (
            .O(N__27935),
            .I(N__27901));
    LocalMux I__5037 (
            .O(N__27930),
            .I(N__27901));
    LocalMux I__5036 (
            .O(N__27927),
            .I(N__27901));
    InMux I__5035 (
            .O(N__27926),
            .I(N__27898));
    LocalMux I__5034 (
            .O(N__27921),
            .I(N__27895));
    InMux I__5033 (
            .O(N__27920),
            .I(N__27892));
    LocalMux I__5032 (
            .O(N__27911),
            .I(N__27889));
    LocalMux I__5031 (
            .O(N__27908),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv12 I__5030 (
            .O(N__27901),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__5029 (
            .O(N__27898),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__5028 (
            .O(N__27895),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__5027 (
            .O(N__27892),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv12 I__5026 (
            .O(N__27889),
            .I(\c0.rx.r_SM_Main_0 ));
    InMux I__5025 (
            .O(N__27876),
            .I(N__27873));
    LocalMux I__5024 (
            .O(N__27873),
            .I(\c0.rx.n4 ));
    CascadeMux I__5023 (
            .O(N__27870),
            .I(\c0.tx.n54_cascade_ ));
    InMux I__5022 (
            .O(N__27867),
            .I(N__27861));
    InMux I__5021 (
            .O(N__27866),
            .I(N__27861));
    LocalMux I__5020 (
            .O(N__27861),
            .I(\c0.tx.n10 ));
    InMux I__5019 (
            .O(N__27858),
            .I(N__27850));
    CascadeMux I__5018 (
            .O(N__27857),
            .I(N__27847));
    InMux I__5017 (
            .O(N__27856),
            .I(N__27842));
    InMux I__5016 (
            .O(N__27855),
            .I(N__27837));
    InMux I__5015 (
            .O(N__27854),
            .I(N__27837));
    InMux I__5014 (
            .O(N__27853),
            .I(N__27834));
    LocalMux I__5013 (
            .O(N__27850),
            .I(N__27831));
    InMux I__5012 (
            .O(N__27847),
            .I(N__27828));
    InMux I__5011 (
            .O(N__27846),
            .I(N__27823));
    InMux I__5010 (
            .O(N__27845),
            .I(N__27823));
    LocalMux I__5009 (
            .O(N__27842),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__5008 (
            .O(N__27837),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__5007 (
            .O(N__27834),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv4 I__5006 (
            .O(N__27831),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__5005 (
            .O(N__27828),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__5004 (
            .O(N__27823),
            .I(\c0.rx.r_Bit_Index_2 ));
    InMux I__5003 (
            .O(N__27810),
            .I(N__27804));
    InMux I__5002 (
            .O(N__27809),
            .I(N__27801));
    InMux I__5001 (
            .O(N__27808),
            .I(N__27798));
    CascadeMux I__5000 (
            .O(N__27807),
            .I(N__27793));
    LocalMux I__4999 (
            .O(N__27804),
            .I(N__27790));
    LocalMux I__4998 (
            .O(N__27801),
            .I(N__27785));
    LocalMux I__4997 (
            .O(N__27798),
            .I(N__27785));
    InMux I__4996 (
            .O(N__27797),
            .I(N__27782));
    InMux I__4995 (
            .O(N__27796),
            .I(N__27779));
    InMux I__4994 (
            .O(N__27793),
            .I(N__27776));
    Span4Mux_v I__4993 (
            .O(N__27790),
            .I(N__27773));
    Span4Mux_v I__4992 (
            .O(N__27785),
            .I(N__27770));
    LocalMux I__4991 (
            .O(N__27782),
            .I(N__27763));
    LocalMux I__4990 (
            .O(N__27779),
            .I(N__27763));
    LocalMux I__4989 (
            .O(N__27776),
            .I(N__27763));
    Span4Mux_h I__4988 (
            .O(N__27773),
            .I(N__27758));
    Span4Mux_h I__4987 (
            .O(N__27770),
            .I(N__27758));
    Odrv12 I__4986 (
            .O(N__27763),
            .I(\c0.rx.n167 ));
    Odrv4 I__4985 (
            .O(N__27758),
            .I(\c0.rx.n167 ));
    InMux I__4984 (
            .O(N__27753),
            .I(N__27749));
    InMux I__4983 (
            .O(N__27752),
            .I(N__27745));
    LocalMux I__4982 (
            .O(N__27749),
            .I(N__27742));
    InMux I__4981 (
            .O(N__27748),
            .I(N__27739));
    LocalMux I__4980 (
            .O(N__27745),
            .I(N__27736));
    Odrv4 I__4979 (
            .O(N__27742),
            .I(n12527));
    LocalMux I__4978 (
            .O(N__27739),
            .I(n12527));
    Odrv4 I__4977 (
            .O(N__27736),
            .I(n12527));
    InMux I__4976 (
            .O(N__27729),
            .I(N__27722));
    InMux I__4975 (
            .O(N__27728),
            .I(N__27722));
    InMux I__4974 (
            .O(N__27727),
            .I(N__27719));
    LocalMux I__4973 (
            .O(N__27722),
            .I(data_in_0_0));
    LocalMux I__4972 (
            .O(N__27719),
            .I(data_in_0_0));
    InMux I__4971 (
            .O(N__27714),
            .I(N__27704));
    InMux I__4970 (
            .O(N__27713),
            .I(N__27704));
    InMux I__4969 (
            .O(N__27712),
            .I(N__27704));
    InMux I__4968 (
            .O(N__27711),
            .I(N__27701));
    LocalMux I__4967 (
            .O(N__27704),
            .I(data_in_3_7));
    LocalMux I__4966 (
            .O(N__27701),
            .I(data_in_3_7));
    InMux I__4965 (
            .O(N__27696),
            .I(N__27693));
    LocalMux I__4964 (
            .O(N__27693),
            .I(\c0.n6_adj_2368 ));
    InMux I__4963 (
            .O(N__27690),
            .I(N__27685));
    InMux I__4962 (
            .O(N__27689),
            .I(N__27680));
    InMux I__4961 (
            .O(N__27688),
            .I(N__27680));
    LocalMux I__4960 (
            .O(N__27685),
            .I(data_in_1_3));
    LocalMux I__4959 (
            .O(N__27680),
            .I(data_in_1_3));
    InMux I__4958 (
            .O(N__27675),
            .I(N__27670));
    InMux I__4957 (
            .O(N__27674),
            .I(N__27665));
    InMux I__4956 (
            .O(N__27673),
            .I(N__27665));
    LocalMux I__4955 (
            .O(N__27670),
            .I(data_in_0_3));
    LocalMux I__4954 (
            .O(N__27665),
            .I(data_in_0_3));
    InMux I__4953 (
            .O(N__27660),
            .I(N__27655));
    InMux I__4952 (
            .O(N__27659),
            .I(N__27650));
    InMux I__4951 (
            .O(N__27658),
            .I(N__27650));
    LocalMux I__4950 (
            .O(N__27655),
            .I(data_in_0_1));
    LocalMux I__4949 (
            .O(N__27650),
            .I(data_in_0_1));
    InMux I__4948 (
            .O(N__27645),
            .I(N__27642));
    LocalMux I__4947 (
            .O(N__27642),
            .I(\c0.rx.n18196 ));
    InMux I__4946 (
            .O(N__27639),
            .I(N__27636));
    LocalMux I__4945 (
            .O(N__27636),
            .I(N__27633));
    Odrv12 I__4944 (
            .O(N__27633),
            .I(\c0.rx.n18194 ));
    CascadeMux I__4943 (
            .O(N__27630),
            .I(\c0.rx.n12552_cascade_ ));
    CascadeMux I__4942 (
            .O(N__27627),
            .I(N__27624));
    InMux I__4941 (
            .O(N__27624),
            .I(N__27617));
    InMux I__4940 (
            .O(N__27623),
            .I(N__27614));
    InMux I__4939 (
            .O(N__27622),
            .I(N__27611));
    InMux I__4938 (
            .O(N__27621),
            .I(N__27608));
    InMux I__4937 (
            .O(N__27620),
            .I(N__27605));
    LocalMux I__4936 (
            .O(N__27617),
            .I(N__27599));
    LocalMux I__4935 (
            .O(N__27614),
            .I(N__27599));
    LocalMux I__4934 (
            .O(N__27611),
            .I(N__27596));
    LocalMux I__4933 (
            .O(N__27608),
            .I(N__27591));
    LocalMux I__4932 (
            .O(N__27605),
            .I(N__27591));
    InMux I__4931 (
            .O(N__27604),
            .I(N__27588));
    Span4Mux_v I__4930 (
            .O(N__27599),
            .I(N__27579));
    Span4Mux_v I__4929 (
            .O(N__27596),
            .I(N__27579));
    Span4Mux_h I__4928 (
            .O(N__27591),
            .I(N__27579));
    LocalMux I__4927 (
            .O(N__27588),
            .I(N__27576));
    InMux I__4926 (
            .O(N__27587),
            .I(N__27573));
    CascadeMux I__4925 (
            .O(N__27586),
            .I(N__27569));
    Span4Mux_v I__4924 (
            .O(N__27579),
            .I(N__27566));
    Span4Mux_v I__4923 (
            .O(N__27576),
            .I(N__27561));
    LocalMux I__4922 (
            .O(N__27573),
            .I(N__27561));
    InMux I__4921 (
            .O(N__27572),
            .I(N__27556));
    InMux I__4920 (
            .O(N__27569),
            .I(N__27556));
    Odrv4 I__4919 (
            .O(N__27566),
            .I(rx_data_6));
    Odrv4 I__4918 (
            .O(N__27561),
            .I(rx_data_6));
    LocalMux I__4917 (
            .O(N__27556),
            .I(rx_data_6));
    InMux I__4916 (
            .O(N__27549),
            .I(N__27544));
    CascadeMux I__4915 (
            .O(N__27548),
            .I(N__27536));
    CascadeMux I__4914 (
            .O(N__27547),
            .I(N__27533));
    LocalMux I__4913 (
            .O(N__27544),
            .I(N__27530));
    InMux I__4912 (
            .O(N__27543),
            .I(N__27523));
    InMux I__4911 (
            .O(N__27542),
            .I(N__27523));
    InMux I__4910 (
            .O(N__27541),
            .I(N__27520));
    CascadeMux I__4909 (
            .O(N__27540),
            .I(N__27517));
    InMux I__4908 (
            .O(N__27539),
            .I(N__27514));
    InMux I__4907 (
            .O(N__27536),
            .I(N__27511));
    InMux I__4906 (
            .O(N__27533),
            .I(N__27507));
    Span4Mux_h I__4905 (
            .O(N__27530),
            .I(N__27504));
    InMux I__4904 (
            .O(N__27529),
            .I(N__27501));
    InMux I__4903 (
            .O(N__27528),
            .I(N__27498));
    LocalMux I__4902 (
            .O(N__27523),
            .I(N__27493));
    LocalMux I__4901 (
            .O(N__27520),
            .I(N__27493));
    InMux I__4900 (
            .O(N__27517),
            .I(N__27490));
    LocalMux I__4899 (
            .O(N__27514),
            .I(N__27487));
    LocalMux I__4898 (
            .O(N__27511),
            .I(N__27484));
    InMux I__4897 (
            .O(N__27510),
            .I(N__27481));
    LocalMux I__4896 (
            .O(N__27507),
            .I(N__27474));
    Span4Mux_v I__4895 (
            .O(N__27504),
            .I(N__27474));
    LocalMux I__4894 (
            .O(N__27501),
            .I(N__27474));
    LocalMux I__4893 (
            .O(N__27498),
            .I(N__27469));
    Span4Mux_h I__4892 (
            .O(N__27493),
            .I(N__27469));
    LocalMux I__4891 (
            .O(N__27490),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv12 I__4890 (
            .O(N__27487),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__4889 (
            .O(N__27484),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__4888 (
            .O(N__27481),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__4887 (
            .O(N__27474),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__4886 (
            .O(N__27469),
            .I(\c0.rx.r_Bit_Index_1 ));
    InMux I__4885 (
            .O(N__27456),
            .I(N__27452));
    InMux I__4884 (
            .O(N__27455),
            .I(N__27444));
    LocalMux I__4883 (
            .O(N__27452),
            .I(N__27441));
    InMux I__4882 (
            .O(N__27451),
            .I(N__27436));
    InMux I__4881 (
            .O(N__27450),
            .I(N__27436));
    CascadeMux I__4880 (
            .O(N__27449),
            .I(N__27431));
    InMux I__4879 (
            .O(N__27448),
            .I(N__27423));
    InMux I__4878 (
            .O(N__27447),
            .I(N__27423));
    LocalMux I__4877 (
            .O(N__27444),
            .I(N__27416));
    Span4Mux_v I__4876 (
            .O(N__27441),
            .I(N__27416));
    LocalMux I__4875 (
            .O(N__27436),
            .I(N__27416));
    InMux I__4874 (
            .O(N__27435),
            .I(N__27411));
    InMux I__4873 (
            .O(N__27434),
            .I(N__27411));
    InMux I__4872 (
            .O(N__27431),
            .I(N__27405));
    InMux I__4871 (
            .O(N__27430),
            .I(N__27405));
    InMux I__4870 (
            .O(N__27429),
            .I(N__27402));
    InMux I__4869 (
            .O(N__27428),
            .I(N__27399));
    LocalMux I__4868 (
            .O(N__27423),
            .I(N__27396));
    Span4Mux_v I__4867 (
            .O(N__27416),
            .I(N__27391));
    LocalMux I__4866 (
            .O(N__27411),
            .I(N__27391));
    InMux I__4865 (
            .O(N__27410),
            .I(N__27388));
    LocalMux I__4864 (
            .O(N__27405),
            .I(N__27385));
    LocalMux I__4863 (
            .O(N__27402),
            .I(\c0.rx.r_SM_Main_2 ));
    LocalMux I__4862 (
            .O(N__27399),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv12 I__4861 (
            .O(N__27396),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv4 I__4860 (
            .O(N__27391),
            .I(\c0.rx.r_SM_Main_2 ));
    LocalMux I__4859 (
            .O(N__27388),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv12 I__4858 (
            .O(N__27385),
            .I(\c0.rx.r_SM_Main_2 ));
    InMux I__4857 (
            .O(N__27372),
            .I(N__27366));
    InMux I__4856 (
            .O(N__27371),
            .I(N__27366));
    LocalMux I__4855 (
            .O(N__27366),
            .I(N__27363));
    Span4Mux_h I__4854 (
            .O(N__27363),
            .I(N__27360));
    Span4Mux_v I__4853 (
            .O(N__27360),
            .I(N__27357));
    Odrv4 I__4852 (
            .O(N__27357),
            .I(n164_adj_2464));
    InMux I__4851 (
            .O(N__27354),
            .I(N__27349));
    InMux I__4850 (
            .O(N__27353),
            .I(N__27346));
    InMux I__4849 (
            .O(N__27352),
            .I(N__27343));
    LocalMux I__4848 (
            .O(N__27349),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__4847 (
            .O(N__27346),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__4846 (
            .O(N__27343),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__4845 (
            .O(N__27336),
            .I(N__27331));
    InMux I__4844 (
            .O(N__27335),
            .I(N__27328));
    InMux I__4843 (
            .O(N__27334),
            .I(N__27325));
    LocalMux I__4842 (
            .O(N__27331),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__4841 (
            .O(N__27328),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__4840 (
            .O(N__27325),
            .I(\c0.rx.r_Clock_Count_2 ));
    CascadeMux I__4839 (
            .O(N__27318),
            .I(N__27313));
    InMux I__4838 (
            .O(N__27317),
            .I(N__27310));
    InMux I__4837 (
            .O(N__27316),
            .I(N__27307));
    InMux I__4836 (
            .O(N__27313),
            .I(N__27304));
    LocalMux I__4835 (
            .O(N__27310),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__4834 (
            .O(N__27307),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__4833 (
            .O(N__27304),
            .I(\c0.rx.r_Clock_Count_3 ));
    CascadeMux I__4832 (
            .O(N__27297),
            .I(\c0.rx.n17990_cascade_ ));
    InMux I__4831 (
            .O(N__27294),
            .I(N__27289));
    InMux I__4830 (
            .O(N__27293),
            .I(N__27286));
    InMux I__4829 (
            .O(N__27292),
            .I(N__27283));
    LocalMux I__4828 (
            .O(N__27289),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__4827 (
            .O(N__27286),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__4826 (
            .O(N__27283),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__4825 (
            .O(N__27276),
            .I(N__27271));
    InMux I__4824 (
            .O(N__27275),
            .I(N__27268));
    InMux I__4823 (
            .O(N__27274),
            .I(N__27265));
    LocalMux I__4822 (
            .O(N__27271),
            .I(data_in_2_6));
    LocalMux I__4821 (
            .O(N__27268),
            .I(data_in_2_6));
    LocalMux I__4820 (
            .O(N__27265),
            .I(data_in_2_6));
    InMux I__4819 (
            .O(N__27258),
            .I(N__27255));
    LocalMux I__4818 (
            .O(N__27255),
            .I(N__27249));
    InMux I__4817 (
            .O(N__27254),
            .I(N__27246));
    InMux I__4816 (
            .O(N__27253),
            .I(N__27241));
    InMux I__4815 (
            .O(N__27252),
            .I(N__27241));
    Odrv4 I__4814 (
            .O(N__27249),
            .I(data_in_1_6));
    LocalMux I__4813 (
            .O(N__27246),
            .I(data_in_1_6));
    LocalMux I__4812 (
            .O(N__27241),
            .I(data_in_1_6));
    InMux I__4811 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4810 (
            .O(N__27231),
            .I(N__27228));
    Span4Mux_h I__4809 (
            .O(N__27228),
            .I(N__27225));
    Span4Mux_h I__4808 (
            .O(N__27225),
            .I(N__27222));
    Odrv4 I__4807 (
            .O(N__27222),
            .I(\c0.rx.n18304 ));
    InMux I__4806 (
            .O(N__27219),
            .I(N__27213));
    InMux I__4805 (
            .O(N__27218),
            .I(N__27206));
    InMux I__4804 (
            .O(N__27217),
            .I(N__27206));
    InMux I__4803 (
            .O(N__27216),
            .I(N__27202));
    LocalMux I__4802 (
            .O(N__27213),
            .I(N__27199));
    InMux I__4801 (
            .O(N__27212),
            .I(N__27194));
    InMux I__4800 (
            .O(N__27211),
            .I(N__27194));
    LocalMux I__4799 (
            .O(N__27206),
            .I(N__27191));
    CascadeMux I__4798 (
            .O(N__27205),
            .I(N__27188));
    LocalMux I__4797 (
            .O(N__27202),
            .I(N__27184));
    Span4Mux_h I__4796 (
            .O(N__27199),
            .I(N__27181));
    LocalMux I__4795 (
            .O(N__27194),
            .I(N__27178));
    Span4Mux_h I__4794 (
            .O(N__27191),
            .I(N__27175));
    InMux I__4793 (
            .O(N__27188),
            .I(N__27172));
    InMux I__4792 (
            .O(N__27187),
            .I(N__27169));
    Odrv4 I__4791 (
            .O(N__27184),
            .I(rx_data_5));
    Odrv4 I__4790 (
            .O(N__27181),
            .I(rx_data_5));
    Odrv12 I__4789 (
            .O(N__27178),
            .I(rx_data_5));
    Odrv4 I__4788 (
            .O(N__27175),
            .I(rx_data_5));
    LocalMux I__4787 (
            .O(N__27172),
            .I(rx_data_5));
    LocalMux I__4786 (
            .O(N__27169),
            .I(rx_data_5));
    CascadeMux I__4785 (
            .O(N__27156),
            .I(N__27152));
    InMux I__4784 (
            .O(N__27155),
            .I(N__27145));
    InMux I__4783 (
            .O(N__27152),
            .I(N__27145));
    InMux I__4782 (
            .O(N__27151),
            .I(N__27140));
    InMux I__4781 (
            .O(N__27150),
            .I(N__27140));
    LocalMux I__4780 (
            .O(N__27145),
            .I(data_in_3_5));
    LocalMux I__4779 (
            .O(N__27140),
            .I(data_in_3_5));
    CascadeMux I__4778 (
            .O(N__27135),
            .I(N__27131));
    InMux I__4777 (
            .O(N__27134),
            .I(N__27128));
    InMux I__4776 (
            .O(N__27131),
            .I(N__27125));
    LocalMux I__4775 (
            .O(N__27128),
            .I(N__27122));
    LocalMux I__4774 (
            .O(N__27125),
            .I(N__27116));
    Span4Mux_v I__4773 (
            .O(N__27122),
            .I(N__27116));
    InMux I__4772 (
            .O(N__27121),
            .I(N__27113));
    Span4Mux_v I__4771 (
            .O(N__27116),
            .I(N__27107));
    LocalMux I__4770 (
            .O(N__27113),
            .I(N__27103));
    InMux I__4769 (
            .O(N__27112),
            .I(N__27100));
    InMux I__4768 (
            .O(N__27111),
            .I(N__27097));
    CascadeMux I__4767 (
            .O(N__27110),
            .I(N__27093));
    Span4Mux_h I__4766 (
            .O(N__27107),
            .I(N__27090));
    InMux I__4765 (
            .O(N__27106),
            .I(N__27087));
    Span4Mux_v I__4764 (
            .O(N__27103),
            .I(N__27080));
    LocalMux I__4763 (
            .O(N__27100),
            .I(N__27080));
    LocalMux I__4762 (
            .O(N__27097),
            .I(N__27080));
    InMux I__4761 (
            .O(N__27096),
            .I(N__27075));
    InMux I__4760 (
            .O(N__27093),
            .I(N__27075));
    Odrv4 I__4759 (
            .O(N__27090),
            .I(rx_data_1));
    LocalMux I__4758 (
            .O(N__27087),
            .I(rx_data_1));
    Odrv4 I__4757 (
            .O(N__27080),
            .I(rx_data_1));
    LocalMux I__4756 (
            .O(N__27075),
            .I(rx_data_1));
    InMux I__4755 (
            .O(N__27066),
            .I(N__27063));
    LocalMux I__4754 (
            .O(N__27063),
            .I(N__27057));
    InMux I__4753 (
            .O(N__27062),
            .I(N__27054));
    InMux I__4752 (
            .O(N__27061),
            .I(N__27051));
    InMux I__4751 (
            .O(N__27060),
            .I(N__27048));
    Odrv4 I__4750 (
            .O(N__27057),
            .I(data_in_3_0));
    LocalMux I__4749 (
            .O(N__27054),
            .I(data_in_3_0));
    LocalMux I__4748 (
            .O(N__27051),
            .I(data_in_3_0));
    LocalMux I__4747 (
            .O(N__27048),
            .I(data_in_3_0));
    InMux I__4746 (
            .O(N__27039),
            .I(N__27036));
    LocalMux I__4745 (
            .O(N__27036),
            .I(N__27032));
    CascadeMux I__4744 (
            .O(N__27035),
            .I(N__27027));
    Span4Mux_v I__4743 (
            .O(N__27032),
            .I(N__27024));
    InMux I__4742 (
            .O(N__27031),
            .I(N__27021));
    InMux I__4741 (
            .O(N__27030),
            .I(N__27016));
    InMux I__4740 (
            .O(N__27027),
            .I(N__27016));
    Odrv4 I__4739 (
            .O(N__27024),
            .I(data_in_2_0));
    LocalMux I__4738 (
            .O(N__27021),
            .I(data_in_2_0));
    LocalMux I__4737 (
            .O(N__27016),
            .I(data_in_2_0));
    InMux I__4736 (
            .O(N__27009),
            .I(N__27005));
    CascadeMux I__4735 (
            .O(N__27008),
            .I(N__27002));
    LocalMux I__4734 (
            .O(N__27005),
            .I(N__26997));
    InMux I__4733 (
            .O(N__27002),
            .I(N__26992));
    InMux I__4732 (
            .O(N__27001),
            .I(N__26992));
    InMux I__4731 (
            .O(N__27000),
            .I(N__26989));
    Odrv4 I__4730 (
            .O(N__26997),
            .I(data_in_1_7));
    LocalMux I__4729 (
            .O(N__26992),
            .I(data_in_1_7));
    LocalMux I__4728 (
            .O(N__26989),
            .I(data_in_1_7));
    InMux I__4727 (
            .O(N__26982),
            .I(N__26979));
    LocalMux I__4726 (
            .O(N__26979),
            .I(\c0.n13693 ));
    InMux I__4725 (
            .O(N__26976),
            .I(N__26971));
    InMux I__4724 (
            .O(N__26975),
            .I(N__26968));
    InMux I__4723 (
            .O(N__26974),
            .I(N__26964));
    LocalMux I__4722 (
            .O(N__26971),
            .I(N__26959));
    LocalMux I__4721 (
            .O(N__26968),
            .I(N__26959));
    InMux I__4720 (
            .O(N__26967),
            .I(N__26951));
    LocalMux I__4719 (
            .O(N__26964),
            .I(N__26946));
    Span4Mux_h I__4718 (
            .O(N__26959),
            .I(N__26946));
    InMux I__4717 (
            .O(N__26958),
            .I(N__26943));
    InMux I__4716 (
            .O(N__26957),
            .I(N__26938));
    InMux I__4715 (
            .O(N__26956),
            .I(N__26938));
    InMux I__4714 (
            .O(N__26955),
            .I(N__26933));
    InMux I__4713 (
            .O(N__26954),
            .I(N__26933));
    LocalMux I__4712 (
            .O(N__26951),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    Odrv4 I__4711 (
            .O(N__26946),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    LocalMux I__4710 (
            .O(N__26943),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    LocalMux I__4709 (
            .O(N__26938),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    LocalMux I__4708 (
            .O(N__26933),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    CascadeMux I__4707 (
            .O(N__26922),
            .I(\c0.rx.n11041_cascade_ ));
    InMux I__4706 (
            .O(N__26919),
            .I(N__26916));
    LocalMux I__4705 (
            .O(N__26916),
            .I(N__26913));
    Odrv4 I__4704 (
            .O(N__26913),
            .I(\c0.n8_adj_2385 ));
    InMux I__4703 (
            .O(N__26910),
            .I(N__26907));
    LocalMux I__4702 (
            .O(N__26907),
            .I(\c0.n15_adj_2372 ));
    InMux I__4701 (
            .O(N__26904),
            .I(N__26896));
    InMux I__4700 (
            .O(N__26903),
            .I(N__26896));
    InMux I__4699 (
            .O(N__26902),
            .I(N__26891));
    InMux I__4698 (
            .O(N__26901),
            .I(N__26891));
    LocalMux I__4697 (
            .O(N__26896),
            .I(data_in_1_2));
    LocalMux I__4696 (
            .O(N__26891),
            .I(data_in_1_2));
    CascadeMux I__4695 (
            .O(N__26886),
            .I(N__26882));
    InMux I__4694 (
            .O(N__26885),
            .I(N__26879));
    InMux I__4693 (
            .O(N__26882),
            .I(N__26876));
    LocalMux I__4692 (
            .O(N__26879),
            .I(data_in_0_7));
    LocalMux I__4691 (
            .O(N__26876),
            .I(data_in_0_7));
    InMux I__4690 (
            .O(N__26871),
            .I(N__26867));
    InMux I__4689 (
            .O(N__26870),
            .I(N__26860));
    LocalMux I__4688 (
            .O(N__26867),
            .I(N__26857));
    InMux I__4687 (
            .O(N__26866),
            .I(N__26852));
    InMux I__4686 (
            .O(N__26865),
            .I(N__26852));
    InMux I__4685 (
            .O(N__26864),
            .I(N__26848));
    InMux I__4684 (
            .O(N__26863),
            .I(N__26845));
    LocalMux I__4683 (
            .O(N__26860),
            .I(N__26842));
    Span4Mux_v I__4682 (
            .O(N__26857),
            .I(N__26837));
    LocalMux I__4681 (
            .O(N__26852),
            .I(N__26837));
    InMux I__4680 (
            .O(N__26851),
            .I(N__26834));
    LocalMux I__4679 (
            .O(N__26848),
            .I(\c0.rx.r_Bit_Index_0 ));
    LocalMux I__4678 (
            .O(N__26845),
            .I(\c0.rx.r_Bit_Index_0 ));
    Odrv4 I__4677 (
            .O(N__26842),
            .I(\c0.rx.r_Bit_Index_0 ));
    Odrv4 I__4676 (
            .O(N__26837),
            .I(\c0.rx.r_Bit_Index_0 ));
    LocalMux I__4675 (
            .O(N__26834),
            .I(\c0.rx.r_Bit_Index_0 ));
    InMux I__4674 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__4673 (
            .O(N__26820),
            .I(N__26817));
    Span12Mux_s9_v I__4672 (
            .O(N__26817),
            .I(N__26814));
    Odrv12 I__4671 (
            .O(N__26814),
            .I(n151));
    CascadeMux I__4670 (
            .O(N__26811),
            .I(n151_cascade_));
    CascadeMux I__4669 (
            .O(N__26808),
            .I(N__26804));
    InMux I__4668 (
            .O(N__26807),
            .I(N__26799));
    InMux I__4667 (
            .O(N__26804),
            .I(N__26796));
    InMux I__4666 (
            .O(N__26803),
            .I(N__26793));
    InMux I__4665 (
            .O(N__26802),
            .I(N__26790));
    LocalMux I__4664 (
            .O(N__26799),
            .I(N__26783));
    LocalMux I__4663 (
            .O(N__26796),
            .I(N__26783));
    LocalMux I__4662 (
            .O(N__26793),
            .I(N__26783));
    LocalMux I__4661 (
            .O(N__26790),
            .I(data_in_2_2));
    Odrv4 I__4660 (
            .O(N__26783),
            .I(data_in_2_2));
    InMux I__4659 (
            .O(N__26778),
            .I(N__26775));
    LocalMux I__4658 (
            .O(N__26775),
            .I(\c0.n18008 ));
    CascadeMux I__4657 (
            .O(N__26772),
            .I(\c0.n8_adj_2369_cascade_ ));
    InMux I__4656 (
            .O(N__26769),
            .I(N__26765));
    InMux I__4655 (
            .O(N__26768),
            .I(N__26762));
    LocalMux I__4654 (
            .O(N__26765),
            .I(\c0.n10493 ));
    LocalMux I__4653 (
            .O(N__26762),
            .I(\c0.n10493 ));
    InMux I__4652 (
            .O(N__26757),
            .I(N__26754));
    LocalMux I__4651 (
            .O(N__26754),
            .I(N__26751));
    Span4Mux_v I__4650 (
            .O(N__26751),
            .I(N__26746));
    InMux I__4649 (
            .O(N__26750),
            .I(N__26743));
    InMux I__4648 (
            .O(N__26749),
            .I(N__26740));
    Odrv4 I__4647 (
            .O(N__26746),
            .I(data_in_1_0));
    LocalMux I__4646 (
            .O(N__26743),
            .I(data_in_1_0));
    LocalMux I__4645 (
            .O(N__26740),
            .I(data_in_1_0));
    InMux I__4644 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__4643 (
            .O(N__26730),
            .I(\c0.rx.n110 ));
    CascadeMux I__4642 (
            .O(N__26727),
            .I(N__26722));
    CascadeMux I__4641 (
            .O(N__26726),
            .I(N__26719));
    InMux I__4640 (
            .O(N__26725),
            .I(N__26715));
    InMux I__4639 (
            .O(N__26722),
            .I(N__26712));
    InMux I__4638 (
            .O(N__26719),
            .I(N__26709));
    InMux I__4637 (
            .O(N__26718),
            .I(N__26706));
    LocalMux I__4636 (
            .O(N__26715),
            .I(N__26700));
    LocalMux I__4635 (
            .O(N__26712),
            .I(N__26693));
    LocalMux I__4634 (
            .O(N__26709),
            .I(N__26693));
    LocalMux I__4633 (
            .O(N__26706),
            .I(N__26693));
    InMux I__4632 (
            .O(N__26705),
            .I(N__26690));
    InMux I__4631 (
            .O(N__26704),
            .I(N__26684));
    InMux I__4630 (
            .O(N__26703),
            .I(N__26684));
    Sp12to4 I__4629 (
            .O(N__26700),
            .I(N__26681));
    Span4Mux_v I__4628 (
            .O(N__26693),
            .I(N__26676));
    LocalMux I__4627 (
            .O(N__26690),
            .I(N__26676));
    InMux I__4626 (
            .O(N__26689),
            .I(N__26673));
    LocalMux I__4625 (
            .O(N__26684),
            .I(rx_data_2));
    Odrv12 I__4624 (
            .O(N__26681),
            .I(rx_data_2));
    Odrv4 I__4623 (
            .O(N__26676),
            .I(rx_data_2));
    LocalMux I__4622 (
            .O(N__26673),
            .I(rx_data_2));
    CascadeMux I__4621 (
            .O(N__26664),
            .I(\c0.rx.r_SM_Main_2_N_2088_2_cascade_ ));
    InMux I__4620 (
            .O(N__26661),
            .I(N__26656));
    InMux I__4619 (
            .O(N__26660),
            .I(N__26651));
    InMux I__4618 (
            .O(N__26659),
            .I(N__26651));
    LocalMux I__4617 (
            .O(N__26656),
            .I(\c0.rx.n161 ));
    LocalMux I__4616 (
            .O(N__26651),
            .I(\c0.rx.n161 ));
    CascadeMux I__4615 (
            .O(N__26646),
            .I(N__26643));
    InMux I__4614 (
            .O(N__26643),
            .I(N__26639));
    CascadeMux I__4613 (
            .O(N__26642),
            .I(N__26634));
    LocalMux I__4612 (
            .O(N__26639),
            .I(N__26630));
    InMux I__4611 (
            .O(N__26638),
            .I(N__26625));
    InMux I__4610 (
            .O(N__26637),
            .I(N__26621));
    InMux I__4609 (
            .O(N__26634),
            .I(N__26616));
    InMux I__4608 (
            .O(N__26633),
            .I(N__26616));
    Span4Mux_h I__4607 (
            .O(N__26630),
            .I(N__26613));
    InMux I__4606 (
            .O(N__26629),
            .I(N__26610));
    InMux I__4605 (
            .O(N__26628),
            .I(N__26607));
    LocalMux I__4604 (
            .O(N__26625),
            .I(N__26604));
    InMux I__4603 (
            .O(N__26624),
            .I(N__26601));
    LocalMux I__4602 (
            .O(N__26621),
            .I(N__26598));
    LocalMux I__4601 (
            .O(N__26616),
            .I(N__26595));
    Sp12to4 I__4600 (
            .O(N__26613),
            .I(N__26592));
    LocalMux I__4599 (
            .O(N__26610),
            .I(N__26585));
    LocalMux I__4598 (
            .O(N__26607),
            .I(N__26585));
    Span4Mux_v I__4597 (
            .O(N__26604),
            .I(N__26585));
    LocalMux I__4596 (
            .O(N__26601),
            .I(rx_data_0));
    Odrv4 I__4595 (
            .O(N__26598),
            .I(rx_data_0));
    Odrv4 I__4594 (
            .O(N__26595),
            .I(rx_data_0));
    Odrv12 I__4593 (
            .O(N__26592),
            .I(rx_data_0));
    Odrv4 I__4592 (
            .O(N__26585),
            .I(rx_data_0));
    CascadeMux I__4591 (
            .O(N__26574),
            .I(N__26568));
    InMux I__4590 (
            .O(N__26573),
            .I(N__26563));
    InMux I__4589 (
            .O(N__26572),
            .I(N__26563));
    InMux I__4588 (
            .O(N__26571),
            .I(N__26560));
    InMux I__4587 (
            .O(N__26568),
            .I(N__26557));
    LocalMux I__4586 (
            .O(N__26563),
            .I(data_in_3_2));
    LocalMux I__4585 (
            .O(N__26560),
            .I(data_in_3_2));
    LocalMux I__4584 (
            .O(N__26557),
            .I(data_in_3_2));
    InMux I__4583 (
            .O(N__26550),
            .I(N__26546));
    InMux I__4582 (
            .O(N__26549),
            .I(N__26542));
    LocalMux I__4581 (
            .O(N__26546),
            .I(N__26539));
    InMux I__4580 (
            .O(N__26545),
            .I(N__26536));
    LocalMux I__4579 (
            .O(N__26542),
            .I(data_in_0_6));
    Odrv4 I__4578 (
            .O(N__26539),
            .I(data_in_0_6));
    LocalMux I__4577 (
            .O(N__26536),
            .I(data_in_0_6));
    CascadeMux I__4576 (
            .O(N__26529),
            .I(N__26524));
    InMux I__4575 (
            .O(N__26528),
            .I(N__26520));
    InMux I__4574 (
            .O(N__26527),
            .I(N__26515));
    InMux I__4573 (
            .O(N__26524),
            .I(N__26515));
    InMux I__4572 (
            .O(N__26523),
            .I(N__26512));
    LocalMux I__4571 (
            .O(N__26520),
            .I(data_in_3_6));
    LocalMux I__4570 (
            .O(N__26515),
            .I(data_in_3_6));
    LocalMux I__4569 (
            .O(N__26512),
            .I(data_in_3_6));
    CascadeMux I__4568 (
            .O(N__26505),
            .I(N__26502));
    InMux I__4567 (
            .O(N__26502),
            .I(N__26497));
    InMux I__4566 (
            .O(N__26501),
            .I(N__26491));
    InMux I__4565 (
            .O(N__26500),
            .I(N__26488));
    LocalMux I__4564 (
            .O(N__26497),
            .I(N__26485));
    InMux I__4563 (
            .O(N__26496),
            .I(N__26482));
    InMux I__4562 (
            .O(N__26495),
            .I(N__26479));
    CascadeMux I__4561 (
            .O(N__26494),
            .I(N__26476));
    LocalMux I__4560 (
            .O(N__26491),
            .I(N__26471));
    LocalMux I__4559 (
            .O(N__26488),
            .I(N__26468));
    Span4Mux_v I__4558 (
            .O(N__26485),
            .I(N__26465));
    LocalMux I__4557 (
            .O(N__26482),
            .I(N__26460));
    LocalMux I__4556 (
            .O(N__26479),
            .I(N__26460));
    InMux I__4555 (
            .O(N__26476),
            .I(N__26455));
    InMux I__4554 (
            .O(N__26475),
            .I(N__26455));
    CascadeMux I__4553 (
            .O(N__26474),
            .I(N__26452));
    Span4Mux_v I__4552 (
            .O(N__26471),
            .I(N__26449));
    Span4Mux_h I__4551 (
            .O(N__26468),
            .I(N__26446));
    Sp12to4 I__4550 (
            .O(N__26465),
            .I(N__26439));
    Span12Mux_v I__4549 (
            .O(N__26460),
            .I(N__26439));
    LocalMux I__4548 (
            .O(N__26455),
            .I(N__26439));
    InMux I__4547 (
            .O(N__26452),
            .I(N__26436));
    Odrv4 I__4546 (
            .O(N__26449),
            .I(rx_data_4));
    Odrv4 I__4545 (
            .O(N__26446),
            .I(rx_data_4));
    Odrv12 I__4544 (
            .O(N__26439),
            .I(rx_data_4));
    LocalMux I__4543 (
            .O(N__26436),
            .I(rx_data_4));
    InMux I__4542 (
            .O(N__26427),
            .I(N__26416));
    InMux I__4541 (
            .O(N__26426),
            .I(N__26416));
    InMux I__4540 (
            .O(N__26425),
            .I(N__26413));
    InMux I__4539 (
            .O(N__26424),
            .I(N__26410));
    InMux I__4538 (
            .O(N__26423),
            .I(N__26403));
    InMux I__4537 (
            .O(N__26422),
            .I(N__26403));
    InMux I__4536 (
            .O(N__26421),
            .I(N__26403));
    LocalMux I__4535 (
            .O(N__26416),
            .I(n120));
    LocalMux I__4534 (
            .O(N__26413),
            .I(n120));
    LocalMux I__4533 (
            .O(N__26410),
            .I(n120));
    LocalMux I__4532 (
            .O(N__26403),
            .I(n120));
    InMux I__4531 (
            .O(N__26394),
            .I(N__26390));
    CascadeMux I__4530 (
            .O(N__26393),
            .I(N__26386));
    LocalMux I__4529 (
            .O(N__26390),
            .I(N__26383));
    InMux I__4528 (
            .O(N__26389),
            .I(N__26378));
    InMux I__4527 (
            .O(N__26386),
            .I(N__26378));
    Odrv12 I__4526 (
            .O(N__26383),
            .I(data_in_frame_2_4));
    LocalMux I__4525 (
            .O(N__26378),
            .I(data_in_frame_2_4));
    CascadeMux I__4524 (
            .O(N__26373),
            .I(\c0.rx.n18729_cascade_ ));
    CascadeMux I__4523 (
            .O(N__26370),
            .I(\c0.rx.n18732_cascade_ ));
    InMux I__4522 (
            .O(N__26367),
            .I(N__26364));
    LocalMux I__4521 (
            .O(N__26364),
            .I(N__26361));
    Odrv4 I__4520 (
            .O(N__26361),
            .I(\c0.rx.n11 ));
    InMux I__4519 (
            .O(N__26358),
            .I(N__26355));
    LocalMux I__4518 (
            .O(N__26355),
            .I(N__26351));
    InMux I__4517 (
            .O(N__26354),
            .I(N__26348));
    Odrv4 I__4516 (
            .O(N__26351),
            .I(n12582));
    LocalMux I__4515 (
            .O(N__26348),
            .I(n12582));
    InMux I__4514 (
            .O(N__26343),
            .I(N__26340));
    LocalMux I__4513 (
            .O(N__26340),
            .I(N__26336));
    InMux I__4512 (
            .O(N__26339),
            .I(N__26333));
    Span4Mux_h I__4511 (
            .O(N__26336),
            .I(N__26328));
    LocalMux I__4510 (
            .O(N__26333),
            .I(N__26328));
    Odrv4 I__4509 (
            .O(N__26328),
            .I(n135_adj_2463));
    CascadeMux I__4508 (
            .O(N__26325),
            .I(n4_adj_2471_cascade_));
    InMux I__4507 (
            .O(N__26322),
            .I(N__26318));
    InMux I__4506 (
            .O(N__26321),
            .I(N__26315));
    LocalMux I__4505 (
            .O(N__26318),
            .I(N__26312));
    LocalMux I__4504 (
            .O(N__26315),
            .I(data_in_frame_5_5));
    Odrv4 I__4503 (
            .O(N__26312),
            .I(data_in_frame_5_5));
    InMux I__4502 (
            .O(N__26307),
            .I(N__26304));
    LocalMux I__4501 (
            .O(N__26304),
            .I(N__26299));
    InMux I__4500 (
            .O(N__26303),
            .I(N__26294));
    InMux I__4499 (
            .O(N__26302),
            .I(N__26291));
    Span4Mux_h I__4498 (
            .O(N__26299),
            .I(N__26288));
    InMux I__4497 (
            .O(N__26298),
            .I(N__26285));
    InMux I__4496 (
            .O(N__26297),
            .I(N__26282));
    LocalMux I__4495 (
            .O(N__26294),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__4494 (
            .O(N__26291),
            .I(\c0.data_in_frame_1_3 ));
    Odrv4 I__4493 (
            .O(N__26288),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__4492 (
            .O(N__26285),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__4491 (
            .O(N__26282),
            .I(\c0.data_in_frame_1_3 ));
    CascadeMux I__4490 (
            .O(N__26271),
            .I(\c0.n16981_cascade_ ));
    InMux I__4489 (
            .O(N__26268),
            .I(N__26265));
    LocalMux I__4488 (
            .O(N__26265),
            .I(\c0.n20_adj_2397 ));
    InMux I__4487 (
            .O(N__26262),
            .I(N__26259));
    LocalMux I__4486 (
            .O(N__26259),
            .I(N__26256));
    Span4Mux_v I__4485 (
            .O(N__26256),
            .I(N__26253));
    Span4Mux_h I__4484 (
            .O(N__26253),
            .I(N__26250));
    Odrv4 I__4483 (
            .O(N__26250),
            .I(\c0.n20_adj_2350 ));
    InMux I__4482 (
            .O(N__26247),
            .I(N__26244));
    LocalMux I__4481 (
            .O(N__26244),
            .I(\c0.n2128 ));
    InMux I__4480 (
            .O(N__26241),
            .I(N__26237));
    InMux I__4479 (
            .O(N__26240),
            .I(N__26234));
    LocalMux I__4478 (
            .O(N__26237),
            .I(N__26231));
    LocalMux I__4477 (
            .O(N__26234),
            .I(data_in_frame_6_4));
    Odrv4 I__4476 (
            .O(N__26231),
            .I(data_in_frame_6_4));
    InMux I__4475 (
            .O(N__26226),
            .I(N__26223));
    LocalMux I__4474 (
            .O(N__26223),
            .I(N__26219));
    InMux I__4473 (
            .O(N__26222),
            .I(N__26216));
    Span4Mux_h I__4472 (
            .O(N__26219),
            .I(N__26213));
    LocalMux I__4471 (
            .O(N__26216),
            .I(data_in_frame_5_0));
    Odrv4 I__4470 (
            .O(N__26213),
            .I(data_in_frame_5_0));
    CascadeMux I__4469 (
            .O(N__26208),
            .I(\c0.n2128_cascade_ ));
    InMux I__4468 (
            .O(N__26205),
            .I(N__26202));
    LocalMux I__4467 (
            .O(N__26202),
            .I(N__26199));
    Odrv4 I__4466 (
            .O(N__26199),
            .I(\c0.n22_adj_2392 ));
    InMux I__4465 (
            .O(N__26196),
            .I(N__26193));
    LocalMux I__4464 (
            .O(N__26193),
            .I(N__26188));
    InMux I__4463 (
            .O(N__26192),
            .I(N__26185));
    InMux I__4462 (
            .O(N__26191),
            .I(N__26182));
    Odrv4 I__4461 (
            .O(N__26188),
            .I(data_in_frame_0_2));
    LocalMux I__4460 (
            .O(N__26185),
            .I(data_in_frame_0_2));
    LocalMux I__4459 (
            .O(N__26182),
            .I(data_in_frame_0_2));
    InMux I__4458 (
            .O(N__26175),
            .I(N__26171));
    CascadeMux I__4457 (
            .O(N__26174),
            .I(N__26167));
    LocalMux I__4456 (
            .O(N__26171),
            .I(N__26164));
    InMux I__4455 (
            .O(N__26170),
            .I(N__26160));
    InMux I__4454 (
            .O(N__26167),
            .I(N__26157));
    Span4Mux_v I__4453 (
            .O(N__26164),
            .I(N__26154));
    InMux I__4452 (
            .O(N__26163),
            .I(N__26151));
    LocalMux I__4451 (
            .O(N__26160),
            .I(data_in_frame_0_3));
    LocalMux I__4450 (
            .O(N__26157),
            .I(data_in_frame_0_3));
    Odrv4 I__4449 (
            .O(N__26154),
            .I(data_in_frame_0_3));
    LocalMux I__4448 (
            .O(N__26151),
            .I(data_in_frame_0_3));
    InMux I__4447 (
            .O(N__26142),
            .I(N__26136));
    InMux I__4446 (
            .O(N__26141),
            .I(N__26136));
    LocalMux I__4445 (
            .O(N__26136),
            .I(\c0.n2120 ));
    InMux I__4444 (
            .O(N__26133),
            .I(N__26128));
    InMux I__4443 (
            .O(N__26132),
            .I(N__26125));
    InMux I__4442 (
            .O(N__26131),
            .I(N__26122));
    LocalMux I__4441 (
            .O(N__26128),
            .I(N__26119));
    LocalMux I__4440 (
            .O(N__26125),
            .I(\c0.n2124 ));
    LocalMux I__4439 (
            .O(N__26122),
            .I(\c0.n2124 ));
    Odrv4 I__4438 (
            .O(N__26119),
            .I(\c0.n2124 ));
    InMux I__4437 (
            .O(N__26112),
            .I(N__26108));
    InMux I__4436 (
            .O(N__26111),
            .I(N__26105));
    LocalMux I__4435 (
            .O(N__26108),
            .I(N__26102));
    LocalMux I__4434 (
            .O(N__26105),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__4433 (
            .O(N__26102),
            .I(\c0.data_in_frame_3_4 ));
    CascadeMux I__4432 (
            .O(N__26097),
            .I(\c0.n2120_cascade_ ));
    InMux I__4431 (
            .O(N__26094),
            .I(N__26090));
    InMux I__4430 (
            .O(N__26093),
            .I(N__26087));
    LocalMux I__4429 (
            .O(N__26090),
            .I(N__26084));
    LocalMux I__4428 (
            .O(N__26087),
            .I(\c0.data_in_frame_3_6 ));
    Odrv4 I__4427 (
            .O(N__26084),
            .I(\c0.data_in_frame_3_6 ));
    InMux I__4426 (
            .O(N__26079),
            .I(N__26076));
    LocalMux I__4425 (
            .O(N__26076),
            .I(N__26073));
    Odrv4 I__4424 (
            .O(N__26073),
            .I(\c0.n19_adj_2415 ));
    InMux I__4423 (
            .O(N__26070),
            .I(N__26063));
    InMux I__4422 (
            .O(N__26069),
            .I(N__26060));
    InMux I__4421 (
            .O(N__26068),
            .I(N__26057));
    InMux I__4420 (
            .O(N__26067),
            .I(N__26052));
    InMux I__4419 (
            .O(N__26066),
            .I(N__26052));
    LocalMux I__4418 (
            .O(N__26063),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__4417 (
            .O(N__26060),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__4416 (
            .O(N__26057),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__4415 (
            .O(N__26052),
            .I(\c0.data_in_frame_1_0 ));
    InMux I__4414 (
            .O(N__26043),
            .I(N__26039));
    InMux I__4413 (
            .O(N__26042),
            .I(N__26033));
    LocalMux I__4412 (
            .O(N__26039),
            .I(N__26030));
    InMux I__4411 (
            .O(N__26038),
            .I(N__26025));
    InMux I__4410 (
            .O(N__26037),
            .I(N__26025));
    InMux I__4409 (
            .O(N__26036),
            .I(N__26022));
    LocalMux I__4408 (
            .O(N__26033),
            .I(\c0.data_in_frame_1_1 ));
    Odrv4 I__4407 (
            .O(N__26030),
            .I(\c0.data_in_frame_1_1 ));
    LocalMux I__4406 (
            .O(N__26025),
            .I(\c0.data_in_frame_1_1 ));
    LocalMux I__4405 (
            .O(N__26022),
            .I(\c0.data_in_frame_1_1 ));
    InMux I__4404 (
            .O(N__26013),
            .I(N__26009));
    InMux I__4403 (
            .O(N__26012),
            .I(N__26005));
    LocalMux I__4402 (
            .O(N__26009),
            .I(N__25999));
    InMux I__4401 (
            .O(N__26008),
            .I(N__25995));
    LocalMux I__4400 (
            .O(N__26005),
            .I(N__25991));
    InMux I__4399 (
            .O(N__26004),
            .I(N__25986));
    InMux I__4398 (
            .O(N__26003),
            .I(N__25986));
    InMux I__4397 (
            .O(N__26002),
            .I(N__25983));
    Span4Mux_h I__4396 (
            .O(N__25999),
            .I(N__25980));
    InMux I__4395 (
            .O(N__25998),
            .I(N__25977));
    LocalMux I__4394 (
            .O(N__25995),
            .I(N__25974));
    InMux I__4393 (
            .O(N__25994),
            .I(N__25971));
    Span4Mux_v I__4392 (
            .O(N__25991),
            .I(N__25966));
    LocalMux I__4391 (
            .O(N__25986),
            .I(N__25966));
    LocalMux I__4390 (
            .O(N__25983),
            .I(data_in_frame_0_7));
    Odrv4 I__4389 (
            .O(N__25980),
            .I(data_in_frame_0_7));
    LocalMux I__4388 (
            .O(N__25977),
            .I(data_in_frame_0_7));
    Odrv4 I__4387 (
            .O(N__25974),
            .I(data_in_frame_0_7));
    LocalMux I__4386 (
            .O(N__25971),
            .I(data_in_frame_0_7));
    Odrv4 I__4385 (
            .O(N__25966),
            .I(data_in_frame_0_7));
    InMux I__4384 (
            .O(N__25953),
            .I(N__25949));
    InMux I__4383 (
            .O(N__25952),
            .I(N__25946));
    LocalMux I__4382 (
            .O(N__25949),
            .I(N__25941));
    LocalMux I__4381 (
            .O(N__25946),
            .I(N__25937));
    InMux I__4380 (
            .O(N__25945),
            .I(N__25932));
    InMux I__4379 (
            .O(N__25944),
            .I(N__25932));
    Span4Mux_h I__4378 (
            .O(N__25941),
            .I(N__25929));
    InMux I__4377 (
            .O(N__25940),
            .I(N__25926));
    Odrv4 I__4376 (
            .O(N__25937),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__4375 (
            .O(N__25932),
            .I(\c0.data_in_frame_1_4 ));
    Odrv4 I__4374 (
            .O(N__25929),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__4373 (
            .O(N__25926),
            .I(\c0.data_in_frame_1_4 ));
    CascadeMux I__4372 (
            .O(N__25917),
            .I(\c0.n17721_cascade_ ));
    InMux I__4371 (
            .O(N__25914),
            .I(N__25910));
    InMux I__4370 (
            .O(N__25913),
            .I(N__25906));
    LocalMux I__4369 (
            .O(N__25910),
            .I(N__25903));
    InMux I__4368 (
            .O(N__25909),
            .I(N__25897));
    LocalMux I__4367 (
            .O(N__25906),
            .I(N__25894));
    Span4Mux_h I__4366 (
            .O(N__25903),
            .I(N__25891));
    InMux I__4365 (
            .O(N__25902),
            .I(N__25888));
    InMux I__4364 (
            .O(N__25901),
            .I(N__25883));
    InMux I__4363 (
            .O(N__25900),
            .I(N__25883));
    LocalMux I__4362 (
            .O(N__25897),
            .I(data_in_frame_0_6));
    Odrv4 I__4361 (
            .O(N__25894),
            .I(data_in_frame_0_6));
    Odrv4 I__4360 (
            .O(N__25891),
            .I(data_in_frame_0_6));
    LocalMux I__4359 (
            .O(N__25888),
            .I(data_in_frame_0_6));
    LocalMux I__4358 (
            .O(N__25883),
            .I(data_in_frame_0_6));
    InMux I__4357 (
            .O(N__25872),
            .I(N__25869));
    LocalMux I__4356 (
            .O(N__25869),
            .I(\c0.n10_adj_2390 ));
    InMux I__4355 (
            .O(N__25866),
            .I(N__25855));
    InMux I__4354 (
            .O(N__25865),
            .I(N__25855));
    InMux I__4353 (
            .O(N__25864),
            .I(N__25852));
    InMux I__4352 (
            .O(N__25863),
            .I(N__25849));
    InMux I__4351 (
            .O(N__25862),
            .I(N__25846));
    InMux I__4350 (
            .O(N__25861),
            .I(N__25841));
    InMux I__4349 (
            .O(N__25860),
            .I(N__25841));
    LocalMux I__4348 (
            .O(N__25855),
            .I(n16797));
    LocalMux I__4347 (
            .O(N__25852),
            .I(n16797));
    LocalMux I__4346 (
            .O(N__25849),
            .I(n16797));
    LocalMux I__4345 (
            .O(N__25846),
            .I(n16797));
    LocalMux I__4344 (
            .O(N__25841),
            .I(n16797));
    InMux I__4343 (
            .O(N__25830),
            .I(N__25827));
    LocalMux I__4342 (
            .O(N__25827),
            .I(N__25823));
    InMux I__4341 (
            .O(N__25826),
            .I(N__25820));
    Span4Mux_h I__4340 (
            .O(N__25823),
            .I(N__25817));
    LocalMux I__4339 (
            .O(N__25820),
            .I(data_in_frame_5_4));
    Odrv4 I__4338 (
            .O(N__25817),
            .I(data_in_frame_5_4));
    InMux I__4337 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__4336 (
            .O(N__25809),
            .I(n158));
    InMux I__4335 (
            .O(N__25806),
            .I(N__25803));
    LocalMux I__4334 (
            .O(N__25803),
            .I(N__25799));
    InMux I__4333 (
            .O(N__25802),
            .I(N__25796));
    Span4Mux_h I__4332 (
            .O(N__25799),
            .I(N__25793));
    LocalMux I__4331 (
            .O(N__25796),
            .I(N__25790));
    Odrv4 I__4330 (
            .O(N__25793),
            .I(n12600));
    Odrv4 I__4329 (
            .O(N__25790),
            .I(n12600));
    CascadeMux I__4328 (
            .O(N__25785),
            .I(N__25776));
    InMux I__4327 (
            .O(N__25784),
            .I(N__25773));
    InMux I__4326 (
            .O(N__25783),
            .I(N__25770));
    CascadeMux I__4325 (
            .O(N__25782),
            .I(N__25767));
    CascadeMux I__4324 (
            .O(N__25781),
            .I(N__25764));
    InMux I__4323 (
            .O(N__25780),
            .I(N__25758));
    InMux I__4322 (
            .O(N__25779),
            .I(N__25758));
    InMux I__4321 (
            .O(N__25776),
            .I(N__25755));
    LocalMux I__4320 (
            .O(N__25773),
            .I(N__25752));
    LocalMux I__4319 (
            .O(N__25770),
            .I(N__25749));
    InMux I__4318 (
            .O(N__25767),
            .I(N__25746));
    InMux I__4317 (
            .O(N__25764),
            .I(N__25743));
    InMux I__4316 (
            .O(N__25763),
            .I(N__25740));
    LocalMux I__4315 (
            .O(N__25758),
            .I(N__25737));
    LocalMux I__4314 (
            .O(N__25755),
            .I(N__25734));
    Sp12to4 I__4313 (
            .O(N__25752),
            .I(N__25729));
    Sp12to4 I__4312 (
            .O(N__25749),
            .I(N__25729));
    LocalMux I__4311 (
            .O(N__25746),
            .I(rx_data_3));
    LocalMux I__4310 (
            .O(N__25743),
            .I(rx_data_3));
    LocalMux I__4309 (
            .O(N__25740),
            .I(rx_data_3));
    Odrv4 I__4308 (
            .O(N__25737),
            .I(rx_data_3));
    Odrv4 I__4307 (
            .O(N__25734),
            .I(rx_data_3));
    Odrv12 I__4306 (
            .O(N__25729),
            .I(rx_data_3));
    CascadeMux I__4305 (
            .O(N__25716),
            .I(N__25707));
    InMux I__4304 (
            .O(N__25715),
            .I(N__25689));
    InMux I__4303 (
            .O(N__25714),
            .I(N__25689));
    InMux I__4302 (
            .O(N__25713),
            .I(N__25689));
    InMux I__4301 (
            .O(N__25712),
            .I(N__25689));
    InMux I__4300 (
            .O(N__25711),
            .I(N__25689));
    InMux I__4299 (
            .O(N__25710),
            .I(N__25686));
    InMux I__4298 (
            .O(N__25707),
            .I(N__25679));
    InMux I__4297 (
            .O(N__25706),
            .I(N__25679));
    InMux I__4296 (
            .O(N__25705),
            .I(N__25679));
    CascadeMux I__4295 (
            .O(N__25704),
            .I(N__25674));
    InMux I__4294 (
            .O(N__25703),
            .I(N__25663));
    InMux I__4293 (
            .O(N__25702),
            .I(N__25663));
    InMux I__4292 (
            .O(N__25701),
            .I(N__25663));
    InMux I__4291 (
            .O(N__25700),
            .I(N__25660));
    LocalMux I__4290 (
            .O(N__25689),
            .I(N__25652));
    LocalMux I__4289 (
            .O(N__25686),
            .I(N__25652));
    LocalMux I__4288 (
            .O(N__25679),
            .I(N__25652));
    InMux I__4287 (
            .O(N__25678),
            .I(N__25649));
    InMux I__4286 (
            .O(N__25677),
            .I(N__25642));
    InMux I__4285 (
            .O(N__25674),
            .I(N__25642));
    InMux I__4284 (
            .O(N__25673),
            .I(N__25635));
    InMux I__4283 (
            .O(N__25672),
            .I(N__25635));
    InMux I__4282 (
            .O(N__25671),
            .I(N__25635));
    InMux I__4281 (
            .O(N__25670),
            .I(N__25632));
    LocalMux I__4280 (
            .O(N__25663),
            .I(N__25627));
    LocalMux I__4279 (
            .O(N__25660),
            .I(N__25627));
    InMux I__4278 (
            .O(N__25659),
            .I(N__25623));
    Span4Mux_v I__4277 (
            .O(N__25652),
            .I(N__25618));
    LocalMux I__4276 (
            .O(N__25649),
            .I(N__25618));
    InMux I__4275 (
            .O(N__25648),
            .I(N__25615));
    InMux I__4274 (
            .O(N__25647),
            .I(N__25612));
    LocalMux I__4273 (
            .O(N__25642),
            .I(N__25607));
    LocalMux I__4272 (
            .O(N__25635),
            .I(N__25607));
    LocalMux I__4271 (
            .O(N__25632),
            .I(N__25602));
    Span4Mux_v I__4270 (
            .O(N__25627),
            .I(N__25602));
    CascadeMux I__4269 (
            .O(N__25626),
            .I(N__25599));
    LocalMux I__4268 (
            .O(N__25623),
            .I(N__25587));
    Span4Mux_v I__4267 (
            .O(N__25618),
            .I(N__25587));
    LocalMux I__4266 (
            .O(N__25615),
            .I(N__25587));
    LocalMux I__4265 (
            .O(N__25612),
            .I(N__25587));
    Span12Mux_h I__4264 (
            .O(N__25607),
            .I(N__25584));
    Span4Mux_h I__4263 (
            .O(N__25602),
            .I(N__25581));
    InMux I__4262 (
            .O(N__25599),
            .I(N__25578));
    InMux I__4261 (
            .O(N__25598),
            .I(N__25571));
    InMux I__4260 (
            .O(N__25597),
            .I(N__25571));
    InMux I__4259 (
            .O(N__25596),
            .I(N__25571));
    Span4Mux_h I__4258 (
            .O(N__25587),
            .I(N__25568));
    Odrv12 I__4257 (
            .O(N__25584),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__4256 (
            .O(N__25581),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__4255 (
            .O(N__25578),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__4254 (
            .O(N__25571),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__4253 (
            .O(N__25568),
            .I(\c0.FRAME_MATCHER_i_1 ));
    InMux I__4252 (
            .O(N__25557),
            .I(N__25540));
    InMux I__4251 (
            .O(N__25556),
            .I(N__25533));
    InMux I__4250 (
            .O(N__25555),
            .I(N__25533));
    InMux I__4249 (
            .O(N__25554),
            .I(N__25533));
    InMux I__4248 (
            .O(N__25553),
            .I(N__25528));
    InMux I__4247 (
            .O(N__25552),
            .I(N__25528));
    InMux I__4246 (
            .O(N__25551),
            .I(N__25523));
    InMux I__4245 (
            .O(N__25550),
            .I(N__25523));
    InMux I__4244 (
            .O(N__25549),
            .I(N__25516));
    InMux I__4243 (
            .O(N__25548),
            .I(N__25516));
    InMux I__4242 (
            .O(N__25547),
            .I(N__25516));
    InMux I__4241 (
            .O(N__25546),
            .I(N__25507));
    InMux I__4240 (
            .O(N__25545),
            .I(N__25507));
    InMux I__4239 (
            .O(N__25544),
            .I(N__25507));
    InMux I__4238 (
            .O(N__25543),
            .I(N__25507));
    LocalMux I__4237 (
            .O(N__25540),
            .I(\c0.rx.n129 ));
    LocalMux I__4236 (
            .O(N__25533),
            .I(\c0.rx.n129 ));
    LocalMux I__4235 (
            .O(N__25528),
            .I(\c0.rx.n129 ));
    LocalMux I__4234 (
            .O(N__25523),
            .I(\c0.rx.n129 ));
    LocalMux I__4233 (
            .O(N__25516),
            .I(\c0.rx.n129 ));
    LocalMux I__4232 (
            .O(N__25507),
            .I(\c0.rx.n129 ));
    InMux I__4231 (
            .O(N__25494),
            .I(N__25490));
    InMux I__4230 (
            .O(N__25493),
            .I(N__25487));
    LocalMux I__4229 (
            .O(N__25490),
            .I(N__25484));
    LocalMux I__4228 (
            .O(N__25487),
            .I(data_in_frame_5_3));
    Odrv4 I__4227 (
            .O(N__25484),
            .I(data_in_frame_5_3));
    InMux I__4226 (
            .O(N__25479),
            .I(N__25472));
    CascadeMux I__4225 (
            .O(N__25478),
            .I(N__25469));
    InMux I__4224 (
            .O(N__25477),
            .I(N__25466));
    InMux I__4223 (
            .O(N__25476),
            .I(N__25463));
    InMux I__4222 (
            .O(N__25475),
            .I(N__25460));
    LocalMux I__4221 (
            .O(N__25472),
            .I(N__25457));
    InMux I__4220 (
            .O(N__25469),
            .I(N__25454));
    LocalMux I__4219 (
            .O(N__25466),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__4218 (
            .O(N__25463),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__4217 (
            .O(N__25460),
            .I(\c0.data_in_frame_1_2 ));
    Odrv4 I__4216 (
            .O(N__25457),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__4215 (
            .O(N__25454),
            .I(\c0.data_in_frame_1_2 ));
    InMux I__4214 (
            .O(N__25443),
            .I(N__25439));
    InMux I__4213 (
            .O(N__25442),
            .I(N__25436));
    LocalMux I__4212 (
            .O(N__25439),
            .I(N__25432));
    LocalMux I__4211 (
            .O(N__25436),
            .I(N__25429));
    InMux I__4210 (
            .O(N__25435),
            .I(N__25426));
    Span4Mux_h I__4209 (
            .O(N__25432),
            .I(N__25423));
    Odrv12 I__4208 (
            .O(N__25429),
            .I(\c0.n2122 ));
    LocalMux I__4207 (
            .O(N__25426),
            .I(\c0.n2122 ));
    Odrv4 I__4206 (
            .O(N__25423),
            .I(\c0.n2122 ));
    InMux I__4205 (
            .O(N__25416),
            .I(N__25412));
    CascadeMux I__4204 (
            .O(N__25415),
            .I(N__25409));
    LocalMux I__4203 (
            .O(N__25412),
            .I(N__25406));
    InMux I__4202 (
            .O(N__25409),
            .I(N__25403));
    Odrv4 I__4201 (
            .O(N__25406),
            .I(data_in_frame_6_5));
    LocalMux I__4200 (
            .O(N__25403),
            .I(data_in_frame_6_5));
    InMux I__4199 (
            .O(N__25398),
            .I(N__25395));
    LocalMux I__4198 (
            .O(N__25395),
            .I(\c0.n16994 ));
    InMux I__4197 (
            .O(N__25392),
            .I(N__25388));
    InMux I__4196 (
            .O(N__25391),
            .I(N__25385));
    LocalMux I__4195 (
            .O(N__25388),
            .I(N__25382));
    LocalMux I__4194 (
            .O(N__25385),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__4193 (
            .O(N__25382),
            .I(\c0.data_in_frame_3_2 ));
    CascadeMux I__4192 (
            .O(N__25377),
            .I(N__25374));
    InMux I__4191 (
            .O(N__25374),
            .I(N__25371));
    LocalMux I__4190 (
            .O(N__25371),
            .I(N__25367));
    InMux I__4189 (
            .O(N__25370),
            .I(N__25364));
    Span4Mux_h I__4188 (
            .O(N__25367),
            .I(N__25361));
    LocalMux I__4187 (
            .O(N__25364),
            .I(data_in_frame_6_6));
    Odrv4 I__4186 (
            .O(N__25361),
            .I(data_in_frame_6_6));
    InMux I__4185 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__4184 (
            .O(N__25353),
            .I(N__25350));
    Span4Mux_v I__4183 (
            .O(N__25350),
            .I(N__25346));
    InMux I__4182 (
            .O(N__25349),
            .I(N__25343));
    Span4Mux_v I__4181 (
            .O(N__25346),
            .I(N__25340));
    LocalMux I__4180 (
            .O(N__25343),
            .I(data_in_frame_5_1));
    Odrv4 I__4179 (
            .O(N__25340),
            .I(data_in_frame_5_1));
    InMux I__4178 (
            .O(N__25335),
            .I(N__25332));
    LocalMux I__4177 (
            .O(N__25332),
            .I(N__25328));
    InMux I__4176 (
            .O(N__25331),
            .I(N__25325));
    Span4Mux_h I__4175 (
            .O(N__25328),
            .I(N__25322));
    LocalMux I__4174 (
            .O(N__25325),
            .I(data_in_frame_6_2));
    Odrv4 I__4173 (
            .O(N__25322),
            .I(data_in_frame_6_2));
    InMux I__4172 (
            .O(N__25317),
            .I(N__25314));
    LocalMux I__4171 (
            .O(N__25314),
            .I(\c0.n18315 ));
    InMux I__4170 (
            .O(N__25311),
            .I(\c0.n16481 ));
    InMux I__4169 (
            .O(N__25308),
            .I(\c0.n16482 ));
    CascadeMux I__4168 (
            .O(N__25305),
            .I(N__25302));
    InMux I__4167 (
            .O(N__25302),
            .I(N__25296));
    InMux I__4166 (
            .O(N__25301),
            .I(N__25293));
    InMux I__4165 (
            .O(N__25300),
            .I(N__25288));
    InMux I__4164 (
            .O(N__25299),
            .I(N__25288));
    LocalMux I__4163 (
            .O(N__25296),
            .I(\c0.byte_transmit_counter2_5 ));
    LocalMux I__4162 (
            .O(N__25293),
            .I(\c0.byte_transmit_counter2_5 ));
    LocalMux I__4161 (
            .O(N__25288),
            .I(\c0.byte_transmit_counter2_5 ));
    InMux I__4160 (
            .O(N__25281),
            .I(N__25278));
    LocalMux I__4159 (
            .O(N__25278),
            .I(N__25275));
    Odrv4 I__4158 (
            .O(N__25275),
            .I(\c0.n18316 ));
    InMux I__4157 (
            .O(N__25272),
            .I(\c0.n16483 ));
    InMux I__4156 (
            .O(N__25269),
            .I(N__25264));
    InMux I__4155 (
            .O(N__25268),
            .I(N__25261));
    InMux I__4154 (
            .O(N__25267),
            .I(N__25257));
    LocalMux I__4153 (
            .O(N__25264),
            .I(N__25254));
    LocalMux I__4152 (
            .O(N__25261),
            .I(N__25251));
    InMux I__4151 (
            .O(N__25260),
            .I(N__25248));
    LocalMux I__4150 (
            .O(N__25257),
            .I(\c0.byte_transmit_counter2_6 ));
    Odrv12 I__4149 (
            .O(N__25254),
            .I(\c0.byte_transmit_counter2_6 ));
    Odrv4 I__4148 (
            .O(N__25251),
            .I(\c0.byte_transmit_counter2_6 ));
    LocalMux I__4147 (
            .O(N__25248),
            .I(\c0.byte_transmit_counter2_6 ));
    InMux I__4146 (
            .O(N__25239),
            .I(N__25236));
    LocalMux I__4145 (
            .O(N__25236),
            .I(N__25233));
    Odrv4 I__4144 (
            .O(N__25233),
            .I(\c0.n18317 ));
    InMux I__4143 (
            .O(N__25230),
            .I(\c0.n16484 ));
    InMux I__4142 (
            .O(N__25227),
            .I(N__25222));
    CascadeMux I__4141 (
            .O(N__25226),
            .I(N__25219));
    InMux I__4140 (
            .O(N__25225),
            .I(N__25215));
    LocalMux I__4139 (
            .O(N__25222),
            .I(N__25212));
    InMux I__4138 (
            .O(N__25219),
            .I(N__25207));
    InMux I__4137 (
            .O(N__25218),
            .I(N__25207));
    LocalMux I__4136 (
            .O(N__25215),
            .I(\c0.byte_transmit_counter2_7 ));
    Odrv4 I__4135 (
            .O(N__25212),
            .I(\c0.byte_transmit_counter2_7 ));
    LocalMux I__4134 (
            .O(N__25207),
            .I(\c0.byte_transmit_counter2_7 ));
    InMux I__4133 (
            .O(N__25200),
            .I(N__25185));
    InMux I__4132 (
            .O(N__25199),
            .I(N__25185));
    InMux I__4131 (
            .O(N__25198),
            .I(N__25185));
    InMux I__4130 (
            .O(N__25197),
            .I(N__25185));
    InMux I__4129 (
            .O(N__25196),
            .I(N__25185));
    LocalMux I__4128 (
            .O(N__25185),
            .I(N__25179));
    InMux I__4127 (
            .O(N__25184),
            .I(N__25172));
    InMux I__4126 (
            .O(N__25183),
            .I(N__25172));
    InMux I__4125 (
            .O(N__25182),
            .I(N__25172));
    Odrv4 I__4124 (
            .O(N__25179),
            .I(\c0.tx2_transmit_N_1996 ));
    LocalMux I__4123 (
            .O(N__25172),
            .I(\c0.tx2_transmit_N_1996 ));
    InMux I__4122 (
            .O(N__25167),
            .I(\c0.n16485 ));
    InMux I__4121 (
            .O(N__25164),
            .I(N__25161));
    LocalMux I__4120 (
            .O(N__25161),
            .I(N__25158));
    Odrv4 I__4119 (
            .O(N__25158),
            .I(\c0.n18318 ));
    CascadeMux I__4118 (
            .O(N__25155),
            .I(\c0.n18100_cascade_ ));
    CascadeMux I__4117 (
            .O(N__25152),
            .I(\c0.n18103_cascade_ ));
    CascadeMux I__4116 (
            .O(N__25149),
            .I(\c0.n13808_cascade_ ));
    CascadeMux I__4115 (
            .O(N__25146),
            .I(\c0.n14064_cascade_ ));
    SRMux I__4114 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__4113 (
            .O(N__25140),
            .I(N__25137));
    Span4Mux_s1_v I__4112 (
            .O(N__25137),
            .I(N__25134));
    Odrv4 I__4111 (
            .O(N__25134),
            .I(\c0.n4_adj_2203 ));
    SRMux I__4110 (
            .O(N__25131),
            .I(N__25128));
    LocalMux I__4109 (
            .O(N__25128),
            .I(\c0.n4_adj_2201 ));
    InMux I__4108 (
            .O(N__25125),
            .I(N__25116));
    InMux I__4107 (
            .O(N__25124),
            .I(N__25116));
    InMux I__4106 (
            .O(N__25123),
            .I(N__25116));
    LocalMux I__4105 (
            .O(N__25116),
            .I(N__25110));
    CascadeMux I__4104 (
            .O(N__25115),
            .I(N__25107));
    CascadeMux I__4103 (
            .O(N__25114),
            .I(N__25104));
    CascadeMux I__4102 (
            .O(N__25113),
            .I(N__25101));
    Span4Mux_h I__4101 (
            .O(N__25110),
            .I(N__25095));
    InMux I__4100 (
            .O(N__25107),
            .I(N__25086));
    InMux I__4099 (
            .O(N__25104),
            .I(N__25086));
    InMux I__4098 (
            .O(N__25101),
            .I(N__25086));
    InMux I__4097 (
            .O(N__25100),
            .I(N__25086));
    InMux I__4096 (
            .O(N__25099),
            .I(N__25081));
    InMux I__4095 (
            .O(N__25098),
            .I(N__25081));
    Odrv4 I__4094 (
            .O(N__25095),
            .I(n17694));
    LocalMux I__4093 (
            .O(N__25086),
            .I(n17694));
    LocalMux I__4092 (
            .O(N__25081),
            .I(n17694));
    CascadeMux I__4091 (
            .O(N__25074),
            .I(N__25070));
    InMux I__4090 (
            .O(N__25073),
            .I(N__25062));
    InMux I__4089 (
            .O(N__25070),
            .I(N__25062));
    InMux I__4088 (
            .O(N__25069),
            .I(N__25062));
    LocalMux I__4087 (
            .O(N__25062),
            .I(N__25059));
    Span4Mux_h I__4086 (
            .O(N__25059),
            .I(N__25049));
    InMux I__4085 (
            .O(N__25058),
            .I(N__25046));
    InMux I__4084 (
            .O(N__25057),
            .I(N__25033));
    InMux I__4083 (
            .O(N__25056),
            .I(N__25033));
    InMux I__4082 (
            .O(N__25055),
            .I(N__25033));
    InMux I__4081 (
            .O(N__25054),
            .I(N__25033));
    InMux I__4080 (
            .O(N__25053),
            .I(N__25033));
    InMux I__4079 (
            .O(N__25052),
            .I(N__25033));
    Odrv4 I__4078 (
            .O(N__25049),
            .I(\c0.n43 ));
    LocalMux I__4077 (
            .O(N__25046),
            .I(\c0.n43 ));
    LocalMux I__4076 (
            .O(N__25033),
            .I(\c0.n43 ));
    SRMux I__4075 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__4074 (
            .O(N__25023),
            .I(N__25020));
    Span4Mux_s0_v I__4073 (
            .O(N__25020),
            .I(N__25017));
    Odrv4 I__4072 (
            .O(N__25017),
            .I(\c0.n4_adj_2199 ));
    InMux I__4071 (
            .O(N__25014),
            .I(bfn_7_3_0_));
    InMux I__4070 (
            .O(N__25011),
            .I(N__25008));
    LocalMux I__4069 (
            .O(N__25008),
            .I(N__25005));
    Span4Mux_h I__4068 (
            .O(N__25005),
            .I(N__25002));
    Span4Mux_v I__4067 (
            .O(N__25002),
            .I(N__24999));
    Odrv4 I__4066 (
            .O(N__24999),
            .I(\c0.n18253 ));
    InMux I__4065 (
            .O(N__24996),
            .I(\c0.n16479 ));
    InMux I__4064 (
            .O(N__24993),
            .I(N__24990));
    LocalMux I__4063 (
            .O(N__24990),
            .I(\c0.n18314 ));
    InMux I__4062 (
            .O(N__24987),
            .I(\c0.n16480 ));
    InMux I__4061 (
            .O(N__24984),
            .I(N__24977));
    InMux I__4060 (
            .O(N__24983),
            .I(N__24977));
    InMux I__4059 (
            .O(N__24982),
            .I(N__24974));
    LocalMux I__4058 (
            .O(N__24977),
            .I(blink_counter_22));
    LocalMux I__4057 (
            .O(N__24974),
            .I(blink_counter_22));
    InMux I__4056 (
            .O(N__24969),
            .I(n16630));
    CascadeMux I__4055 (
            .O(N__24966),
            .I(N__24962));
    InMux I__4054 (
            .O(N__24965),
            .I(N__24956));
    InMux I__4053 (
            .O(N__24962),
            .I(N__24956));
    InMux I__4052 (
            .O(N__24961),
            .I(N__24953));
    LocalMux I__4051 (
            .O(N__24956),
            .I(blink_counter_23));
    LocalMux I__4050 (
            .O(N__24953),
            .I(blink_counter_23));
    InMux I__4049 (
            .O(N__24948),
            .I(n16631));
    InMux I__4048 (
            .O(N__24945),
            .I(N__24938));
    InMux I__4047 (
            .O(N__24944),
            .I(N__24938));
    InMux I__4046 (
            .O(N__24943),
            .I(N__24935));
    LocalMux I__4045 (
            .O(N__24938),
            .I(blink_counter_24));
    LocalMux I__4044 (
            .O(N__24935),
            .I(blink_counter_24));
    InMux I__4043 (
            .O(N__24930),
            .I(bfn_6_24_0_));
    InMux I__4042 (
            .O(N__24927),
            .I(n16633));
    InMux I__4041 (
            .O(N__24924),
            .I(N__24920));
    InMux I__4040 (
            .O(N__24923),
            .I(N__24917));
    LocalMux I__4039 (
            .O(N__24920),
            .I(blink_counter_25));
    LocalMux I__4038 (
            .O(N__24917),
            .I(blink_counter_25));
    CEMux I__4037 (
            .O(N__24912),
            .I(N__24909));
    LocalMux I__4036 (
            .O(N__24909),
            .I(N__24906));
    Odrv4 I__4035 (
            .O(N__24906),
            .I(\control.n11 ));
    IoInMux I__4034 (
            .O(N__24903),
            .I(N__24900));
    LocalMux I__4033 (
            .O(N__24900),
            .I(N__24897));
    Span4Mux_s3_v I__4032 (
            .O(N__24897),
            .I(N__24894));
    Odrv4 I__4031 (
            .O(N__24894),
            .I(PIN_1_c_0));
    InMux I__4030 (
            .O(N__24891),
            .I(N__24888));
    LocalMux I__4029 (
            .O(N__24888),
            .I(n12));
    InMux I__4028 (
            .O(N__24885),
            .I(n16622));
    InMux I__4027 (
            .O(N__24882),
            .I(N__24879));
    LocalMux I__4026 (
            .O(N__24879),
            .I(n11));
    InMux I__4025 (
            .O(N__24876),
            .I(n16623));
    InMux I__4024 (
            .O(N__24873),
            .I(N__24870));
    LocalMux I__4023 (
            .O(N__24870),
            .I(n10_adj_2467));
    InMux I__4022 (
            .O(N__24867),
            .I(bfn_6_23_0_));
    InMux I__4021 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__4020 (
            .O(N__24861),
            .I(n9));
    InMux I__4019 (
            .O(N__24858),
            .I(n16625));
    InMux I__4018 (
            .O(N__24855),
            .I(N__24852));
    LocalMux I__4017 (
            .O(N__24852),
            .I(n8));
    InMux I__4016 (
            .O(N__24849),
            .I(n16626));
    InMux I__4015 (
            .O(N__24846),
            .I(N__24843));
    LocalMux I__4014 (
            .O(N__24843),
            .I(n7_adj_2476));
    InMux I__4013 (
            .O(N__24840),
            .I(n16627));
    InMux I__4012 (
            .O(N__24837),
            .I(N__24834));
    LocalMux I__4011 (
            .O(N__24834),
            .I(n6));
    InMux I__4010 (
            .O(N__24831),
            .I(n16628));
    CascadeMux I__4009 (
            .O(N__24828),
            .I(N__24825));
    InMux I__4008 (
            .O(N__24825),
            .I(N__24818));
    InMux I__4007 (
            .O(N__24824),
            .I(N__24818));
    InMux I__4006 (
            .O(N__24823),
            .I(N__24815));
    LocalMux I__4005 (
            .O(N__24818),
            .I(blink_counter_21));
    LocalMux I__4004 (
            .O(N__24815),
            .I(blink_counter_21));
    InMux I__4003 (
            .O(N__24810),
            .I(n16629));
    InMux I__4002 (
            .O(N__24807),
            .I(n16613));
    InMux I__4001 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__4000 (
            .O(N__24801),
            .I(n20));
    InMux I__3999 (
            .O(N__24798),
            .I(n16614));
    InMux I__3998 (
            .O(N__24795),
            .I(N__24792));
    LocalMux I__3997 (
            .O(N__24792),
            .I(n19));
    InMux I__3996 (
            .O(N__24789),
            .I(n16615));
    InMux I__3995 (
            .O(N__24786),
            .I(N__24783));
    LocalMux I__3994 (
            .O(N__24783),
            .I(n18_adj_2480));
    InMux I__3993 (
            .O(N__24780),
            .I(bfn_6_22_0_));
    InMux I__3992 (
            .O(N__24777),
            .I(N__24774));
    LocalMux I__3991 (
            .O(N__24774),
            .I(n17));
    InMux I__3990 (
            .O(N__24771),
            .I(n16617));
    InMux I__3989 (
            .O(N__24768),
            .I(N__24765));
    LocalMux I__3988 (
            .O(N__24765),
            .I(n16));
    InMux I__3987 (
            .O(N__24762),
            .I(n16618));
    InMux I__3986 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__3985 (
            .O(N__24756),
            .I(n15_adj_2479));
    InMux I__3984 (
            .O(N__24753),
            .I(n16619));
    InMux I__3983 (
            .O(N__24750),
            .I(N__24747));
    LocalMux I__3982 (
            .O(N__24747),
            .I(n14_adj_2478));
    InMux I__3981 (
            .O(N__24744),
            .I(n16620));
    InMux I__3980 (
            .O(N__24741),
            .I(N__24738));
    LocalMux I__3979 (
            .O(N__24738),
            .I(n13));
    InMux I__3978 (
            .O(N__24735),
            .I(n16621));
    CascadeMux I__3977 (
            .O(N__24732),
            .I(\c0.rx.n12_cascade_ ));
    CEMux I__3976 (
            .O(N__24729),
            .I(N__24726));
    LocalMux I__3975 (
            .O(N__24726),
            .I(N__24723));
    Span4Mux_h I__3974 (
            .O(N__24723),
            .I(N__24720));
    Odrv4 I__3973 (
            .O(N__24720),
            .I(\c0.rx.n11082 ));
    InMux I__3972 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__3971 (
            .O(N__24714),
            .I(N__24711));
    Span4Mux_v I__3970 (
            .O(N__24711),
            .I(N__24708));
    Odrv4 I__3969 (
            .O(N__24708),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_18 ));
    InMux I__3968 (
            .O(N__24705),
            .I(N__24700));
    CascadeMux I__3967 (
            .O(N__24704),
            .I(N__24696));
    InMux I__3966 (
            .O(N__24703),
            .I(N__24693));
    LocalMux I__3965 (
            .O(N__24700),
            .I(N__24690));
    InMux I__3964 (
            .O(N__24699),
            .I(N__24687));
    InMux I__3963 (
            .O(N__24696),
            .I(N__24684));
    LocalMux I__3962 (
            .O(N__24693),
            .I(N__24681));
    Span4Mux_v I__3961 (
            .O(N__24690),
            .I(N__24678));
    LocalMux I__3960 (
            .O(N__24687),
            .I(N__24673));
    LocalMux I__3959 (
            .O(N__24684),
            .I(N__24673));
    Span4Mux_h I__3958 (
            .O(N__24681),
            .I(N__24670));
    Span4Mux_h I__3957 (
            .O(N__24678),
            .I(N__24665));
    Span4Mux_h I__3956 (
            .O(N__24673),
            .I(N__24665));
    Odrv4 I__3955 (
            .O(N__24670),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__3954 (
            .O(N__24665),
            .I(\c0.FRAME_MATCHER_i_18 ));
    SRMux I__3953 (
            .O(N__24660),
            .I(N__24657));
    LocalMux I__3952 (
            .O(N__24657),
            .I(N__24654));
    Span4Mux_h I__3951 (
            .O(N__24654),
            .I(N__24651));
    Span4Mux_v I__3950 (
            .O(N__24651),
            .I(N__24648));
    Odrv4 I__3949 (
            .O(N__24648),
            .I(\c0.n3_adj_2305 ));
    InMux I__3948 (
            .O(N__24645),
            .I(N__24640));
    InMux I__3947 (
            .O(N__24644),
            .I(N__24637));
    InMux I__3946 (
            .O(N__24643),
            .I(N__24634));
    LocalMux I__3945 (
            .O(N__24640),
            .I(N__24617));
    LocalMux I__3944 (
            .O(N__24637),
            .I(N__24612));
    LocalMux I__3943 (
            .O(N__24634),
            .I(N__24612));
    InMux I__3942 (
            .O(N__24633),
            .I(N__24609));
    InMux I__3941 (
            .O(N__24632),
            .I(N__24606));
    InMux I__3940 (
            .O(N__24631),
            .I(N__24603));
    InMux I__3939 (
            .O(N__24630),
            .I(N__24600));
    InMux I__3938 (
            .O(N__24629),
            .I(N__24596));
    InMux I__3937 (
            .O(N__24628),
            .I(N__24593));
    InMux I__3936 (
            .O(N__24627),
            .I(N__24590));
    InMux I__3935 (
            .O(N__24626),
            .I(N__24587));
    InMux I__3934 (
            .O(N__24625),
            .I(N__24582));
    InMux I__3933 (
            .O(N__24624),
            .I(N__24579));
    InMux I__3932 (
            .O(N__24623),
            .I(N__24576));
    InMux I__3931 (
            .O(N__24622),
            .I(N__24573));
    InMux I__3930 (
            .O(N__24621),
            .I(N__24570));
    InMux I__3929 (
            .O(N__24620),
            .I(N__24562));
    Span4Mux_h I__3928 (
            .O(N__24617),
            .I(N__24549));
    Span4Mux_v I__3927 (
            .O(N__24612),
            .I(N__24549));
    LocalMux I__3926 (
            .O(N__24609),
            .I(N__24549));
    LocalMux I__3925 (
            .O(N__24606),
            .I(N__24549));
    LocalMux I__3924 (
            .O(N__24603),
            .I(N__24549));
    LocalMux I__3923 (
            .O(N__24600),
            .I(N__24549));
    InMux I__3922 (
            .O(N__24599),
            .I(N__24546));
    LocalMux I__3921 (
            .O(N__24596),
            .I(N__24537));
    LocalMux I__3920 (
            .O(N__24593),
            .I(N__24537));
    LocalMux I__3919 (
            .O(N__24590),
            .I(N__24537));
    LocalMux I__3918 (
            .O(N__24587),
            .I(N__24537));
    InMux I__3917 (
            .O(N__24586),
            .I(N__24534));
    InMux I__3916 (
            .O(N__24585),
            .I(N__24530));
    LocalMux I__3915 (
            .O(N__24582),
            .I(N__24519));
    LocalMux I__3914 (
            .O(N__24579),
            .I(N__24519));
    LocalMux I__3913 (
            .O(N__24576),
            .I(N__24519));
    LocalMux I__3912 (
            .O(N__24573),
            .I(N__24519));
    LocalMux I__3911 (
            .O(N__24570),
            .I(N__24519));
    InMux I__3910 (
            .O(N__24569),
            .I(N__24516));
    InMux I__3909 (
            .O(N__24568),
            .I(N__24513));
    InMux I__3908 (
            .O(N__24567),
            .I(N__24510));
    InMux I__3907 (
            .O(N__24566),
            .I(N__24507));
    InMux I__3906 (
            .O(N__24565),
            .I(N__24504));
    LocalMux I__3905 (
            .O(N__24562),
            .I(N__24495));
    Span4Mux_v I__3904 (
            .O(N__24549),
            .I(N__24490));
    LocalMux I__3903 (
            .O(N__24546),
            .I(N__24490));
    Span4Mux_v I__3902 (
            .O(N__24537),
            .I(N__24485));
    LocalMux I__3901 (
            .O(N__24534),
            .I(N__24485));
    InMux I__3900 (
            .O(N__24533),
            .I(N__24482));
    LocalMux I__3899 (
            .O(N__24530),
            .I(N__24469));
    Span4Mux_v I__3898 (
            .O(N__24519),
            .I(N__24469));
    LocalMux I__3897 (
            .O(N__24516),
            .I(N__24469));
    LocalMux I__3896 (
            .O(N__24513),
            .I(N__24469));
    LocalMux I__3895 (
            .O(N__24510),
            .I(N__24469));
    LocalMux I__3894 (
            .O(N__24507),
            .I(N__24469));
    LocalMux I__3893 (
            .O(N__24504),
            .I(N__24466));
    InMux I__3892 (
            .O(N__24503),
            .I(N__24463));
    InMux I__3891 (
            .O(N__24502),
            .I(N__24460));
    InMux I__3890 (
            .O(N__24501),
            .I(N__24457));
    InMux I__3889 (
            .O(N__24500),
            .I(N__24454));
    InMux I__3888 (
            .O(N__24499),
            .I(N__24449));
    InMux I__3887 (
            .O(N__24498),
            .I(N__24449));
    Span12Mux_v I__3886 (
            .O(N__24495),
            .I(N__24443));
    Span4Mux_v I__3885 (
            .O(N__24490),
            .I(N__24438));
    Span4Mux_v I__3884 (
            .O(N__24485),
            .I(N__24438));
    LocalMux I__3883 (
            .O(N__24482),
            .I(N__24435));
    Span4Mux_v I__3882 (
            .O(N__24469),
            .I(N__24428));
    Span4Mux_s2_h I__3881 (
            .O(N__24466),
            .I(N__24428));
    LocalMux I__3880 (
            .O(N__24463),
            .I(N__24428));
    LocalMux I__3879 (
            .O(N__24460),
            .I(N__24425));
    LocalMux I__3878 (
            .O(N__24457),
            .I(N__24418));
    LocalMux I__3877 (
            .O(N__24454),
            .I(N__24418));
    LocalMux I__3876 (
            .O(N__24449),
            .I(N__24418));
    InMux I__3875 (
            .O(N__24448),
            .I(N__24415));
    InMux I__3874 (
            .O(N__24447),
            .I(N__24410));
    InMux I__3873 (
            .O(N__24446),
            .I(N__24410));
    Odrv12 I__3872 (
            .O(N__24443),
            .I(n1166));
    Odrv4 I__3871 (
            .O(N__24438),
            .I(n1166));
    Odrv4 I__3870 (
            .O(N__24435),
            .I(n1166));
    Odrv4 I__3869 (
            .O(N__24428),
            .I(n1166));
    Odrv4 I__3868 (
            .O(N__24425),
            .I(n1166));
    Odrv12 I__3867 (
            .O(N__24418),
            .I(n1166));
    LocalMux I__3866 (
            .O(N__24415),
            .I(n1166));
    LocalMux I__3865 (
            .O(N__24410),
            .I(n1166));
    InMux I__3864 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__3863 (
            .O(N__24390),
            .I(N__24387));
    Span4Mux_v I__3862 (
            .O(N__24387),
            .I(N__24384));
    Odrv4 I__3861 (
            .O(N__24384),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_13 ));
    CascadeMux I__3860 (
            .O(N__24381),
            .I(N__24375));
    CascadeMux I__3859 (
            .O(N__24380),
            .I(N__24372));
    InMux I__3858 (
            .O(N__24379),
            .I(N__24369));
    InMux I__3857 (
            .O(N__24378),
            .I(N__24366));
    InMux I__3856 (
            .O(N__24375),
            .I(N__24363));
    InMux I__3855 (
            .O(N__24372),
            .I(N__24360));
    LocalMux I__3854 (
            .O(N__24369),
            .I(N__24351));
    LocalMux I__3853 (
            .O(N__24366),
            .I(N__24351));
    LocalMux I__3852 (
            .O(N__24363),
            .I(N__24351));
    LocalMux I__3851 (
            .O(N__24360),
            .I(N__24351));
    Span4Mux_h I__3850 (
            .O(N__24351),
            .I(N__24348));
    Odrv4 I__3849 (
            .O(N__24348),
            .I(\c0.FRAME_MATCHER_i_13 ));
    SRMux I__3848 (
            .O(N__24345),
            .I(N__24342));
    LocalMux I__3847 (
            .O(N__24342),
            .I(N__24339));
    Span4Mux_h I__3846 (
            .O(N__24339),
            .I(N__24336));
    Span4Mux_v I__3845 (
            .O(N__24336),
            .I(N__24333));
    Odrv4 I__3844 (
            .O(N__24333),
            .I(\c0.n3_adj_2317 ));
    InMux I__3843 (
            .O(N__24330),
            .I(N__24327));
    LocalMux I__3842 (
            .O(N__24327),
            .I(n26));
    InMux I__3841 (
            .O(N__24324),
            .I(bfn_6_21_0_));
    InMux I__3840 (
            .O(N__24321),
            .I(N__24318));
    LocalMux I__3839 (
            .O(N__24318),
            .I(n25));
    InMux I__3838 (
            .O(N__24315),
            .I(n16609));
    InMux I__3837 (
            .O(N__24312),
            .I(N__24309));
    LocalMux I__3836 (
            .O(N__24309),
            .I(n24));
    InMux I__3835 (
            .O(N__24306),
            .I(n16610));
    InMux I__3834 (
            .O(N__24303),
            .I(N__24300));
    LocalMux I__3833 (
            .O(N__24300),
            .I(n23));
    InMux I__3832 (
            .O(N__24297),
            .I(n16611));
    InMux I__3831 (
            .O(N__24294),
            .I(N__24291));
    LocalMux I__3830 (
            .O(N__24291),
            .I(n22_adj_2481));
    InMux I__3829 (
            .O(N__24288),
            .I(n16612));
    InMux I__3828 (
            .O(N__24285),
            .I(N__24282));
    LocalMux I__3827 (
            .O(N__24282),
            .I(n21));
    InMux I__3826 (
            .O(N__24279),
            .I(\c0.rx.n16536 ));
    InMux I__3825 (
            .O(N__24276),
            .I(\c0.rx.n16537 ));
    InMux I__3824 (
            .O(N__24273),
            .I(\c0.rx.n16538 ));
    SRMux I__3823 (
            .O(N__24270),
            .I(N__24267));
    LocalMux I__3822 (
            .O(N__24267),
            .I(N__24264));
    Odrv4 I__3821 (
            .O(N__24264),
            .I(\c0.rx.n12819 ));
    CascadeMux I__3820 (
            .O(N__24261),
            .I(\c0.n18225_cascade_ ));
    InMux I__3819 (
            .O(N__24258),
            .I(N__24255));
    LocalMux I__3818 (
            .O(N__24255),
            .I(N__24252));
    Span4Mux_v I__3817 (
            .O(N__24252),
            .I(N__24249));
    Span4Mux_h I__3816 (
            .O(N__24249),
            .I(N__24246));
    Odrv4 I__3815 (
            .O(N__24246),
            .I(\c0.rx.n5 ));
    InMux I__3814 (
            .O(N__24243),
            .I(N__24240));
    LocalMux I__3813 (
            .O(N__24240),
            .I(N__24237));
    Span4Mux_v I__3812 (
            .O(N__24237),
            .I(N__24234));
    Span4Mux_h I__3811 (
            .O(N__24234),
            .I(N__24231));
    Odrv4 I__3810 (
            .O(N__24231),
            .I(\c0.rx.n57 ));
    CascadeMux I__3809 (
            .O(N__24228),
            .I(\c0.rx.n15905_cascade_ ));
    CascadeMux I__3808 (
            .O(N__24225),
            .I(\c0.rx.n6_cascade_ ));
    InMux I__3807 (
            .O(N__24222),
            .I(N__24219));
    LocalMux I__3806 (
            .O(N__24219),
            .I(\c0.rx.n12 ));
    InMux I__3805 (
            .O(N__24216),
            .I(N__24208));
    InMux I__3804 (
            .O(N__24215),
            .I(N__24208));
    InMux I__3803 (
            .O(N__24214),
            .I(N__24203));
    InMux I__3802 (
            .O(N__24213),
            .I(N__24203));
    LocalMux I__3801 (
            .O(N__24208),
            .I(data_in_2_7));
    LocalMux I__3800 (
            .O(N__24203),
            .I(data_in_2_7));
    InMux I__3799 (
            .O(N__24198),
            .I(N__24192));
    InMux I__3798 (
            .O(N__24197),
            .I(N__24185));
    InMux I__3797 (
            .O(N__24196),
            .I(N__24185));
    InMux I__3796 (
            .O(N__24195),
            .I(N__24185));
    LocalMux I__3795 (
            .O(N__24192),
            .I(data_in_2_5));
    LocalMux I__3794 (
            .O(N__24185),
            .I(data_in_2_5));
    CascadeMux I__3793 (
            .O(N__24180),
            .I(N__24174));
    InMux I__3792 (
            .O(N__24179),
            .I(N__24171));
    InMux I__3791 (
            .O(N__24178),
            .I(N__24166));
    InMux I__3790 (
            .O(N__24177),
            .I(N__24166));
    InMux I__3789 (
            .O(N__24174),
            .I(N__24162));
    LocalMux I__3788 (
            .O(N__24171),
            .I(N__24159));
    LocalMux I__3787 (
            .O(N__24166),
            .I(N__24156));
    CascadeMux I__3786 (
            .O(N__24165),
            .I(N__24150));
    LocalMux I__3785 (
            .O(N__24162),
            .I(N__24147));
    Span4Mux_v I__3784 (
            .O(N__24159),
            .I(N__24142));
    Span4Mux_v I__3783 (
            .O(N__24156),
            .I(N__24142));
    InMux I__3782 (
            .O(N__24155),
            .I(N__24139));
    InMux I__3781 (
            .O(N__24154),
            .I(N__24136));
    InMux I__3780 (
            .O(N__24153),
            .I(N__24133));
    InMux I__3779 (
            .O(N__24150),
            .I(N__24130));
    Odrv12 I__3778 (
            .O(N__24147),
            .I(rx_data_7));
    Odrv4 I__3777 (
            .O(N__24142),
            .I(rx_data_7));
    LocalMux I__3776 (
            .O(N__24139),
            .I(rx_data_7));
    LocalMux I__3775 (
            .O(N__24136),
            .I(rx_data_7));
    LocalMux I__3774 (
            .O(N__24133),
            .I(rx_data_7));
    LocalMux I__3773 (
            .O(N__24130),
            .I(rx_data_7));
    InMux I__3772 (
            .O(N__24117),
            .I(bfn_6_13_0_));
    InMux I__3771 (
            .O(N__24114),
            .I(\c0.rx.n16532 ));
    InMux I__3770 (
            .O(N__24111),
            .I(\c0.rx.n16533 ));
    InMux I__3769 (
            .O(N__24108),
            .I(\c0.rx.n16534 ));
    InMux I__3768 (
            .O(N__24105),
            .I(\c0.rx.n16535 ));
    InMux I__3767 (
            .O(N__24102),
            .I(N__24098));
    InMux I__3766 (
            .O(N__24101),
            .I(N__24094));
    LocalMux I__3765 (
            .O(N__24098),
            .I(N__24091));
    InMux I__3764 (
            .O(N__24097),
            .I(N__24088));
    LocalMux I__3763 (
            .O(N__24094),
            .I(data_in_1_5));
    Odrv4 I__3762 (
            .O(N__24091),
            .I(data_in_1_5));
    LocalMux I__3761 (
            .O(N__24088),
            .I(data_in_1_5));
    CascadeMux I__3760 (
            .O(N__24081),
            .I(N__24076));
    InMux I__3759 (
            .O(N__24080),
            .I(N__24073));
    InMux I__3758 (
            .O(N__24079),
            .I(N__24070));
    InMux I__3757 (
            .O(N__24076),
            .I(N__24067));
    LocalMux I__3756 (
            .O(N__24073),
            .I(data_in_2_4));
    LocalMux I__3755 (
            .O(N__24070),
            .I(data_in_2_4));
    LocalMux I__3754 (
            .O(N__24067),
            .I(data_in_2_4));
    InMux I__3753 (
            .O(N__24060),
            .I(N__24057));
    LocalMux I__3752 (
            .O(N__24057),
            .I(\c0.n18_adj_2370 ));
    CascadeMux I__3751 (
            .O(N__24054),
            .I(N__24051));
    InMux I__3750 (
            .O(N__24051),
            .I(N__24048));
    LocalMux I__3749 (
            .O(N__24048),
            .I(\c0.n13_adj_2380 ));
    InMux I__3748 (
            .O(N__24045),
            .I(N__24042));
    LocalMux I__3747 (
            .O(N__24042),
            .I(N__24038));
    InMux I__3746 (
            .O(N__24041),
            .I(N__24035));
    Odrv4 I__3745 (
            .O(N__24038),
            .I(\c0.rx.n10988 ));
    LocalMux I__3744 (
            .O(N__24035),
            .I(\c0.rx.n10988 ));
    CascadeMux I__3743 (
            .O(N__24030),
            .I(\c0.n18006_cascade_ ));
    InMux I__3742 (
            .O(N__24027),
            .I(N__24024));
    LocalMux I__3741 (
            .O(N__24024),
            .I(N__24021));
    Odrv4 I__3740 (
            .O(N__24021),
            .I(\c0.n14_adj_2375 ));
    CascadeMux I__3739 (
            .O(N__24018),
            .I(\c0.n20_adj_2371_cascade_ ));
    InMux I__3738 (
            .O(N__24015),
            .I(N__24012));
    LocalMux I__3737 (
            .O(N__24012),
            .I(\c0.n10516 ));
    CascadeMux I__3736 (
            .O(N__24009),
            .I(\c0.n10516_cascade_ ));
    InMux I__3735 (
            .O(N__24006),
            .I(N__24003));
    LocalMux I__3734 (
            .O(N__24003),
            .I(\c0.n10367 ));
    InMux I__3733 (
            .O(N__24000),
            .I(N__23995));
    InMux I__3732 (
            .O(N__23999),
            .I(N__23990));
    InMux I__3731 (
            .O(N__23998),
            .I(N__23990));
    LocalMux I__3730 (
            .O(N__23995),
            .I(data_in_0_5));
    LocalMux I__3729 (
            .O(N__23990),
            .I(data_in_0_5));
    CascadeMux I__3728 (
            .O(N__23985),
            .I(\c0.n10367_cascade_ ));
    InMux I__3727 (
            .O(N__23982),
            .I(N__23979));
    LocalMux I__3726 (
            .O(N__23979),
            .I(\c0.n15_adj_2389 ));
    CascadeMux I__3725 (
            .O(N__23976),
            .I(N__23973));
    InMux I__3724 (
            .O(N__23973),
            .I(N__23969));
    InMux I__3723 (
            .O(N__23972),
            .I(N__23964));
    LocalMux I__3722 (
            .O(N__23969),
            .I(N__23961));
    InMux I__3721 (
            .O(N__23968),
            .I(N__23956));
    InMux I__3720 (
            .O(N__23967),
            .I(N__23956));
    LocalMux I__3719 (
            .O(N__23964),
            .I(data_in_1_4));
    Odrv4 I__3718 (
            .O(N__23961),
            .I(data_in_1_4));
    LocalMux I__3717 (
            .O(N__23956),
            .I(data_in_1_4));
    InMux I__3716 (
            .O(N__23949),
            .I(N__23943));
    InMux I__3715 (
            .O(N__23948),
            .I(N__23943));
    LocalMux I__3714 (
            .O(N__23943),
            .I(data_in_0_4));
    InMux I__3713 (
            .O(N__23940),
            .I(N__23932));
    InMux I__3712 (
            .O(N__23939),
            .I(N__23932));
    InMux I__3711 (
            .O(N__23938),
            .I(N__23927));
    InMux I__3710 (
            .O(N__23937),
            .I(N__23927));
    LocalMux I__3709 (
            .O(N__23932),
            .I(data_in_3_4));
    LocalMux I__3708 (
            .O(N__23927),
            .I(data_in_3_4));
    InMux I__3707 (
            .O(N__23922),
            .I(N__23919));
    LocalMux I__3706 (
            .O(N__23919),
            .I(\c0.n14_adj_2388 ));
    CascadeMux I__3705 (
            .O(N__23916),
            .I(N__23902));
    CascadeMux I__3704 (
            .O(N__23915),
            .I(N__23898));
    CascadeMux I__3703 (
            .O(N__23914),
            .I(N__23894));
    CascadeMux I__3702 (
            .O(N__23913),
            .I(N__23890));
    CascadeMux I__3701 (
            .O(N__23912),
            .I(N__23887));
    CascadeMux I__3700 (
            .O(N__23911),
            .I(N__23882));
    CascadeMux I__3699 (
            .O(N__23910),
            .I(N__23878));
    CascadeMux I__3698 (
            .O(N__23909),
            .I(N__23872));
    CascadeMux I__3697 (
            .O(N__23908),
            .I(N__23868));
    CascadeMux I__3696 (
            .O(N__23907),
            .I(N__23864));
    CascadeMux I__3695 (
            .O(N__23906),
            .I(N__23860));
    InMux I__3694 (
            .O(N__23905),
            .I(N__23846));
    InMux I__3693 (
            .O(N__23902),
            .I(N__23846));
    InMux I__3692 (
            .O(N__23901),
            .I(N__23846));
    InMux I__3691 (
            .O(N__23898),
            .I(N__23835));
    InMux I__3690 (
            .O(N__23897),
            .I(N__23835));
    InMux I__3689 (
            .O(N__23894),
            .I(N__23835));
    InMux I__3688 (
            .O(N__23893),
            .I(N__23835));
    InMux I__3687 (
            .O(N__23890),
            .I(N__23835));
    InMux I__3686 (
            .O(N__23887),
            .I(N__23824));
    InMux I__3685 (
            .O(N__23886),
            .I(N__23824));
    InMux I__3684 (
            .O(N__23885),
            .I(N__23824));
    InMux I__3683 (
            .O(N__23882),
            .I(N__23824));
    InMux I__3682 (
            .O(N__23881),
            .I(N__23824));
    InMux I__3681 (
            .O(N__23878),
            .I(N__23817));
    InMux I__3680 (
            .O(N__23877),
            .I(N__23817));
    InMux I__3679 (
            .O(N__23876),
            .I(N__23817));
    InMux I__3678 (
            .O(N__23875),
            .I(N__23800));
    InMux I__3677 (
            .O(N__23872),
            .I(N__23800));
    InMux I__3676 (
            .O(N__23871),
            .I(N__23800));
    InMux I__3675 (
            .O(N__23868),
            .I(N__23800));
    InMux I__3674 (
            .O(N__23867),
            .I(N__23800));
    InMux I__3673 (
            .O(N__23864),
            .I(N__23800));
    InMux I__3672 (
            .O(N__23863),
            .I(N__23800));
    InMux I__3671 (
            .O(N__23860),
            .I(N__23800));
    CascadeMux I__3670 (
            .O(N__23859),
            .I(N__23797));
    CascadeMux I__3669 (
            .O(N__23858),
            .I(N__23794));
    CascadeMux I__3668 (
            .O(N__23857),
            .I(N__23791));
    CascadeMux I__3667 (
            .O(N__23856),
            .I(N__23787));
    CascadeMux I__3666 (
            .O(N__23855),
            .I(N__23784));
    CascadeMux I__3665 (
            .O(N__23854),
            .I(N__23781));
    CascadeMux I__3664 (
            .O(N__23853),
            .I(N__23778));
    LocalMux I__3663 (
            .O(N__23846),
            .I(N__23775));
    LocalMux I__3662 (
            .O(N__23835),
            .I(N__23772));
    LocalMux I__3661 (
            .O(N__23824),
            .I(N__23767));
    LocalMux I__3660 (
            .O(N__23817),
            .I(N__23767));
    LocalMux I__3659 (
            .O(N__23800),
            .I(N__23764));
    InMux I__3658 (
            .O(N__23797),
            .I(N__23753));
    InMux I__3657 (
            .O(N__23794),
            .I(N__23753));
    InMux I__3656 (
            .O(N__23791),
            .I(N__23753));
    InMux I__3655 (
            .O(N__23790),
            .I(N__23753));
    InMux I__3654 (
            .O(N__23787),
            .I(N__23753));
    InMux I__3653 (
            .O(N__23784),
            .I(N__23746));
    InMux I__3652 (
            .O(N__23781),
            .I(N__23746));
    InMux I__3651 (
            .O(N__23778),
            .I(N__23746));
    Span4Mux_h I__3650 (
            .O(N__23775),
            .I(N__23743));
    Span4Mux_h I__3649 (
            .O(N__23772),
            .I(N__23740));
    Span12Mux_s5_h I__3648 (
            .O(N__23767),
            .I(N__23737));
    Span4Mux_h I__3647 (
            .O(N__23764),
            .I(N__23734));
    LocalMux I__3646 (
            .O(N__23753),
            .I(N__23729));
    LocalMux I__3645 (
            .O(N__23746),
            .I(N__23729));
    Odrv4 I__3644 (
            .O(N__23743),
            .I(\c0.n18631 ));
    Odrv4 I__3643 (
            .O(N__23740),
            .I(\c0.n18631 ));
    Odrv12 I__3642 (
            .O(N__23737),
            .I(\c0.n18631 ));
    Odrv4 I__3641 (
            .O(N__23734),
            .I(\c0.n18631 ));
    Odrv4 I__3640 (
            .O(N__23729),
            .I(\c0.n18631 ));
    CascadeMux I__3639 (
            .O(N__23718),
            .I(\c0.n18002_cascade_ ));
    InMux I__3638 (
            .O(N__23715),
            .I(N__23709));
    InMux I__3637 (
            .O(N__23714),
            .I(N__23709));
    LocalMux I__3636 (
            .O(N__23709),
            .I(\c0.n10498 ));
    CascadeMux I__3635 (
            .O(N__23706),
            .I(\c0.rx.n10988_cascade_ ));
    CascadeMux I__3634 (
            .O(N__23703),
            .I(\c0.rx.n12624_cascade_ ));
    InMux I__3633 (
            .O(N__23700),
            .I(N__23694));
    InMux I__3632 (
            .O(N__23699),
            .I(N__23694));
    LocalMux I__3631 (
            .O(N__23694),
            .I(data_in_0_2));
    InMux I__3630 (
            .O(N__23691),
            .I(N__23687));
    InMux I__3629 (
            .O(N__23690),
            .I(N__23684));
    LocalMux I__3628 (
            .O(N__23687),
            .I(data_in_frame_5_7));
    LocalMux I__3627 (
            .O(N__23684),
            .I(data_in_frame_5_7));
    InMux I__3626 (
            .O(N__23679),
            .I(N__23675));
    CascadeMux I__3625 (
            .O(N__23678),
            .I(N__23671));
    LocalMux I__3624 (
            .O(N__23675),
            .I(N__23668));
    InMux I__3623 (
            .O(N__23674),
            .I(N__23665));
    InMux I__3622 (
            .O(N__23671),
            .I(N__23662));
    Span4Mux_h I__3621 (
            .O(N__23668),
            .I(N__23659));
    LocalMux I__3620 (
            .O(N__23665),
            .I(data_in_frame_2_7));
    LocalMux I__3619 (
            .O(N__23662),
            .I(data_in_frame_2_7));
    Odrv4 I__3618 (
            .O(N__23659),
            .I(data_in_frame_2_7));
    CascadeMux I__3617 (
            .O(N__23652),
            .I(\c0.rx.n17702_cascade_ ));
    CascadeMux I__3616 (
            .O(N__23649),
            .I(N__23646));
    InMux I__3615 (
            .O(N__23646),
            .I(N__23643));
    LocalMux I__3614 (
            .O(N__23643),
            .I(\c0.rx.n17702 ));
    CascadeMux I__3613 (
            .O(N__23640),
            .I(\c0.rx.n17704_cascade_ ));
    InMux I__3612 (
            .O(N__23637),
            .I(N__23630));
    InMux I__3611 (
            .O(N__23636),
            .I(N__23627));
    InMux I__3610 (
            .O(N__23635),
            .I(N__23622));
    InMux I__3609 (
            .O(N__23634),
            .I(N__23617));
    InMux I__3608 (
            .O(N__23633),
            .I(N__23617));
    LocalMux I__3607 (
            .O(N__23630),
            .I(N__23614));
    LocalMux I__3606 (
            .O(N__23627),
            .I(N__23611));
    InMux I__3605 (
            .O(N__23626),
            .I(N__23608));
    InMux I__3604 (
            .O(N__23625),
            .I(N__23605));
    LocalMux I__3603 (
            .O(N__23622),
            .I(n11058));
    LocalMux I__3602 (
            .O(N__23617),
            .I(n11058));
    Odrv4 I__3601 (
            .O(N__23614),
            .I(n11058));
    Odrv4 I__3600 (
            .O(N__23611),
            .I(n11058));
    LocalMux I__3599 (
            .O(N__23608),
            .I(n11058));
    LocalMux I__3598 (
            .O(N__23605),
            .I(n11058));
    InMux I__3597 (
            .O(N__23592),
            .I(N__23583));
    InMux I__3596 (
            .O(N__23591),
            .I(N__23580));
    InMux I__3595 (
            .O(N__23590),
            .I(N__23575));
    InMux I__3594 (
            .O(N__23589),
            .I(N__23575));
    InMux I__3593 (
            .O(N__23588),
            .I(N__23570));
    InMux I__3592 (
            .O(N__23587),
            .I(N__23570));
    InMux I__3591 (
            .O(N__23586),
            .I(N__23567));
    LocalMux I__3590 (
            .O(N__23583),
            .I(n16802));
    LocalMux I__3589 (
            .O(N__23580),
            .I(n16802));
    LocalMux I__3588 (
            .O(N__23575),
            .I(n16802));
    LocalMux I__3587 (
            .O(N__23570),
            .I(n16802));
    LocalMux I__3586 (
            .O(N__23567),
            .I(n16802));
    InMux I__3585 (
            .O(N__23556),
            .I(N__23551));
    InMux I__3584 (
            .O(N__23555),
            .I(N__23548));
    InMux I__3583 (
            .O(N__23554),
            .I(N__23545));
    LocalMux I__3582 (
            .O(N__23551),
            .I(\c0.n10569 ));
    LocalMux I__3581 (
            .O(N__23548),
            .I(\c0.n10569 ));
    LocalMux I__3580 (
            .O(N__23545),
            .I(\c0.n10569 ));
    InMux I__3579 (
            .O(N__23538),
            .I(N__23534));
    InMux I__3578 (
            .O(N__23537),
            .I(N__23531));
    LocalMux I__3577 (
            .O(N__23534),
            .I(N__23528));
    LocalMux I__3576 (
            .O(N__23531),
            .I(data_in_frame_6_3));
    Odrv4 I__3575 (
            .O(N__23528),
            .I(data_in_frame_6_3));
    CascadeMux I__3574 (
            .O(N__23523),
            .I(\c0.n17734_cascade_ ));
    CascadeMux I__3573 (
            .O(N__23520),
            .I(N__23516));
    InMux I__3572 (
            .O(N__23519),
            .I(N__23511));
    InMux I__3571 (
            .O(N__23516),
            .I(N__23508));
    InMux I__3570 (
            .O(N__23515),
            .I(N__23503));
    InMux I__3569 (
            .O(N__23514),
            .I(N__23503));
    LocalMux I__3568 (
            .O(N__23511),
            .I(\c0.data_in_frame_1_7 ));
    LocalMux I__3567 (
            .O(N__23508),
            .I(\c0.data_in_frame_1_7 ));
    LocalMux I__3566 (
            .O(N__23503),
            .I(\c0.data_in_frame_1_7 ));
    InMux I__3565 (
            .O(N__23496),
            .I(N__23493));
    LocalMux I__3564 (
            .O(N__23493),
            .I(\c0.n19_adj_2400 ));
    InMux I__3563 (
            .O(N__23490),
            .I(N__23487));
    LocalMux I__3562 (
            .O(N__23487),
            .I(\c0.n18_adj_2398 ));
    CascadeMux I__3561 (
            .O(N__23484),
            .I(\c0.n18000_cascade_ ));
    InMux I__3560 (
            .O(N__23481),
            .I(N__23477));
    InMux I__3559 (
            .O(N__23480),
            .I(N__23474));
    LocalMux I__3558 (
            .O(N__23477),
            .I(N__23471));
    LocalMux I__3557 (
            .O(N__23474),
            .I(data_in_frame_5_2));
    Odrv4 I__3556 (
            .O(N__23471),
            .I(data_in_frame_5_2));
    InMux I__3555 (
            .O(N__23466),
            .I(N__23463));
    LocalMux I__3554 (
            .O(N__23463),
            .I(N__23457));
    InMux I__3553 (
            .O(N__23462),
            .I(N__23454));
    InMux I__3552 (
            .O(N__23461),
            .I(N__23450));
    InMux I__3551 (
            .O(N__23460),
            .I(N__23447));
    Span4Mux_v I__3550 (
            .O(N__23457),
            .I(N__23440));
    LocalMux I__3549 (
            .O(N__23454),
            .I(N__23440));
    InMux I__3548 (
            .O(N__23453),
            .I(N__23437));
    LocalMux I__3547 (
            .O(N__23450),
            .I(N__23434));
    LocalMux I__3546 (
            .O(N__23447),
            .I(N__23431));
    InMux I__3545 (
            .O(N__23446),
            .I(N__23428));
    InMux I__3544 (
            .O(N__23445),
            .I(N__23424));
    Span4Mux_v I__3543 (
            .O(N__23440),
            .I(N__23421));
    LocalMux I__3542 (
            .O(N__23437),
            .I(N__23414));
    Span4Mux_v I__3541 (
            .O(N__23434),
            .I(N__23414));
    Span4Mux_v I__3540 (
            .O(N__23431),
            .I(N__23414));
    LocalMux I__3539 (
            .O(N__23428),
            .I(N__23411));
    InMux I__3538 (
            .O(N__23427),
            .I(N__23408));
    LocalMux I__3537 (
            .O(N__23424),
            .I(N__23405));
    Sp12to4 I__3536 (
            .O(N__23421),
            .I(N__23398));
    Span4Mux_h I__3535 (
            .O(N__23414),
            .I(N__23393));
    Span4Mux_h I__3534 (
            .O(N__23411),
            .I(N__23393));
    LocalMux I__3533 (
            .O(N__23408),
            .I(N__23388));
    Span4Mux_s2_h I__3532 (
            .O(N__23405),
            .I(N__23388));
    InMux I__3531 (
            .O(N__23404),
            .I(N__23381));
    InMux I__3530 (
            .O(N__23403),
            .I(N__23381));
    InMux I__3529 (
            .O(N__23402),
            .I(N__23381));
    InMux I__3528 (
            .O(N__23401),
            .I(N__23378));
    Odrv12 I__3527 (
            .O(N__23398),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__3526 (
            .O(N__23393),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__3525 (
            .O(N__23388),
            .I(\c0.FRAME_MATCHER_i_0 ));
    LocalMux I__3524 (
            .O(N__23381),
            .I(\c0.FRAME_MATCHER_i_0 ));
    LocalMux I__3523 (
            .O(N__23378),
            .I(\c0.FRAME_MATCHER_i_0 ));
    CascadeMux I__3522 (
            .O(N__23367),
            .I(N__23363));
    CascadeMux I__3521 (
            .O(N__23366),
            .I(N__23357));
    InMux I__3520 (
            .O(N__23363),
            .I(N__23353));
    CascadeMux I__3519 (
            .O(N__23362),
            .I(N__23350));
    CascadeMux I__3518 (
            .O(N__23361),
            .I(N__23346));
    InMux I__3517 (
            .O(N__23360),
            .I(N__23343));
    InMux I__3516 (
            .O(N__23357),
            .I(N__23339));
    InMux I__3515 (
            .O(N__23356),
            .I(N__23332));
    LocalMux I__3514 (
            .O(N__23353),
            .I(N__23328));
    InMux I__3513 (
            .O(N__23350),
            .I(N__23325));
    CascadeMux I__3512 (
            .O(N__23349),
            .I(N__23322));
    InMux I__3511 (
            .O(N__23346),
            .I(N__23319));
    LocalMux I__3510 (
            .O(N__23343),
            .I(N__23316));
    CascadeMux I__3509 (
            .O(N__23342),
            .I(N__23313));
    LocalMux I__3508 (
            .O(N__23339),
            .I(N__23310));
    InMux I__3507 (
            .O(N__23338),
            .I(N__23305));
    InMux I__3506 (
            .O(N__23337),
            .I(N__23305));
    CascadeMux I__3505 (
            .O(N__23336),
            .I(N__23302));
    CascadeMux I__3504 (
            .O(N__23335),
            .I(N__23299));
    LocalMux I__3503 (
            .O(N__23332),
            .I(N__23296));
    CascadeMux I__3502 (
            .O(N__23331),
            .I(N__23291));
    Span4Mux_v I__3501 (
            .O(N__23328),
            .I(N__23285));
    LocalMux I__3500 (
            .O(N__23325),
            .I(N__23285));
    InMux I__3499 (
            .O(N__23322),
            .I(N__23282));
    LocalMux I__3498 (
            .O(N__23319),
            .I(N__23277));
    Span4Mux_v I__3497 (
            .O(N__23316),
            .I(N__23277));
    InMux I__3496 (
            .O(N__23313),
            .I(N__23274));
    Span4Mux_h I__3495 (
            .O(N__23310),
            .I(N__23269));
    LocalMux I__3494 (
            .O(N__23305),
            .I(N__23269));
    InMux I__3493 (
            .O(N__23302),
            .I(N__23266));
    InMux I__3492 (
            .O(N__23299),
            .I(N__23263));
    Span4Mux_h I__3491 (
            .O(N__23296),
            .I(N__23260));
    InMux I__3490 (
            .O(N__23295),
            .I(N__23251));
    InMux I__3489 (
            .O(N__23294),
            .I(N__23251));
    InMux I__3488 (
            .O(N__23291),
            .I(N__23251));
    InMux I__3487 (
            .O(N__23290),
            .I(N__23251));
    Span4Mux_v I__3486 (
            .O(N__23285),
            .I(N__23240));
    LocalMux I__3485 (
            .O(N__23282),
            .I(N__23240));
    Span4Mux_h I__3484 (
            .O(N__23277),
            .I(N__23240));
    LocalMux I__3483 (
            .O(N__23274),
            .I(N__23240));
    Span4Mux_v I__3482 (
            .O(N__23269),
            .I(N__23240));
    LocalMux I__3481 (
            .O(N__23266),
            .I(N__23231));
    LocalMux I__3480 (
            .O(N__23263),
            .I(N__23231));
    Sp12to4 I__3479 (
            .O(N__23260),
            .I(N__23231));
    LocalMux I__3478 (
            .O(N__23251),
            .I(N__23231));
    Odrv4 I__3477 (
            .O(N__23240),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv12 I__3476 (
            .O(N__23231),
            .I(\c0.FRAME_MATCHER_i_2 ));
    InMux I__3475 (
            .O(N__23226),
            .I(N__23223));
    LocalMux I__3474 (
            .O(N__23223),
            .I(N__23217));
    InMux I__3473 (
            .O(N__23222),
            .I(N__23214));
    InMux I__3472 (
            .O(N__23221),
            .I(N__23211));
    InMux I__3471 (
            .O(N__23220),
            .I(N__23207));
    Span4Mux_h I__3470 (
            .O(N__23217),
            .I(N__23200));
    LocalMux I__3469 (
            .O(N__23214),
            .I(N__23200));
    LocalMux I__3468 (
            .O(N__23211),
            .I(N__23200));
    InMux I__3467 (
            .O(N__23210),
            .I(N__23197));
    LocalMux I__3466 (
            .O(N__23207),
            .I(N__23194));
    Span4Mux_v I__3465 (
            .O(N__23200),
            .I(N__23187));
    LocalMux I__3464 (
            .O(N__23197),
            .I(N__23187));
    Span4Mux_v I__3463 (
            .O(N__23194),
            .I(N__23187));
    Odrv4 I__3462 (
            .O(N__23187),
            .I(\c0.rx.n12963 ));
    CascadeMux I__3461 (
            .O(N__23184),
            .I(n120_cascade_));
    InMux I__3460 (
            .O(N__23181),
            .I(N__23174));
    InMux I__3459 (
            .O(N__23180),
            .I(N__23174));
    InMux I__3458 (
            .O(N__23179),
            .I(N__23171));
    LocalMux I__3457 (
            .O(N__23174),
            .I(N__23168));
    LocalMux I__3456 (
            .O(N__23171),
            .I(data_in_frame_2_3));
    Odrv4 I__3455 (
            .O(N__23168),
            .I(data_in_frame_2_3));
    InMux I__3454 (
            .O(N__23163),
            .I(N__23160));
    LocalMux I__3453 (
            .O(N__23160),
            .I(N__23154));
    InMux I__3452 (
            .O(N__23159),
            .I(N__23151));
    InMux I__3451 (
            .O(N__23158),
            .I(N__23146));
    InMux I__3450 (
            .O(N__23157),
            .I(N__23146));
    Odrv4 I__3449 (
            .O(N__23154),
            .I(data_in_frame_0_4));
    LocalMux I__3448 (
            .O(N__23151),
            .I(data_in_frame_0_4));
    LocalMux I__3447 (
            .O(N__23146),
            .I(data_in_frame_0_4));
    CascadeMux I__3446 (
            .O(N__23139),
            .I(N__23136));
    InMux I__3445 (
            .O(N__23136),
            .I(N__23133));
    LocalMux I__3444 (
            .O(N__23133),
            .I(N__23127));
    InMux I__3443 (
            .O(N__23132),
            .I(N__23124));
    InMux I__3442 (
            .O(N__23131),
            .I(N__23121));
    InMux I__3441 (
            .O(N__23130),
            .I(N__23118));
    Odrv4 I__3440 (
            .O(N__23127),
            .I(data_in_frame_0_5));
    LocalMux I__3439 (
            .O(N__23124),
            .I(data_in_frame_0_5));
    LocalMux I__3438 (
            .O(N__23121),
            .I(data_in_frame_0_5));
    LocalMux I__3437 (
            .O(N__23118),
            .I(data_in_frame_0_5));
    InMux I__3436 (
            .O(N__23109),
            .I(N__23104));
    InMux I__3435 (
            .O(N__23108),
            .I(N__23101));
    InMux I__3434 (
            .O(N__23107),
            .I(N__23098));
    LocalMux I__3433 (
            .O(N__23104),
            .I(data_in_frame_2_6));
    LocalMux I__3432 (
            .O(N__23101),
            .I(data_in_frame_2_6));
    LocalMux I__3431 (
            .O(N__23098),
            .I(data_in_frame_2_6));
    InMux I__3430 (
            .O(N__23091),
            .I(N__23088));
    LocalMux I__3429 (
            .O(N__23088),
            .I(\c0.n15_adj_2416 ));
    InMux I__3428 (
            .O(N__23085),
            .I(N__23079));
    InMux I__3427 (
            .O(N__23084),
            .I(N__23076));
    InMux I__3426 (
            .O(N__23083),
            .I(N__23073));
    InMux I__3425 (
            .O(N__23082),
            .I(N__23070));
    LocalMux I__3424 (
            .O(N__23079),
            .I(\c0.n2138 ));
    LocalMux I__3423 (
            .O(N__23076),
            .I(\c0.n2138 ));
    LocalMux I__3422 (
            .O(N__23073),
            .I(\c0.n2138 ));
    LocalMux I__3421 (
            .O(N__23070),
            .I(\c0.n2138 ));
    InMux I__3420 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__3419 (
            .O(N__23058),
            .I(N__23055));
    Odrv4 I__3418 (
            .O(N__23055),
            .I(\c0.n22_adj_2419 ));
    InMux I__3417 (
            .O(N__23052),
            .I(N__23048));
    InMux I__3416 (
            .O(N__23051),
            .I(N__23045));
    LocalMux I__3415 (
            .O(N__23048),
            .I(data_in_frame_6_7));
    LocalMux I__3414 (
            .O(N__23045),
            .I(data_in_frame_6_7));
    InMux I__3413 (
            .O(N__23040),
            .I(N__23036));
    InMux I__3412 (
            .O(N__23039),
            .I(N__23033));
    LocalMux I__3411 (
            .O(N__23036),
            .I(\c0.n17813 ));
    LocalMux I__3410 (
            .O(N__23033),
            .I(\c0.n17813 ));
    InMux I__3409 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__3408 (
            .O(N__23025),
            .I(\c0.n10761 ));
    InMux I__3407 (
            .O(N__23022),
            .I(N__23013));
    InMux I__3406 (
            .O(N__23021),
            .I(N__23013));
    InMux I__3405 (
            .O(N__23020),
            .I(N__23013));
    LocalMux I__3404 (
            .O(N__23013),
            .I(N__23007));
    InMux I__3403 (
            .O(N__23012),
            .I(N__23002));
    InMux I__3402 (
            .O(N__23011),
            .I(N__23002));
    InMux I__3401 (
            .O(N__23010),
            .I(N__22999));
    Odrv4 I__3400 (
            .O(N__23007),
            .I(data_in_frame_0_0));
    LocalMux I__3399 (
            .O(N__23002),
            .I(data_in_frame_0_0));
    LocalMux I__3398 (
            .O(N__22999),
            .I(data_in_frame_0_0));
    CascadeMux I__3397 (
            .O(N__22992),
            .I(\c0.n10761_cascade_ ));
    InMux I__3396 (
            .O(N__22989),
            .I(N__22986));
    LocalMux I__3395 (
            .O(N__22986),
            .I(N__22982));
    CascadeMux I__3394 (
            .O(N__22985),
            .I(N__22978));
    Span4Mux_h I__3393 (
            .O(N__22982),
            .I(N__22973));
    InMux I__3392 (
            .O(N__22981),
            .I(N__22970));
    InMux I__3391 (
            .O(N__22978),
            .I(N__22965));
    InMux I__3390 (
            .O(N__22977),
            .I(N__22965));
    InMux I__3389 (
            .O(N__22976),
            .I(N__22962));
    Odrv4 I__3388 (
            .O(N__22973),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__3387 (
            .O(N__22970),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__3386 (
            .O(N__22965),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__3385 (
            .O(N__22962),
            .I(\c0.data_in_frame_1_5 ));
    CascadeMux I__3384 (
            .O(N__22953),
            .I(\c0.n17733_cascade_ ));
    InMux I__3383 (
            .O(N__22950),
            .I(N__22946));
    InMux I__3382 (
            .O(N__22949),
            .I(N__22943));
    LocalMux I__3381 (
            .O(N__22946),
            .I(data_in_frame_6_0));
    LocalMux I__3380 (
            .O(N__22943),
            .I(data_in_frame_6_0));
    InMux I__3379 (
            .O(N__22938),
            .I(N__22935));
    LocalMux I__3378 (
            .O(N__22935),
            .I(\c0.n17735 ));
    CascadeMux I__3377 (
            .O(N__22932),
            .I(N__22928));
    InMux I__3376 (
            .O(N__22931),
            .I(N__22923));
    InMux I__3375 (
            .O(N__22928),
            .I(N__22919));
    InMux I__3374 (
            .O(N__22927),
            .I(N__22914));
    InMux I__3373 (
            .O(N__22926),
            .I(N__22914));
    LocalMux I__3372 (
            .O(N__22923),
            .I(N__22911));
    InMux I__3371 (
            .O(N__22922),
            .I(N__22908));
    LocalMux I__3370 (
            .O(N__22919),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__3369 (
            .O(N__22914),
            .I(\c0.data_in_frame_1_6 ));
    Odrv4 I__3368 (
            .O(N__22911),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__3367 (
            .O(N__22908),
            .I(\c0.data_in_frame_1_6 ));
    InMux I__3366 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__3365 (
            .O(N__22896),
            .I(\c0.n17733 ));
    InMux I__3364 (
            .O(N__22893),
            .I(N__22890));
    LocalMux I__3363 (
            .O(N__22890),
            .I(\c0.n21_adj_2421 ));
    InMux I__3362 (
            .O(N__22887),
            .I(N__22884));
    LocalMux I__3361 (
            .O(N__22884),
            .I(N__22881));
    Span4Mux_h I__3360 (
            .O(N__22881),
            .I(N__22878));
    Odrv4 I__3359 (
            .O(N__22878),
            .I(\c0.n24_adj_2418 ));
    CascadeMux I__3358 (
            .O(N__22875),
            .I(\c0.n23_adj_2420_cascade_ ));
    CascadeMux I__3357 (
            .O(N__22872),
            .I(n16797_cascade_));
    InMux I__3356 (
            .O(N__22869),
            .I(N__22865));
    InMux I__3355 (
            .O(N__22868),
            .I(N__22862));
    LocalMux I__3354 (
            .O(N__22865),
            .I(N__22859));
    LocalMux I__3353 (
            .O(N__22862),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__3352 (
            .O(N__22859),
            .I(\c0.data_in_frame_3_5 ));
    CascadeMux I__3351 (
            .O(N__22854),
            .I(\c0.rx.n129_cascade_ ));
    InMux I__3350 (
            .O(N__22851),
            .I(N__22847));
    InMux I__3349 (
            .O(N__22850),
            .I(N__22844));
    LocalMux I__3348 (
            .O(N__22847),
            .I(N__22841));
    LocalMux I__3347 (
            .O(N__22844),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__3346 (
            .O(N__22841),
            .I(\c0.data_in_frame_3_7 ));
    CascadeMux I__3345 (
            .O(N__22836),
            .I(N__22832));
    InMux I__3344 (
            .O(N__22835),
            .I(N__22829));
    InMux I__3343 (
            .O(N__22832),
            .I(N__22826));
    LocalMux I__3342 (
            .O(N__22829),
            .I(data_in_frame_6_1));
    LocalMux I__3341 (
            .O(N__22826),
            .I(data_in_frame_6_1));
    InMux I__3340 (
            .O(N__22821),
            .I(N__22818));
    LocalMux I__3339 (
            .O(N__22818),
            .I(n18043));
    InMux I__3338 (
            .O(N__22815),
            .I(N__22812));
    LocalMux I__3337 (
            .O(N__22812),
            .I(n18044));
    IoInMux I__3336 (
            .O(N__22809),
            .I(N__22806));
    LocalMux I__3335 (
            .O(N__22806),
            .I(N__22803));
    Span12Mux_s8_v I__3334 (
            .O(N__22803),
            .I(N__22800));
    Odrv12 I__3333 (
            .O(N__22800),
            .I(LED_c));
    IoInMux I__3332 (
            .O(N__22797),
            .I(N__22794));
    LocalMux I__3331 (
            .O(N__22794),
            .I(N__22791));
    Span4Mux_s3_h I__3330 (
            .O(N__22791),
            .I(N__22788));
    Odrv4 I__3329 (
            .O(N__22788),
            .I(PIN_3_c_2));
    SRMux I__3328 (
            .O(N__22785),
            .I(N__22782));
    LocalMux I__3327 (
            .O(N__22782),
            .I(N__22779));
    Span4Mux_h I__3326 (
            .O(N__22779),
            .I(N__22776));
    Span4Mux_s1_v I__3325 (
            .O(N__22776),
            .I(N__22773));
    Odrv4 I__3324 (
            .O(N__22773),
            .I(\c0.n4_adj_2225 ));
    InMux I__3323 (
            .O(N__22770),
            .I(N__22766));
    IoInMux I__3322 (
            .O(N__22769),
            .I(N__22763));
    LocalMux I__3321 (
            .O(N__22766),
            .I(N__22760));
    LocalMux I__3320 (
            .O(N__22763),
            .I(N__22757));
    Span4Mux_s2_v I__3319 (
            .O(N__22760),
            .I(N__22754));
    Span4Mux_s2_v I__3318 (
            .O(N__22757),
            .I(N__22751));
    Span4Mux_v I__3317 (
            .O(N__22754),
            .I(N__22748));
    Span4Mux_v I__3316 (
            .O(N__22751),
            .I(N__22742));
    Span4Mux_v I__3315 (
            .O(N__22748),
            .I(N__22742));
    InMux I__3314 (
            .O(N__22747),
            .I(N__22739));
    Odrv4 I__3313 (
            .O(N__22742),
            .I(tx2_o));
    LocalMux I__3312 (
            .O(N__22739),
            .I(tx2_o));
    IoInMux I__3311 (
            .O(N__22734),
            .I(N__22731));
    LocalMux I__3310 (
            .O(N__22731),
            .I(N__22728));
    Span4Mux_s1_v I__3309 (
            .O(N__22728),
            .I(N__22725));
    Odrv4 I__3308 (
            .O(N__22725),
            .I(tx2_enable));
    SRMux I__3307 (
            .O(N__22722),
            .I(N__22719));
    LocalMux I__3306 (
            .O(N__22719),
            .I(N__22716));
    Span4Mux_h I__3305 (
            .O(N__22716),
            .I(N__22713));
    Span4Mux_s2_h I__3304 (
            .O(N__22713),
            .I(N__22710));
    Odrv4 I__3303 (
            .O(N__22710),
            .I(\c0.n4_adj_2216 ));
    InMux I__3302 (
            .O(N__22707),
            .I(N__22703));
    InMux I__3301 (
            .O(N__22706),
            .I(N__22700));
    LocalMux I__3300 (
            .O(N__22703),
            .I(N__22697));
    LocalMux I__3299 (
            .O(N__22700),
            .I(\c0.data_in_frame_3_3 ));
    Odrv4 I__3298 (
            .O(N__22697),
            .I(\c0.data_in_frame_3_3 ));
    InMux I__3297 (
            .O(N__22692),
            .I(N__22688));
    CascadeMux I__3296 (
            .O(N__22691),
            .I(N__22685));
    LocalMux I__3295 (
            .O(N__22688),
            .I(N__22681));
    InMux I__3294 (
            .O(N__22685),
            .I(N__22678));
    InMux I__3293 (
            .O(N__22684),
            .I(N__22675));
    Span4Mux_v I__3292 (
            .O(N__22681),
            .I(N__22672));
    LocalMux I__3291 (
            .O(N__22678),
            .I(N__22669));
    LocalMux I__3290 (
            .O(N__22675),
            .I(data_in_frame_2_2));
    Odrv4 I__3289 (
            .O(N__22672),
            .I(data_in_frame_2_2));
    Odrv12 I__3288 (
            .O(N__22669),
            .I(data_in_frame_2_2));
    InMux I__3287 (
            .O(N__22662),
            .I(N__22659));
    LocalMux I__3286 (
            .O(N__22659),
            .I(\c0.n18_adj_2417 ));
    CascadeMux I__3285 (
            .O(N__22656),
            .I(N__22653));
    InMux I__3284 (
            .O(N__22653),
            .I(N__22649));
    CascadeMux I__3283 (
            .O(N__22652),
            .I(N__22646));
    LocalMux I__3282 (
            .O(N__22649),
            .I(N__22642));
    InMux I__3281 (
            .O(N__22646),
            .I(N__22639));
    InMux I__3280 (
            .O(N__22645),
            .I(N__22636));
    Span4Mux_h I__3279 (
            .O(N__22642),
            .I(N__22631));
    LocalMux I__3278 (
            .O(N__22639),
            .I(N__22631));
    LocalMux I__3277 (
            .O(N__22636),
            .I(data_in_frame_2_1));
    Odrv4 I__3276 (
            .O(N__22631),
            .I(data_in_frame_2_1));
    CascadeMux I__3275 (
            .O(N__22626),
            .I(N__22623));
    InMux I__3274 (
            .O(N__22623),
            .I(N__22620));
    LocalMux I__3273 (
            .O(N__22620),
            .I(N__22614));
    InMux I__3272 (
            .O(N__22619),
            .I(N__22611));
    InMux I__3271 (
            .O(N__22618),
            .I(N__22608));
    InMux I__3270 (
            .O(N__22617),
            .I(N__22605));
    Span4Mux_h I__3269 (
            .O(N__22614),
            .I(N__22602));
    LocalMux I__3268 (
            .O(N__22611),
            .I(N__22595));
    LocalMux I__3267 (
            .O(N__22608),
            .I(N__22595));
    LocalMux I__3266 (
            .O(N__22605),
            .I(N__22595));
    Span4Mux_s0_h I__3265 (
            .O(N__22602),
            .I(N__22592));
    Span4Mux_v I__3264 (
            .O(N__22595),
            .I(N__22589));
    Odrv4 I__3263 (
            .O(N__22592),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv4 I__3262 (
            .O(N__22589),
            .I(\c0.FRAME_MATCHER_i_12 ));
    InMux I__3261 (
            .O(N__22584),
            .I(N__22581));
    LocalMux I__3260 (
            .O(N__22581),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_12 ));
    InMux I__3259 (
            .O(N__22578),
            .I(N__22575));
    LocalMux I__3258 (
            .O(N__22575),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_27 ));
    InMux I__3257 (
            .O(N__22572),
            .I(N__22556));
    InMux I__3256 (
            .O(N__22571),
            .I(N__22556));
    InMux I__3255 (
            .O(N__22570),
            .I(N__22547));
    InMux I__3254 (
            .O(N__22569),
            .I(N__22547));
    InMux I__3253 (
            .O(N__22568),
            .I(N__22547));
    InMux I__3252 (
            .O(N__22567),
            .I(N__22547));
    InMux I__3251 (
            .O(N__22566),
            .I(N__22544));
    InMux I__3250 (
            .O(N__22565),
            .I(N__22533));
    InMux I__3249 (
            .O(N__22564),
            .I(N__22533));
    InMux I__3248 (
            .O(N__22563),
            .I(N__22533));
    InMux I__3247 (
            .O(N__22562),
            .I(N__22533));
    InMux I__3246 (
            .O(N__22561),
            .I(N__22533));
    LocalMux I__3245 (
            .O(N__22556),
            .I(N__22525));
    LocalMux I__3244 (
            .O(N__22547),
            .I(N__22522));
    LocalMux I__3243 (
            .O(N__22544),
            .I(N__22519));
    LocalMux I__3242 (
            .O(N__22533),
            .I(N__22516));
    InMux I__3241 (
            .O(N__22532),
            .I(N__22505));
    InMux I__3240 (
            .O(N__22531),
            .I(N__22505));
    InMux I__3239 (
            .O(N__22530),
            .I(N__22505));
    InMux I__3238 (
            .O(N__22529),
            .I(N__22505));
    InMux I__3237 (
            .O(N__22528),
            .I(N__22505));
    Span4Mux_v I__3236 (
            .O(N__22525),
            .I(N__22488));
    Span4Mux_v I__3235 (
            .O(N__22522),
            .I(N__22488));
    Span4Mux_h I__3234 (
            .O(N__22519),
            .I(N__22481));
    Span4Mux_v I__3233 (
            .O(N__22516),
            .I(N__22481));
    LocalMux I__3232 (
            .O(N__22505),
            .I(N__22481));
    InMux I__3231 (
            .O(N__22504),
            .I(N__22472));
    InMux I__3230 (
            .O(N__22503),
            .I(N__22472));
    InMux I__3229 (
            .O(N__22502),
            .I(N__22472));
    InMux I__3228 (
            .O(N__22501),
            .I(N__22472));
    InMux I__3227 (
            .O(N__22500),
            .I(N__22463));
    InMux I__3226 (
            .O(N__22499),
            .I(N__22463));
    InMux I__3225 (
            .O(N__22498),
            .I(N__22463));
    InMux I__3224 (
            .O(N__22497),
            .I(N__22463));
    InMux I__3223 (
            .O(N__22496),
            .I(N__22460));
    InMux I__3222 (
            .O(N__22495),
            .I(N__22453));
    InMux I__3221 (
            .O(N__22494),
            .I(N__22453));
    InMux I__3220 (
            .O(N__22493),
            .I(N__22453));
    Odrv4 I__3219 (
            .O(N__22488),
            .I(\c0.n13033 ));
    Odrv4 I__3218 (
            .O(N__22481),
            .I(\c0.n13033 ));
    LocalMux I__3217 (
            .O(N__22472),
            .I(\c0.n13033 ));
    LocalMux I__3216 (
            .O(N__22463),
            .I(\c0.n13033 ));
    LocalMux I__3215 (
            .O(N__22460),
            .I(\c0.n13033 ));
    LocalMux I__3214 (
            .O(N__22453),
            .I(\c0.n13033 ));
    InMux I__3213 (
            .O(N__22440),
            .I(N__22435));
    InMux I__3212 (
            .O(N__22439),
            .I(N__22431));
    InMux I__3211 (
            .O(N__22438),
            .I(N__22428));
    LocalMux I__3210 (
            .O(N__22435),
            .I(N__22425));
    InMux I__3209 (
            .O(N__22434),
            .I(N__22422));
    LocalMux I__3208 (
            .O(N__22431),
            .I(N__22419));
    LocalMux I__3207 (
            .O(N__22428),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__3206 (
            .O(N__22425),
            .I(\c0.FRAME_MATCHER_i_26 ));
    LocalMux I__3205 (
            .O(N__22422),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__3204 (
            .O(N__22419),
            .I(\c0.FRAME_MATCHER_i_26 ));
    InMux I__3203 (
            .O(N__22410),
            .I(N__22407));
    LocalMux I__3202 (
            .O(N__22407),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_26 ));
    InMux I__3201 (
            .O(N__22404),
            .I(N__22401));
    LocalMux I__3200 (
            .O(N__22401),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_27 ));
    CascadeMux I__3199 (
            .O(N__22398),
            .I(N__22394));
    InMux I__3198 (
            .O(N__22397),
            .I(N__22391));
    InMux I__3197 (
            .O(N__22394),
            .I(N__22388));
    LocalMux I__3196 (
            .O(N__22391),
            .I(N__22385));
    LocalMux I__3195 (
            .O(N__22388),
            .I(N__22378));
    Span4Mux_v I__3194 (
            .O(N__22385),
            .I(N__22378));
    InMux I__3193 (
            .O(N__22384),
            .I(N__22373));
    InMux I__3192 (
            .O(N__22383),
            .I(N__22373));
    Odrv4 I__3191 (
            .O(N__22378),
            .I(\c0.FRAME_MATCHER_i_27 ));
    LocalMux I__3190 (
            .O(N__22373),
            .I(\c0.FRAME_MATCHER_i_27 ));
    SRMux I__3189 (
            .O(N__22368),
            .I(N__22365));
    LocalMux I__3188 (
            .O(N__22365),
            .I(N__22362));
    Span4Mux_h I__3187 (
            .O(N__22362),
            .I(N__22359));
    Odrv4 I__3186 (
            .O(N__22359),
            .I(\c0.n3_adj_2287 ));
    InMux I__3185 (
            .O(N__22356),
            .I(N__22353));
    LocalMux I__3184 (
            .O(N__22353),
            .I(N__22350));
    Span4Mux_v I__3183 (
            .O(N__22350),
            .I(N__22347));
    Odrv4 I__3182 (
            .O(N__22347),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_3 ));
    InMux I__3181 (
            .O(N__22344),
            .I(N__22340));
    CascadeMux I__3180 (
            .O(N__22343),
            .I(N__22337));
    LocalMux I__3179 (
            .O(N__22340),
            .I(N__22332));
    InMux I__3178 (
            .O(N__22337),
            .I(N__22329));
    InMux I__3177 (
            .O(N__22336),
            .I(N__22326));
    InMux I__3176 (
            .O(N__22335),
            .I(N__22323));
    Span4Mux_h I__3175 (
            .O(N__22332),
            .I(N__22320));
    LocalMux I__3174 (
            .O(N__22329),
            .I(N__22313));
    LocalMux I__3173 (
            .O(N__22326),
            .I(N__22313));
    LocalMux I__3172 (
            .O(N__22323),
            .I(N__22313));
    Odrv4 I__3171 (
            .O(N__22320),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__3170 (
            .O(N__22313),
            .I(\c0.FRAME_MATCHER_i_3 ));
    SRMux I__3169 (
            .O(N__22308),
            .I(N__22305));
    LocalMux I__3168 (
            .O(N__22305),
            .I(N__22302));
    Span4Mux_v I__3167 (
            .O(N__22302),
            .I(N__22299));
    Odrv4 I__3166 (
            .O(N__22299),
            .I(\c0.n3_adj_2340 ));
    InMux I__3165 (
            .O(N__22296),
            .I(N__22293));
    LocalMux I__3164 (
            .O(N__22293),
            .I(N__22290));
    Odrv4 I__3163 (
            .O(N__22290),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_28 ));
    CascadeMux I__3162 (
            .O(N__22287),
            .I(N__22284));
    InMux I__3161 (
            .O(N__22284),
            .I(N__22279));
    CascadeMux I__3160 (
            .O(N__22283),
            .I(N__22276));
    InMux I__3159 (
            .O(N__22282),
            .I(N__22272));
    LocalMux I__3158 (
            .O(N__22279),
            .I(N__22269));
    InMux I__3157 (
            .O(N__22276),
            .I(N__22266));
    InMux I__3156 (
            .O(N__22275),
            .I(N__22263));
    LocalMux I__3155 (
            .O(N__22272),
            .I(N__22260));
    Span4Mux_h I__3154 (
            .O(N__22269),
            .I(N__22253));
    LocalMux I__3153 (
            .O(N__22266),
            .I(N__22253));
    LocalMux I__3152 (
            .O(N__22263),
            .I(N__22253));
    Odrv12 I__3151 (
            .O(N__22260),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__3150 (
            .O(N__22253),
            .I(\c0.FRAME_MATCHER_i_28 ));
    SRMux I__3149 (
            .O(N__22248),
            .I(N__22245));
    LocalMux I__3148 (
            .O(N__22245),
            .I(N__22242));
    Span4Mux_h I__3147 (
            .O(N__22242),
            .I(N__22239));
    Span4Mux_v I__3146 (
            .O(N__22239),
            .I(N__22236));
    Odrv4 I__3145 (
            .O(N__22236),
            .I(\c0.n3_adj_2285 ));
    InMux I__3144 (
            .O(N__22233),
            .I(N__22230));
    LocalMux I__3143 (
            .O(N__22230),
            .I(N__22227));
    Odrv4 I__3142 (
            .O(N__22227),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_13 ));
    InMux I__3141 (
            .O(N__22224),
            .I(N__22218));
    InMux I__3140 (
            .O(N__22223),
            .I(N__22215));
    InMux I__3139 (
            .O(N__22222),
            .I(N__22212));
    InMux I__3138 (
            .O(N__22221),
            .I(N__22209));
    LocalMux I__3137 (
            .O(N__22218),
            .I(N__22204));
    LocalMux I__3136 (
            .O(N__22215),
            .I(N__22204));
    LocalMux I__3135 (
            .O(N__22212),
            .I(N__22201));
    LocalMux I__3134 (
            .O(N__22209),
            .I(N__22196));
    Span4Mux_h I__3133 (
            .O(N__22204),
            .I(N__22196));
    Span4Mux_s2_h I__3132 (
            .O(N__22201),
            .I(N__22193));
    Odrv4 I__3131 (
            .O(N__22196),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv4 I__3130 (
            .O(N__22193),
            .I(\c0.FRAME_MATCHER_i_10 ));
    InMux I__3129 (
            .O(N__22188),
            .I(N__22185));
    LocalMux I__3128 (
            .O(N__22185),
            .I(N__22182));
    Odrv4 I__3127 (
            .O(N__22182),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_10 ));
    CascadeMux I__3126 (
            .O(N__22179),
            .I(N__22175));
    InMux I__3125 (
            .O(N__22178),
            .I(N__22172));
    InMux I__3124 (
            .O(N__22175),
            .I(N__22169));
    LocalMux I__3123 (
            .O(N__22172),
            .I(N__22165));
    LocalMux I__3122 (
            .O(N__22169),
            .I(N__22162));
    InMux I__3121 (
            .O(N__22168),
            .I(N__22159));
    Span4Mux_h I__3120 (
            .O(N__22165),
            .I(N__22153));
    Span4Mux_v I__3119 (
            .O(N__22162),
            .I(N__22153));
    LocalMux I__3118 (
            .O(N__22159),
            .I(N__22150));
    InMux I__3117 (
            .O(N__22158),
            .I(N__22147));
    Span4Mux_v I__3116 (
            .O(N__22153),
            .I(N__22144));
    Span4Mux_h I__3115 (
            .O(N__22150),
            .I(N__22141));
    LocalMux I__3114 (
            .O(N__22147),
            .I(N__22138));
    Span4Mux_s1_h I__3113 (
            .O(N__22144),
            .I(N__22135));
    Odrv4 I__3112 (
            .O(N__22141),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv12 I__3111 (
            .O(N__22138),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv4 I__3110 (
            .O(N__22135),
            .I(\c0.FRAME_MATCHER_i_6 ));
    InMux I__3109 (
            .O(N__22128),
            .I(N__22125));
    LocalMux I__3108 (
            .O(N__22125),
            .I(N__22122));
    Span4Mux_h I__3107 (
            .O(N__22122),
            .I(N__22119));
    Odrv4 I__3106 (
            .O(N__22119),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_6 ));
    InMux I__3105 (
            .O(N__22116),
            .I(N__22113));
    LocalMux I__3104 (
            .O(N__22113),
            .I(N__22110));
    Span4Mux_h I__3103 (
            .O(N__22110),
            .I(N__22107));
    Odrv4 I__3102 (
            .O(N__22107),
            .I(\c0.n109 ));
    InMux I__3101 (
            .O(N__22104),
            .I(N__22101));
    LocalMux I__3100 (
            .O(N__22101),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_11 ));
    SRMux I__3099 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__3098 (
            .O(N__22095),
            .I(N__22092));
    Span4Mux_h I__3097 (
            .O(N__22092),
            .I(N__22089));
    Odrv4 I__3096 (
            .O(N__22089),
            .I(\c0.n3_adj_2324 ));
    CascadeMux I__3095 (
            .O(N__22086),
            .I(\c0.n26_adj_2379_cascade_ ));
    InMux I__3094 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__3093 (
            .O(N__22080),
            .I(N__22077));
    Span12Mux_s4_h I__3092 (
            .O(N__22077),
            .I(N__22074));
    Odrv12 I__3091 (
            .O(N__22074),
            .I(\c0.n44_adj_2382 ));
    CascadeMux I__3090 (
            .O(N__22071),
            .I(N__22067));
    CascadeMux I__3089 (
            .O(N__22070),
            .I(N__22064));
    InMux I__3088 (
            .O(N__22067),
            .I(N__22061));
    InMux I__3087 (
            .O(N__22064),
            .I(N__22058));
    LocalMux I__3086 (
            .O(N__22061),
            .I(N__22053));
    LocalMux I__3085 (
            .O(N__22058),
            .I(N__22050));
    InMux I__3084 (
            .O(N__22057),
            .I(N__22045));
    InMux I__3083 (
            .O(N__22056),
            .I(N__22045));
    Odrv12 I__3082 (
            .O(N__22053),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv4 I__3081 (
            .O(N__22050),
            .I(\c0.FRAME_MATCHER_i_11 ));
    LocalMux I__3080 (
            .O(N__22045),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__3079 (
            .O(N__22038),
            .I(N__22035));
    LocalMux I__3078 (
            .O(N__22035),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_11 ));
    CascadeMux I__3077 (
            .O(N__22032),
            .I(N__22029));
    InMux I__3076 (
            .O(N__22029),
            .I(N__22023));
    InMux I__3075 (
            .O(N__22028),
            .I(N__22018));
    InMux I__3074 (
            .O(N__22027),
            .I(N__22018));
    CascadeMux I__3073 (
            .O(N__22026),
            .I(N__22015));
    LocalMux I__3072 (
            .O(N__22023),
            .I(N__22010));
    LocalMux I__3071 (
            .O(N__22018),
            .I(N__22010));
    InMux I__3070 (
            .O(N__22015),
            .I(N__22007));
    Span4Mux_v I__3069 (
            .O(N__22010),
            .I(N__22004));
    LocalMux I__3068 (
            .O(N__22007),
            .I(\c0.FRAME_MATCHER_i_20 ));
    Odrv4 I__3067 (
            .O(N__22004),
            .I(\c0.FRAME_MATCHER_i_20 ));
    InMux I__3066 (
            .O(N__21999),
            .I(N__21996));
    LocalMux I__3065 (
            .O(N__21996),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_20 ));
    InMux I__3064 (
            .O(N__21993),
            .I(N__21990));
    LocalMux I__3063 (
            .O(N__21990),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_5 ));
    SRMux I__3062 (
            .O(N__21987),
            .I(N__21984));
    LocalMux I__3061 (
            .O(N__21984),
            .I(N__21981));
    Odrv4 I__3060 (
            .O(N__21981),
            .I(\c0.n3_adj_2336 ));
    CascadeMux I__3059 (
            .O(N__21978),
            .I(N__21975));
    InMux I__3058 (
            .O(N__21975),
            .I(N__21972));
    LocalMux I__3057 (
            .O(N__21972),
            .I(N__21966));
    InMux I__3056 (
            .O(N__21971),
            .I(N__21963));
    InMux I__3055 (
            .O(N__21970),
            .I(N__21958));
    InMux I__3054 (
            .O(N__21969),
            .I(N__21958));
    Odrv4 I__3053 (
            .O(N__21966),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__3052 (
            .O(N__21963),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__3051 (
            .O(N__21958),
            .I(\c0.FRAME_MATCHER_i_5 ));
    InMux I__3050 (
            .O(N__21951),
            .I(N__21948));
    LocalMux I__3049 (
            .O(N__21948),
            .I(N__21944));
    InMux I__3048 (
            .O(N__21947),
            .I(N__21941));
    Span4Mux_h I__3047 (
            .O(N__21944),
            .I(N__21938));
    LocalMux I__3046 (
            .O(N__21941),
            .I(N__21935));
    Odrv4 I__3045 (
            .O(N__21938),
            .I(\c0.n10_adj_2378 ));
    Odrv12 I__3044 (
            .O(N__21935),
            .I(\c0.n10_adj_2378 ));
    InMux I__3043 (
            .O(N__21930),
            .I(N__21927));
    LocalMux I__3042 (
            .O(N__21927),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_4 ));
    CascadeMux I__3041 (
            .O(N__21924),
            .I(N__21908));
    CascadeMux I__3040 (
            .O(N__21923),
            .I(N__21905));
    CascadeMux I__3039 (
            .O(N__21922),
            .I(N__21899));
    CascadeMux I__3038 (
            .O(N__21921),
            .I(N__21894));
    CascadeMux I__3037 (
            .O(N__21920),
            .I(N__21891));
    CascadeMux I__3036 (
            .O(N__21919),
            .I(N__21888));
    InMux I__3035 (
            .O(N__21918),
            .I(N__21876));
    InMux I__3034 (
            .O(N__21917),
            .I(N__21876));
    InMux I__3033 (
            .O(N__21916),
            .I(N__21871));
    InMux I__3032 (
            .O(N__21915),
            .I(N__21871));
    InMux I__3031 (
            .O(N__21914),
            .I(N__21863));
    InMux I__3030 (
            .O(N__21913),
            .I(N__21863));
    InMux I__3029 (
            .O(N__21912),
            .I(N__21863));
    InMux I__3028 (
            .O(N__21911),
            .I(N__21860));
    InMux I__3027 (
            .O(N__21908),
            .I(N__21847));
    InMux I__3026 (
            .O(N__21905),
            .I(N__21847));
    InMux I__3025 (
            .O(N__21904),
            .I(N__21847));
    InMux I__3024 (
            .O(N__21903),
            .I(N__21847));
    InMux I__3023 (
            .O(N__21902),
            .I(N__21847));
    InMux I__3022 (
            .O(N__21899),
            .I(N__21847));
    InMux I__3021 (
            .O(N__21898),
            .I(N__21834));
    InMux I__3020 (
            .O(N__21897),
            .I(N__21834));
    InMux I__3019 (
            .O(N__21894),
            .I(N__21834));
    InMux I__3018 (
            .O(N__21891),
            .I(N__21834));
    InMux I__3017 (
            .O(N__21888),
            .I(N__21834));
    InMux I__3016 (
            .O(N__21887),
            .I(N__21834));
    InMux I__3015 (
            .O(N__21886),
            .I(N__21821));
    InMux I__3014 (
            .O(N__21885),
            .I(N__21821));
    InMux I__3013 (
            .O(N__21884),
            .I(N__21821));
    InMux I__3012 (
            .O(N__21883),
            .I(N__21821));
    InMux I__3011 (
            .O(N__21882),
            .I(N__21821));
    InMux I__3010 (
            .O(N__21881),
            .I(N__21821));
    LocalMux I__3009 (
            .O(N__21876),
            .I(N__21818));
    LocalMux I__3008 (
            .O(N__21871),
            .I(N__21815));
    CascadeMux I__3007 (
            .O(N__21870),
            .I(N__21807));
    LocalMux I__3006 (
            .O(N__21863),
            .I(N__21802));
    LocalMux I__3005 (
            .O(N__21860),
            .I(N__21802));
    LocalMux I__3004 (
            .O(N__21847),
            .I(N__21797));
    LocalMux I__3003 (
            .O(N__21834),
            .I(N__21797));
    LocalMux I__3002 (
            .O(N__21821),
            .I(N__21794));
    Span4Mux_h I__3001 (
            .O(N__21818),
            .I(N__21789));
    Span4Mux_h I__3000 (
            .O(N__21815),
            .I(N__21789));
    InMux I__2999 (
            .O(N__21814),
            .I(N__21781));
    InMux I__2998 (
            .O(N__21813),
            .I(N__21781));
    InMux I__2997 (
            .O(N__21812),
            .I(N__21781));
    InMux I__2996 (
            .O(N__21811),
            .I(N__21774));
    InMux I__2995 (
            .O(N__21810),
            .I(N__21774));
    InMux I__2994 (
            .O(N__21807),
            .I(N__21774));
    Span12Mux_v I__2993 (
            .O(N__21802),
            .I(N__21771));
    Span4Mux_h I__2992 (
            .O(N__21797),
            .I(N__21768));
    Span4Mux_h I__2991 (
            .O(N__21794),
            .I(N__21763));
    Span4Mux_v I__2990 (
            .O(N__21789),
            .I(N__21763));
    InMux I__2989 (
            .O(N__21788),
            .I(N__21760));
    LocalMux I__2988 (
            .O(N__21781),
            .I(\c0.n7199 ));
    LocalMux I__2987 (
            .O(N__21774),
            .I(\c0.n7199 ));
    Odrv12 I__2986 (
            .O(N__21771),
            .I(\c0.n7199 ));
    Odrv4 I__2985 (
            .O(N__21768),
            .I(\c0.n7199 ));
    Odrv4 I__2984 (
            .O(N__21763),
            .I(\c0.n7199 ));
    LocalMux I__2983 (
            .O(N__21760),
            .I(\c0.n7199 ));
    InMux I__2982 (
            .O(N__21747),
            .I(N__21742));
    InMux I__2981 (
            .O(N__21746),
            .I(N__21739));
    CascadeMux I__2980 (
            .O(N__21745),
            .I(N__21736));
    LocalMux I__2979 (
            .O(N__21742),
            .I(N__21730));
    LocalMux I__2978 (
            .O(N__21739),
            .I(N__21730));
    InMux I__2977 (
            .O(N__21736),
            .I(N__21725));
    InMux I__2976 (
            .O(N__21735),
            .I(N__21725));
    Sp12to4 I__2975 (
            .O(N__21730),
            .I(N__21720));
    LocalMux I__2974 (
            .O(N__21725),
            .I(N__21720));
    Odrv12 I__2973 (
            .O(N__21720),
            .I(\c0.FRAME_MATCHER_i_4 ));
    CascadeMux I__2972 (
            .O(N__21717),
            .I(N__21705));
    CascadeMux I__2971 (
            .O(N__21716),
            .I(N__21702));
    CascadeMux I__2970 (
            .O(N__21715),
            .I(N__21692));
    CascadeMux I__2969 (
            .O(N__21714),
            .I(N__21689));
    CascadeMux I__2968 (
            .O(N__21713),
            .I(N__21686));
    InMux I__2967 (
            .O(N__21712),
            .I(N__21679));
    InMux I__2966 (
            .O(N__21711),
            .I(N__21679));
    CascadeMux I__2965 (
            .O(N__21710),
            .I(N__21675));
    CascadeMux I__2964 (
            .O(N__21709),
            .I(N__21672));
    CascadeMux I__2963 (
            .O(N__21708),
            .I(N__21666));
    InMux I__2962 (
            .O(N__21705),
            .I(N__21656));
    InMux I__2961 (
            .O(N__21702),
            .I(N__21656));
    InMux I__2960 (
            .O(N__21701),
            .I(N__21656));
    CascadeMux I__2959 (
            .O(N__21700),
            .I(N__21653));
    CascadeMux I__2958 (
            .O(N__21699),
            .I(N__21650));
    InMux I__2957 (
            .O(N__21698),
            .I(N__21643));
    CascadeMux I__2956 (
            .O(N__21697),
            .I(N__21640));
    CascadeMux I__2955 (
            .O(N__21696),
            .I(N__21636));
    InMux I__2954 (
            .O(N__21695),
            .I(N__21623));
    InMux I__2953 (
            .O(N__21692),
            .I(N__21623));
    InMux I__2952 (
            .O(N__21689),
            .I(N__21623));
    InMux I__2951 (
            .O(N__21686),
            .I(N__21623));
    InMux I__2950 (
            .O(N__21685),
            .I(N__21623));
    InMux I__2949 (
            .O(N__21684),
            .I(N__21623));
    LocalMux I__2948 (
            .O(N__21679),
            .I(N__21620));
    InMux I__2947 (
            .O(N__21678),
            .I(N__21611));
    InMux I__2946 (
            .O(N__21675),
            .I(N__21611));
    InMux I__2945 (
            .O(N__21672),
            .I(N__21611));
    InMux I__2944 (
            .O(N__21671),
            .I(N__21611));
    InMux I__2943 (
            .O(N__21670),
            .I(N__21598));
    InMux I__2942 (
            .O(N__21669),
            .I(N__21598));
    InMux I__2941 (
            .O(N__21666),
            .I(N__21598));
    InMux I__2940 (
            .O(N__21665),
            .I(N__21598));
    InMux I__2939 (
            .O(N__21664),
            .I(N__21598));
    InMux I__2938 (
            .O(N__21663),
            .I(N__21598));
    LocalMux I__2937 (
            .O(N__21656),
            .I(N__21595));
    InMux I__2936 (
            .O(N__21653),
            .I(N__21582));
    InMux I__2935 (
            .O(N__21650),
            .I(N__21582));
    InMux I__2934 (
            .O(N__21649),
            .I(N__21582));
    InMux I__2933 (
            .O(N__21648),
            .I(N__21582));
    InMux I__2932 (
            .O(N__21647),
            .I(N__21582));
    InMux I__2931 (
            .O(N__21646),
            .I(N__21582));
    LocalMux I__2930 (
            .O(N__21643),
            .I(N__21579));
    InMux I__2929 (
            .O(N__21640),
            .I(N__21572));
    InMux I__2928 (
            .O(N__21639),
            .I(N__21572));
    InMux I__2927 (
            .O(N__21636),
            .I(N__21572));
    LocalMux I__2926 (
            .O(N__21623),
            .I(N__21567));
    Span4Mux_v I__2925 (
            .O(N__21620),
            .I(N__21567));
    LocalMux I__2924 (
            .O(N__21611),
            .I(\c0.n10353 ));
    LocalMux I__2923 (
            .O(N__21598),
            .I(\c0.n10353 ));
    Odrv4 I__2922 (
            .O(N__21595),
            .I(\c0.n10353 ));
    LocalMux I__2921 (
            .O(N__21582),
            .I(\c0.n10353 ));
    Odrv12 I__2920 (
            .O(N__21579),
            .I(\c0.n10353 ));
    LocalMux I__2919 (
            .O(N__21572),
            .I(\c0.n10353 ));
    Odrv4 I__2918 (
            .O(N__21567),
            .I(\c0.n10353 ));
    SRMux I__2917 (
            .O(N__21552),
            .I(N__21549));
    LocalMux I__2916 (
            .O(N__21549),
            .I(N__21546));
    Odrv12 I__2915 (
            .O(N__21546),
            .I(\c0.n3_adj_2338 ));
    CascadeMux I__2914 (
            .O(N__21543),
            .I(N__21539));
    InMux I__2913 (
            .O(N__21542),
            .I(N__21536));
    InMux I__2912 (
            .O(N__21539),
            .I(N__21532));
    LocalMux I__2911 (
            .O(N__21536),
            .I(N__21512));
    InMux I__2910 (
            .O(N__21535),
            .I(N__21500));
    LocalMux I__2909 (
            .O(N__21532),
            .I(N__21497));
    InMux I__2908 (
            .O(N__21531),
            .I(N__21486));
    InMux I__2907 (
            .O(N__21530),
            .I(N__21486));
    InMux I__2906 (
            .O(N__21529),
            .I(N__21486));
    InMux I__2905 (
            .O(N__21528),
            .I(N__21486));
    InMux I__2904 (
            .O(N__21527),
            .I(N__21486));
    InMux I__2903 (
            .O(N__21526),
            .I(N__21473));
    InMux I__2902 (
            .O(N__21525),
            .I(N__21473));
    InMux I__2901 (
            .O(N__21524),
            .I(N__21473));
    InMux I__2900 (
            .O(N__21523),
            .I(N__21473));
    InMux I__2899 (
            .O(N__21522),
            .I(N__21473));
    InMux I__2898 (
            .O(N__21521),
            .I(N__21473));
    InMux I__2897 (
            .O(N__21520),
            .I(N__21460));
    InMux I__2896 (
            .O(N__21519),
            .I(N__21460));
    InMux I__2895 (
            .O(N__21518),
            .I(N__21460));
    InMux I__2894 (
            .O(N__21517),
            .I(N__21460));
    InMux I__2893 (
            .O(N__21516),
            .I(N__21460));
    InMux I__2892 (
            .O(N__21515),
            .I(N__21460));
    Span4Mux_h I__2891 (
            .O(N__21512),
            .I(N__21457));
    InMux I__2890 (
            .O(N__21511),
            .I(N__21439));
    InMux I__2889 (
            .O(N__21510),
            .I(N__21439));
    InMux I__2888 (
            .O(N__21509),
            .I(N__21439));
    InMux I__2887 (
            .O(N__21508),
            .I(N__21439));
    InMux I__2886 (
            .O(N__21507),
            .I(N__21436));
    InMux I__2885 (
            .O(N__21506),
            .I(N__21427));
    InMux I__2884 (
            .O(N__21505),
            .I(N__21427));
    InMux I__2883 (
            .O(N__21504),
            .I(N__21427));
    InMux I__2882 (
            .O(N__21503),
            .I(N__21427));
    LocalMux I__2881 (
            .O(N__21500),
            .I(N__21424));
    Span4Mux_s2_h I__2880 (
            .O(N__21497),
            .I(N__21412));
    LocalMux I__2879 (
            .O(N__21486),
            .I(N__21412));
    LocalMux I__2878 (
            .O(N__21473),
            .I(N__21412));
    LocalMux I__2877 (
            .O(N__21460),
            .I(N__21412));
    Span4Mux_v I__2876 (
            .O(N__21457),
            .I(N__21409));
    InMux I__2875 (
            .O(N__21456),
            .I(N__21402));
    InMux I__2874 (
            .O(N__21455),
            .I(N__21402));
    InMux I__2873 (
            .O(N__21454),
            .I(N__21402));
    InMux I__2872 (
            .O(N__21453),
            .I(N__21399));
    InMux I__2871 (
            .O(N__21452),
            .I(N__21385));
    InMux I__2870 (
            .O(N__21451),
            .I(N__21385));
    InMux I__2869 (
            .O(N__21450),
            .I(N__21385));
    InMux I__2868 (
            .O(N__21449),
            .I(N__21385));
    InMux I__2867 (
            .O(N__21448),
            .I(N__21385));
    LocalMux I__2866 (
            .O(N__21439),
            .I(N__21382));
    LocalMux I__2865 (
            .O(N__21436),
            .I(N__21379));
    LocalMux I__2864 (
            .O(N__21427),
            .I(N__21376));
    Span4Mux_v I__2863 (
            .O(N__21424),
            .I(N__21367));
    InMux I__2862 (
            .O(N__21423),
            .I(N__21360));
    InMux I__2861 (
            .O(N__21422),
            .I(N__21360));
    InMux I__2860 (
            .O(N__21421),
            .I(N__21360));
    Span4Mux_v I__2859 (
            .O(N__21412),
            .I(N__21357));
    Span4Mux_v I__2858 (
            .O(N__21409),
            .I(N__21354));
    LocalMux I__2857 (
            .O(N__21402),
            .I(N__21349));
    LocalMux I__2856 (
            .O(N__21399),
            .I(N__21349));
    InMux I__2855 (
            .O(N__21398),
            .I(N__21342));
    InMux I__2854 (
            .O(N__21397),
            .I(N__21342));
    InMux I__2853 (
            .O(N__21396),
            .I(N__21342));
    LocalMux I__2852 (
            .O(N__21385),
            .I(N__21335));
    Span4Mux_h I__2851 (
            .O(N__21382),
            .I(N__21335));
    Span4Mux_h I__2850 (
            .O(N__21379),
            .I(N__21335));
    Span4Mux_h I__2849 (
            .O(N__21376),
            .I(N__21332));
    InMux I__2848 (
            .O(N__21375),
            .I(N__21323));
    InMux I__2847 (
            .O(N__21374),
            .I(N__21323));
    InMux I__2846 (
            .O(N__21373),
            .I(N__21323));
    InMux I__2845 (
            .O(N__21372),
            .I(N__21323));
    InMux I__2844 (
            .O(N__21371),
            .I(N__21318));
    InMux I__2843 (
            .O(N__21370),
            .I(N__21318));
    Odrv4 I__2842 (
            .O(N__21367),
            .I(n63));
    LocalMux I__2841 (
            .O(N__21360),
            .I(n63));
    Odrv4 I__2840 (
            .O(N__21357),
            .I(n63));
    Odrv4 I__2839 (
            .O(N__21354),
            .I(n63));
    Odrv12 I__2838 (
            .O(N__21349),
            .I(n63));
    LocalMux I__2837 (
            .O(N__21342),
            .I(n63));
    Odrv4 I__2836 (
            .O(N__21335),
            .I(n63));
    Odrv4 I__2835 (
            .O(N__21332),
            .I(n63));
    LocalMux I__2834 (
            .O(N__21323),
            .I(n63));
    LocalMux I__2833 (
            .O(N__21318),
            .I(n63));
    InMux I__2832 (
            .O(N__21297),
            .I(N__21292));
    InMux I__2831 (
            .O(N__21296),
            .I(N__21286));
    InMux I__2830 (
            .O(N__21295),
            .I(N__21283));
    LocalMux I__2829 (
            .O(N__21292),
            .I(N__21280));
    InMux I__2828 (
            .O(N__21291),
            .I(N__21277));
    CascadeMux I__2827 (
            .O(N__21290),
            .I(N__21273));
    CascadeMux I__2826 (
            .O(N__21289),
            .I(N__21268));
    LocalMux I__2825 (
            .O(N__21286),
            .I(N__21265));
    LocalMux I__2824 (
            .O(N__21283),
            .I(N__21262));
    Span4Mux_h I__2823 (
            .O(N__21280),
            .I(N__21259));
    LocalMux I__2822 (
            .O(N__21277),
            .I(N__21256));
    InMux I__2821 (
            .O(N__21276),
            .I(N__21247));
    InMux I__2820 (
            .O(N__21273),
            .I(N__21247));
    InMux I__2819 (
            .O(N__21272),
            .I(N__21244));
    InMux I__2818 (
            .O(N__21271),
            .I(N__21239));
    InMux I__2817 (
            .O(N__21268),
            .I(N__21239));
    Span4Mux_v I__2816 (
            .O(N__21265),
            .I(N__21234));
    Span4Mux_v I__2815 (
            .O(N__21262),
            .I(N__21234));
    Span4Mux_v I__2814 (
            .O(N__21259),
            .I(N__21229));
    Span4Mux_h I__2813 (
            .O(N__21256),
            .I(N__21229));
    InMux I__2812 (
            .O(N__21255),
            .I(N__21224));
    InMux I__2811 (
            .O(N__21254),
            .I(N__21224));
    InMux I__2810 (
            .O(N__21253),
            .I(N__21219));
    InMux I__2809 (
            .O(N__21252),
            .I(N__21219));
    LocalMux I__2808 (
            .O(N__21247),
            .I(\c0.n63_adj_2262 ));
    LocalMux I__2807 (
            .O(N__21244),
            .I(\c0.n63_adj_2262 ));
    LocalMux I__2806 (
            .O(N__21239),
            .I(\c0.n63_adj_2262 ));
    Odrv4 I__2805 (
            .O(N__21234),
            .I(\c0.n63_adj_2262 ));
    Odrv4 I__2804 (
            .O(N__21229),
            .I(\c0.n63_adj_2262 ));
    LocalMux I__2803 (
            .O(N__21224),
            .I(\c0.n63_adj_2262 ));
    LocalMux I__2802 (
            .O(N__21219),
            .I(\c0.n63_adj_2262 ));
    InMux I__2801 (
            .O(N__21204),
            .I(N__21198));
    InMux I__2800 (
            .O(N__21203),
            .I(N__21198));
    LocalMux I__2799 (
            .O(N__21198),
            .I(N__21192));
    InMux I__2798 (
            .O(N__21197),
            .I(N__21189));
    InMux I__2797 (
            .O(N__21196),
            .I(N__21186));
    InMux I__2796 (
            .O(N__21195),
            .I(N__21183));
    Span4Mux_v I__2795 (
            .O(N__21192),
            .I(N__21178));
    LocalMux I__2794 (
            .O(N__21189),
            .I(N__21178));
    LocalMux I__2793 (
            .O(N__21186),
            .I(N__21175));
    LocalMux I__2792 (
            .O(N__21183),
            .I(N__21170));
    Span4Mux_h I__2791 (
            .O(N__21178),
            .I(N__21158));
    Span4Mux_h I__2790 (
            .O(N__21175),
            .I(N__21158));
    InMux I__2789 (
            .O(N__21174),
            .I(N__21153));
    InMux I__2788 (
            .O(N__21173),
            .I(N__21153));
    Span4Mux_h I__2787 (
            .O(N__21170),
            .I(N__21150));
    InMux I__2786 (
            .O(N__21169),
            .I(N__21147));
    InMux I__2785 (
            .O(N__21168),
            .I(N__21140));
    InMux I__2784 (
            .O(N__21167),
            .I(N__21140));
    InMux I__2783 (
            .O(N__21166),
            .I(N__21140));
    InMux I__2782 (
            .O(N__21165),
            .I(N__21137));
    InMux I__2781 (
            .O(N__21164),
            .I(N__21132));
    InMux I__2780 (
            .O(N__21163),
            .I(N__21132));
    Odrv4 I__2779 (
            .O(N__21158),
            .I(n63_adj_2534));
    LocalMux I__2778 (
            .O(N__21153),
            .I(n63_adj_2534));
    Odrv4 I__2777 (
            .O(N__21150),
            .I(n63_adj_2534));
    LocalMux I__2776 (
            .O(N__21147),
            .I(n63_adj_2534));
    LocalMux I__2775 (
            .O(N__21140),
            .I(n63_adj_2534));
    LocalMux I__2774 (
            .O(N__21137),
            .I(n63_adj_2534));
    LocalMux I__2773 (
            .O(N__21132),
            .I(n63_adj_2534));
    InMux I__2772 (
            .O(N__21117),
            .I(N__21114));
    LocalMux I__2771 (
            .O(N__21114),
            .I(N__21111));
    Odrv4 I__2770 (
            .O(N__21111),
            .I(\c0.n113 ));
    CascadeMux I__2769 (
            .O(N__21108),
            .I(N__21105));
    InMux I__2768 (
            .O(N__21105),
            .I(N__21100));
    InMux I__2767 (
            .O(N__21104),
            .I(N__21097));
    InMux I__2766 (
            .O(N__21103),
            .I(N__21094));
    LocalMux I__2765 (
            .O(N__21100),
            .I(N__21090));
    LocalMux I__2764 (
            .O(N__21097),
            .I(N__21085));
    LocalMux I__2763 (
            .O(N__21094),
            .I(N__21085));
    InMux I__2762 (
            .O(N__21093),
            .I(N__21082));
    Span4Mux_h I__2761 (
            .O(N__21090),
            .I(N__21077));
    Span4Mux_h I__2760 (
            .O(N__21085),
            .I(N__21077));
    LocalMux I__2759 (
            .O(N__21082),
            .I(N__21074));
    Odrv4 I__2758 (
            .O(N__21077),
            .I(\c0.FRAME_MATCHER_i_14 ));
    Odrv12 I__2757 (
            .O(N__21074),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__2756 (
            .O(N__21069),
            .I(N__21066));
    LocalMux I__2755 (
            .O(N__21066),
            .I(N__21063));
    Odrv4 I__2754 (
            .O(N__21063),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_14 ));
    InMux I__2753 (
            .O(N__21060),
            .I(N__21057));
    LocalMux I__2752 (
            .O(N__21057),
            .I(N__21054));
    Span4Mux_v I__2751 (
            .O(N__21054),
            .I(N__21051));
    Odrv4 I__2750 (
            .O(N__21051),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_28 ));
    CascadeMux I__2749 (
            .O(N__21048),
            .I(N__21043));
    InMux I__2748 (
            .O(N__21047),
            .I(N__21040));
    CascadeMux I__2747 (
            .O(N__21046),
            .I(N__21037));
    InMux I__2746 (
            .O(N__21043),
            .I(N__21033));
    LocalMux I__2745 (
            .O(N__21040),
            .I(N__21030));
    InMux I__2744 (
            .O(N__21037),
            .I(N__21027));
    CascadeMux I__2743 (
            .O(N__21036),
            .I(N__21024));
    LocalMux I__2742 (
            .O(N__21033),
            .I(N__21021));
    Span4Mux_h I__2741 (
            .O(N__21030),
            .I(N__21018));
    LocalMux I__2740 (
            .O(N__21027),
            .I(N__21015));
    InMux I__2739 (
            .O(N__21024),
            .I(N__21012));
    Span4Mux_h I__2738 (
            .O(N__21021),
            .I(N__21009));
    Span4Mux_v I__2737 (
            .O(N__21018),
            .I(N__21004));
    Span4Mux_v I__2736 (
            .O(N__21015),
            .I(N__21004));
    LocalMux I__2735 (
            .O(N__21012),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__2734 (
            .O(N__21009),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__2733 (
            .O(N__21004),
            .I(\c0.FRAME_MATCHER_i_19 ));
    InMux I__2732 (
            .O(N__20997),
            .I(N__20994));
    LocalMux I__2731 (
            .O(N__20994),
            .I(N__20991));
    Span4Mux_v I__2730 (
            .O(N__20991),
            .I(N__20988));
    Odrv4 I__2729 (
            .O(N__20988),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_19 ));
    CascadeMux I__2728 (
            .O(N__20985),
            .I(N__20978));
    InMux I__2727 (
            .O(N__20984),
            .I(N__20972));
    InMux I__2726 (
            .O(N__20983),
            .I(N__20965));
    InMux I__2725 (
            .O(N__20982),
            .I(N__20965));
    InMux I__2724 (
            .O(N__20981),
            .I(N__20965));
    InMux I__2723 (
            .O(N__20978),
            .I(N__20962));
    InMux I__2722 (
            .O(N__20977),
            .I(N__20959));
    InMux I__2721 (
            .O(N__20976),
            .I(N__20956));
    CascadeMux I__2720 (
            .O(N__20975),
            .I(N__20953));
    LocalMux I__2719 (
            .O(N__20972),
            .I(N__20946));
    LocalMux I__2718 (
            .O(N__20965),
            .I(N__20943));
    LocalMux I__2717 (
            .O(N__20962),
            .I(N__20936));
    LocalMux I__2716 (
            .O(N__20959),
            .I(N__20936));
    LocalMux I__2715 (
            .O(N__20956),
            .I(N__20936));
    InMux I__2714 (
            .O(N__20953),
            .I(N__20927));
    InMux I__2713 (
            .O(N__20952),
            .I(N__20927));
    InMux I__2712 (
            .O(N__20951),
            .I(N__20927));
    InMux I__2711 (
            .O(N__20950),
            .I(N__20927));
    InMux I__2710 (
            .O(N__20949),
            .I(N__20924));
    Span4Mux_h I__2709 (
            .O(N__20946),
            .I(N__20921));
    Span4Mux_s2_h I__2708 (
            .O(N__20943),
            .I(N__20914));
    Span4Mux_h I__2707 (
            .O(N__20936),
            .I(N__20914));
    LocalMux I__2706 (
            .O(N__20927),
            .I(N__20914));
    LocalMux I__2705 (
            .O(N__20924),
            .I(N__20911));
    Span4Mux_v I__2704 (
            .O(N__20921),
            .I(N__20908));
    Span4Mux_v I__2703 (
            .O(N__20914),
            .I(N__20905));
    Odrv4 I__2702 (
            .O(N__20911),
            .I(FRAME_MATCHER_i_31));
    Odrv4 I__2701 (
            .O(N__20908),
            .I(FRAME_MATCHER_i_31));
    Odrv4 I__2700 (
            .O(N__20905),
            .I(FRAME_MATCHER_i_31));
    CascadeMux I__2699 (
            .O(N__20898),
            .I(N__20895));
    InMux I__2698 (
            .O(N__20895),
            .I(N__20892));
    LocalMux I__2697 (
            .O(N__20892),
            .I(N__20889));
    Span4Mux_v I__2696 (
            .O(N__20889),
            .I(N__20886));
    Odrv4 I__2695 (
            .O(N__20886),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_31 ));
    CascadeMux I__2694 (
            .O(N__20883),
            .I(n63_adj_2534_cascade_));
    InMux I__2693 (
            .O(N__20880),
            .I(N__20877));
    LocalMux I__2692 (
            .O(N__20877),
            .I(N__20874));
    Odrv4 I__2691 (
            .O(N__20874),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_18 ));
    CascadeMux I__2690 (
            .O(N__20871),
            .I(\c0.n63_adj_2262_cascade_ ));
    InMux I__2689 (
            .O(N__20868),
            .I(N__20865));
    LocalMux I__2688 (
            .O(N__20865),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_5 ));
    CascadeMux I__2687 (
            .O(N__20862),
            .I(n11058_cascade_));
    InMux I__2686 (
            .O(N__20859),
            .I(N__20856));
    LocalMux I__2685 (
            .O(N__20856),
            .I(N__20853));
    Span4Mux_v I__2684 (
            .O(N__20853),
            .I(N__20850));
    Odrv4 I__2683 (
            .O(N__20850),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_3 ));
    InMux I__2682 (
            .O(N__20847),
            .I(N__20844));
    LocalMux I__2681 (
            .O(N__20844),
            .I(N__20840));
    InMux I__2680 (
            .O(N__20843),
            .I(N__20837));
    Span4Mux_h I__2679 (
            .O(N__20840),
            .I(N__20833));
    LocalMux I__2678 (
            .O(N__20837),
            .I(N__20830));
    InMux I__2677 (
            .O(N__20836),
            .I(N__20827));
    Odrv4 I__2676 (
            .O(N__20833),
            .I(\c0.n1502 ));
    Odrv4 I__2675 (
            .O(N__20830),
            .I(\c0.n1502 ));
    LocalMux I__2674 (
            .O(N__20827),
            .I(\c0.n1502 ));
    CascadeMux I__2673 (
            .O(N__20820),
            .I(\c0.n1502_cascade_ ));
    InMux I__2672 (
            .O(N__20817),
            .I(N__20811));
    InMux I__2671 (
            .O(N__20816),
            .I(N__20808));
    InMux I__2670 (
            .O(N__20815),
            .I(N__20803));
    InMux I__2669 (
            .O(N__20814),
            .I(N__20803));
    LocalMux I__2668 (
            .O(N__20811),
            .I(N__20798));
    LocalMux I__2667 (
            .O(N__20808),
            .I(N__20798));
    LocalMux I__2666 (
            .O(N__20803),
            .I(N__20792));
    Span4Mux_v I__2665 (
            .O(N__20798),
            .I(N__20789));
    InMux I__2664 (
            .O(N__20797),
            .I(N__20782));
    InMux I__2663 (
            .O(N__20796),
            .I(N__20782));
    InMux I__2662 (
            .O(N__20795),
            .I(N__20782));
    Odrv4 I__2661 (
            .O(N__20792),
            .I(\c0.n10522 ));
    Odrv4 I__2660 (
            .O(N__20789),
            .I(\c0.n10522 ));
    LocalMux I__2659 (
            .O(N__20782),
            .I(\c0.n10522 ));
    InMux I__2658 (
            .O(N__20775),
            .I(N__20772));
    LocalMux I__2657 (
            .O(N__20772),
            .I(\c0.n4_adj_2266 ));
    CascadeMux I__2656 (
            .O(N__20769),
            .I(\c0.n13033_cascade_ ));
    InMux I__2655 (
            .O(N__20766),
            .I(N__20762));
    InMux I__2654 (
            .O(N__20765),
            .I(N__20759));
    LocalMux I__2653 (
            .O(N__20762),
            .I(N__20756));
    LocalMux I__2652 (
            .O(N__20759),
            .I(N__20753));
    Span4Mux_v I__2651 (
            .O(N__20756),
            .I(N__20748));
    Span4Mux_h I__2650 (
            .O(N__20753),
            .I(N__20745));
    InMux I__2649 (
            .O(N__20752),
            .I(N__20740));
    InMux I__2648 (
            .O(N__20751),
            .I(N__20740));
    Odrv4 I__2647 (
            .O(N__20748),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__2646 (
            .O(N__20745),
            .I(\c0.FRAME_MATCHER_i_30 ));
    LocalMux I__2645 (
            .O(N__20740),
            .I(\c0.FRAME_MATCHER_i_30 ));
    InMux I__2644 (
            .O(N__20733),
            .I(N__20730));
    LocalMux I__2643 (
            .O(N__20730),
            .I(N__20727));
    Span4Mux_v I__2642 (
            .O(N__20727),
            .I(N__20724));
    Odrv4 I__2641 (
            .O(N__20724),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_30 ));
    InMux I__2640 (
            .O(N__20721),
            .I(N__20718));
    LocalMux I__2639 (
            .O(N__20718),
            .I(N__20713));
    CascadeMux I__2638 (
            .O(N__20717),
            .I(N__20709));
    InMux I__2637 (
            .O(N__20716),
            .I(N__20706));
    Span4Mux_v I__2636 (
            .O(N__20713),
            .I(N__20703));
    InMux I__2635 (
            .O(N__20712),
            .I(N__20698));
    InMux I__2634 (
            .O(N__20709),
            .I(N__20698));
    LocalMux I__2633 (
            .O(N__20706),
            .I(N__20695));
    Span4Mux_v I__2632 (
            .O(N__20703),
            .I(N__20692));
    LocalMux I__2631 (
            .O(N__20698),
            .I(N__20689));
    Odrv12 I__2630 (
            .O(N__20695),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__2629 (
            .O(N__20692),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__2628 (
            .O(N__20689),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__2627 (
            .O(N__20682),
            .I(N__20679));
    LocalMux I__2626 (
            .O(N__20679),
            .I(N__20676));
    Span4Mux_v I__2625 (
            .O(N__20676),
            .I(N__20673));
    Odrv4 I__2624 (
            .O(N__20673),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_29 ));
    CascadeMux I__2623 (
            .O(N__20670),
            .I(n16802_cascade_));
    CascadeMux I__2622 (
            .O(N__20667),
            .I(\c0.n10569_cascade_ ));
    InMux I__2621 (
            .O(N__20664),
            .I(N__20655));
    InMux I__2620 (
            .O(N__20663),
            .I(N__20655));
    InMux I__2619 (
            .O(N__20662),
            .I(N__20655));
    LocalMux I__2618 (
            .O(N__20655),
            .I(N__20650));
    InMux I__2617 (
            .O(N__20654),
            .I(N__20645));
    InMux I__2616 (
            .O(N__20653),
            .I(N__20645));
    Odrv12 I__2615 (
            .O(N__20650),
            .I(data_in_frame_0_1));
    LocalMux I__2614 (
            .O(N__20645),
            .I(data_in_frame_0_1));
    InMux I__2613 (
            .O(N__20640),
            .I(N__20637));
    LocalMux I__2612 (
            .O(N__20637),
            .I(N__20634));
    Span4Mux_h I__2611 (
            .O(N__20634),
            .I(N__20631));
    Span4Mux_v I__2610 (
            .O(N__20631),
            .I(N__20628));
    Odrv4 I__2609 (
            .O(N__20628),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__2608 (
            .O(N__20625),
            .I(N__20621));
    CascadeMux I__2607 (
            .O(N__20624),
            .I(N__20618));
    InMux I__2606 (
            .O(N__20621),
            .I(N__20615));
    InMux I__2605 (
            .O(N__20618),
            .I(N__20612));
    LocalMux I__2604 (
            .O(N__20615),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__2603 (
            .O(N__20612),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__2602 (
            .O(N__20607),
            .I(N__20603));
    InMux I__2601 (
            .O(N__20606),
            .I(N__20600));
    LocalMux I__2600 (
            .O(N__20603),
            .I(\c0.n2137_adj_2237 ));
    LocalMux I__2599 (
            .O(N__20600),
            .I(\c0.n2137_adj_2237 ));
    CascadeMux I__2598 (
            .O(N__20595),
            .I(\c0.n2137_adj_2237_cascade_ ));
    CascadeMux I__2597 (
            .O(N__20592),
            .I(N__20587));
    InMux I__2596 (
            .O(N__20591),
            .I(N__20584));
    InMux I__2595 (
            .O(N__20590),
            .I(N__20579));
    InMux I__2594 (
            .O(N__20587),
            .I(N__20579));
    LocalMux I__2593 (
            .O(N__20584),
            .I(data_in_frame_2_0));
    LocalMux I__2592 (
            .O(N__20579),
            .I(data_in_frame_2_0));
    InMux I__2591 (
            .O(N__20574),
            .I(N__20569));
    CascadeMux I__2590 (
            .O(N__20573),
            .I(N__20566));
    InMux I__2589 (
            .O(N__20572),
            .I(N__20563));
    LocalMux I__2588 (
            .O(N__20569),
            .I(N__20560));
    InMux I__2587 (
            .O(N__20566),
            .I(N__20557));
    LocalMux I__2586 (
            .O(N__20563),
            .I(data_in_frame_2_5));
    Odrv4 I__2585 (
            .O(N__20560),
            .I(data_in_frame_2_5));
    LocalMux I__2584 (
            .O(N__20557),
            .I(data_in_frame_2_5));
    CascadeMux I__2583 (
            .O(N__20550),
            .I(N__20547));
    InMux I__2582 (
            .O(N__20547),
            .I(N__20543));
    InMux I__2581 (
            .O(N__20546),
            .I(N__20540));
    LocalMux I__2580 (
            .O(N__20543),
            .I(N__20537));
    LocalMux I__2579 (
            .O(N__20540),
            .I(data_in_frame_5_6));
    Odrv4 I__2578 (
            .O(N__20537),
            .I(data_in_frame_5_6));
    CascadeMux I__2577 (
            .O(N__20532),
            .I(N__20528));
    InMux I__2576 (
            .O(N__20531),
            .I(N__20523));
    InMux I__2575 (
            .O(N__20528),
            .I(N__20523));
    LocalMux I__2574 (
            .O(N__20523),
            .I(\c0.data_in_frame_3_0 ));
    InMux I__2573 (
            .O(N__20520),
            .I(N__20516));
    InMux I__2572 (
            .O(N__20519),
            .I(N__20513));
    LocalMux I__2571 (
            .O(N__20516),
            .I(\c0.n2126 ));
    LocalMux I__2570 (
            .O(N__20513),
            .I(\c0.n2126 ));
    SRMux I__2569 (
            .O(N__20508),
            .I(N__20505));
    LocalMux I__2568 (
            .O(N__20505),
            .I(N__20502));
    Odrv4 I__2567 (
            .O(N__20502),
            .I(\c0.n8_adj_2249 ));
    InMux I__2566 (
            .O(N__20499),
            .I(N__20492));
    CascadeMux I__2565 (
            .O(N__20498),
            .I(N__20488));
    InMux I__2564 (
            .O(N__20497),
            .I(N__20485));
    InMux I__2563 (
            .O(N__20496),
            .I(N__20482));
    InMux I__2562 (
            .O(N__20495),
            .I(N__20479));
    LocalMux I__2561 (
            .O(N__20492),
            .I(N__20476));
    InMux I__2560 (
            .O(N__20491),
            .I(N__20473));
    InMux I__2559 (
            .O(N__20488),
            .I(N__20470));
    LocalMux I__2558 (
            .O(N__20485),
            .I(N__20465));
    LocalMux I__2557 (
            .O(N__20482),
            .I(N__20465));
    LocalMux I__2556 (
            .O(N__20479),
            .I(N__20462));
    Span4Mux_h I__2555 (
            .O(N__20476),
            .I(N__20457));
    LocalMux I__2554 (
            .O(N__20473),
            .I(N__20457));
    LocalMux I__2553 (
            .O(N__20470),
            .I(N__20454));
    Span4Mux_h I__2552 (
            .O(N__20465),
            .I(N__20449));
    Span4Mux_s0_v I__2551 (
            .O(N__20462),
            .I(N__20449));
    Span4Mux_h I__2550 (
            .O(N__20457),
            .I(N__20446));
    Span4Mux_v I__2549 (
            .O(N__20454),
            .I(N__20443));
    Odrv4 I__2548 (
            .O(N__20449),
            .I(\c0.n4_adj_2349 ));
    Odrv4 I__2547 (
            .O(N__20446),
            .I(\c0.n4_adj_2349 ));
    Odrv4 I__2546 (
            .O(N__20443),
            .I(\c0.n4_adj_2349 ));
    SRMux I__2545 (
            .O(N__20436),
            .I(N__20433));
    LocalMux I__2544 (
            .O(N__20433),
            .I(N__20430));
    Span4Mux_h I__2543 (
            .O(N__20430),
            .I(N__20427));
    Odrv4 I__2542 (
            .O(N__20427),
            .I(\c0.n8_adj_2244 ));
    InMux I__2541 (
            .O(N__20424),
            .I(N__20419));
    InMux I__2540 (
            .O(N__20423),
            .I(N__20416));
    InMux I__2539 (
            .O(N__20422),
            .I(N__20413));
    LocalMux I__2538 (
            .O(N__20419),
            .I(\c0.FRAME_MATCHER_state_20 ));
    LocalMux I__2537 (
            .O(N__20416),
            .I(\c0.FRAME_MATCHER_state_20 ));
    LocalMux I__2536 (
            .O(N__20413),
            .I(\c0.FRAME_MATCHER_state_20 ));
    CascadeMux I__2535 (
            .O(N__20406),
            .I(N__20403));
    InMux I__2534 (
            .O(N__20403),
            .I(N__20400));
    LocalMux I__2533 (
            .O(N__20400),
            .I(N__20397));
    Span4Mux_h I__2532 (
            .O(N__20397),
            .I(N__20392));
    InMux I__2531 (
            .O(N__20396),
            .I(N__20387));
    InMux I__2530 (
            .O(N__20395),
            .I(N__20387));
    Odrv4 I__2529 (
            .O(N__20392),
            .I(\c0.FRAME_MATCHER_state_29 ));
    LocalMux I__2528 (
            .O(N__20387),
            .I(\c0.FRAME_MATCHER_state_29 ));
    CascadeMux I__2527 (
            .O(N__20382),
            .I(N__20379));
    InMux I__2526 (
            .O(N__20379),
            .I(N__20375));
    InMux I__2525 (
            .O(N__20378),
            .I(N__20372));
    LocalMux I__2524 (
            .O(N__20375),
            .I(N__20368));
    LocalMux I__2523 (
            .O(N__20372),
            .I(N__20365));
    InMux I__2522 (
            .O(N__20371),
            .I(N__20362));
    Span4Mux_h I__2521 (
            .O(N__20368),
            .I(N__20359));
    Span4Mux_h I__2520 (
            .O(N__20365),
            .I(N__20356));
    LocalMux I__2519 (
            .O(N__20362),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__2518 (
            .O(N__20359),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__2517 (
            .O(N__20356),
            .I(\c0.FRAME_MATCHER_state_5 ));
    InMux I__2516 (
            .O(N__20349),
            .I(N__20346));
    LocalMux I__2515 (
            .O(N__20346),
            .I(N__20343));
    Span4Mux_h I__2514 (
            .O(N__20343),
            .I(N__20338));
    InMux I__2513 (
            .O(N__20342),
            .I(N__20335));
    InMux I__2512 (
            .O(N__20341),
            .I(N__20332));
    Sp12to4 I__2511 (
            .O(N__20338),
            .I(N__20327));
    LocalMux I__2510 (
            .O(N__20335),
            .I(N__20327));
    LocalMux I__2509 (
            .O(N__20332),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv12 I__2508 (
            .O(N__20327),
            .I(\c0.FRAME_MATCHER_state_16 ));
    CascadeMux I__2507 (
            .O(N__20322),
            .I(\c0.n30_adj_2355_cascade_ ));
    InMux I__2506 (
            .O(N__20319),
            .I(N__20315));
    InMux I__2505 (
            .O(N__20318),
            .I(N__20312));
    LocalMux I__2504 (
            .O(N__20315),
            .I(N__20309));
    LocalMux I__2503 (
            .O(N__20312),
            .I(N__20305));
    Span4Mux_v I__2502 (
            .O(N__20309),
            .I(N__20302));
    InMux I__2501 (
            .O(N__20308),
            .I(N__20299));
    Span4Mux_v I__2500 (
            .O(N__20305),
            .I(N__20296));
    Span4Mux_s0_v I__2499 (
            .O(N__20302),
            .I(N__20293));
    LocalMux I__2498 (
            .O(N__20299),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__2497 (
            .O(N__20296),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__2496 (
            .O(N__20293),
            .I(\c0.FRAME_MATCHER_state_4 ));
    InMux I__2495 (
            .O(N__20286),
            .I(N__20283));
    LocalMux I__2494 (
            .O(N__20283),
            .I(\c0.n51 ));
    CascadeMux I__2493 (
            .O(N__20280),
            .I(\c0.n10613_cascade_ ));
    InMux I__2492 (
            .O(N__20277),
            .I(N__20274));
    LocalMux I__2491 (
            .O(N__20274),
            .I(\c0.n22_adj_2346 ));
    InMux I__2490 (
            .O(N__20271),
            .I(N__20268));
    LocalMux I__2489 (
            .O(N__20268),
            .I(N__20265));
    Span4Mux_s3_h I__2488 (
            .O(N__20265),
            .I(N__20262));
    Odrv4 I__2487 (
            .O(N__20262),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_30 ));
    InMux I__2486 (
            .O(N__20259),
            .I(\c0.n16515 ));
    InMux I__2485 (
            .O(N__20256),
            .I(\c0.n16516 ));
    InMux I__2484 (
            .O(N__20253),
            .I(N__20250));
    LocalMux I__2483 (
            .O(N__20250),
            .I(N__20247));
    Odrv4 I__2482 (
            .O(N__20247),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_31 ));
    InMux I__2481 (
            .O(N__20244),
            .I(N__20241));
    LocalMux I__2480 (
            .O(N__20241),
            .I(N__20238));
    Odrv12 I__2479 (
            .O(N__20238),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_9 ));
    CascadeMux I__2478 (
            .O(N__20235),
            .I(N__20230));
    InMux I__2477 (
            .O(N__20234),
            .I(N__20224));
    InMux I__2476 (
            .O(N__20233),
            .I(N__20224));
    InMux I__2475 (
            .O(N__20230),
            .I(N__20221));
    InMux I__2474 (
            .O(N__20229),
            .I(N__20218));
    LocalMux I__2473 (
            .O(N__20224),
            .I(N__20213));
    LocalMux I__2472 (
            .O(N__20221),
            .I(N__20213));
    LocalMux I__2471 (
            .O(N__20218),
            .I(N__20210));
    Span4Mux_v I__2470 (
            .O(N__20213),
            .I(N__20207));
    Span4Mux_s3_h I__2469 (
            .O(N__20210),
            .I(N__20204));
    Odrv4 I__2468 (
            .O(N__20207),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv4 I__2467 (
            .O(N__20204),
            .I(\c0.FRAME_MATCHER_i_9 ));
    SRMux I__2466 (
            .O(N__20199),
            .I(N__20196));
    LocalMux I__2465 (
            .O(N__20196),
            .I(N__20193));
    Span4Mux_v I__2464 (
            .O(N__20193),
            .I(N__20190));
    Span4Mux_v I__2463 (
            .O(N__20190),
            .I(N__20187));
    Odrv4 I__2462 (
            .O(N__20187),
            .I(\c0.n3_adj_2328 ));
    InMux I__2461 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__2460 (
            .O(N__20181),
            .I(N__20178));
    Odrv12 I__2459 (
            .O(N__20178),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_6 ));
    SRMux I__2458 (
            .O(N__20175),
            .I(N__20172));
    LocalMux I__2457 (
            .O(N__20172),
            .I(N__20169));
    Span4Mux_v I__2456 (
            .O(N__20169),
            .I(N__20166));
    Odrv4 I__2455 (
            .O(N__20166),
            .I(\c0.n3_adj_2334 ));
    CEMux I__2454 (
            .O(N__20163),
            .I(N__20160));
    LocalMux I__2453 (
            .O(N__20160),
            .I(N__20157));
    Span4Mux_v I__2452 (
            .O(N__20157),
            .I(N__20154));
    Odrv4 I__2451 (
            .O(N__20154),
            .I(\control.n18909 ));
    SRMux I__2450 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__2449 (
            .O(N__20148),
            .I(N__20145));
    Span4Mux_s1_v I__2448 (
            .O(N__20145),
            .I(N__20142));
    Span4Mux_h I__2447 (
            .O(N__20142),
            .I(N__20139));
    Odrv4 I__2446 (
            .O(N__20139),
            .I(\c0.n8_adj_2254 ));
    InMux I__2445 (
            .O(N__20136),
            .I(N__20133));
    LocalMux I__2444 (
            .O(N__20133),
            .I(N__20129));
    InMux I__2443 (
            .O(N__20132),
            .I(N__20126));
    Span4Mux_s3_v I__2442 (
            .O(N__20129),
            .I(N__20120));
    LocalMux I__2441 (
            .O(N__20126),
            .I(N__20120));
    InMux I__2440 (
            .O(N__20125),
            .I(N__20117));
    Span4Mux_h I__2439 (
            .O(N__20120),
            .I(N__20114));
    LocalMux I__2438 (
            .O(N__20117),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv4 I__2437 (
            .O(N__20114),
            .I(\c0.FRAME_MATCHER_state_19 ));
    SRMux I__2436 (
            .O(N__20109),
            .I(N__20106));
    LocalMux I__2435 (
            .O(N__20106),
            .I(\c0.n8_adj_2250 ));
    InMux I__2434 (
            .O(N__20103),
            .I(N__20093));
    InMux I__2433 (
            .O(N__20102),
            .I(N__20084));
    InMux I__2432 (
            .O(N__20101),
            .I(N__20081));
    InMux I__2431 (
            .O(N__20100),
            .I(N__20078));
    InMux I__2430 (
            .O(N__20099),
            .I(N__20075));
    InMux I__2429 (
            .O(N__20098),
            .I(N__20072));
    InMux I__2428 (
            .O(N__20097),
            .I(N__20069));
    InMux I__2427 (
            .O(N__20096),
            .I(N__20066));
    LocalMux I__2426 (
            .O(N__20093),
            .I(N__20062));
    InMux I__2425 (
            .O(N__20092),
            .I(N__20059));
    InMux I__2424 (
            .O(N__20091),
            .I(N__20056));
    InMux I__2423 (
            .O(N__20090),
            .I(N__20052));
    InMux I__2422 (
            .O(N__20089),
            .I(N__20049));
    InMux I__2421 (
            .O(N__20088),
            .I(N__20046));
    InMux I__2420 (
            .O(N__20087),
            .I(N__20043));
    LocalMux I__2419 (
            .O(N__20084),
            .I(N__20038));
    LocalMux I__2418 (
            .O(N__20081),
            .I(N__20035));
    LocalMux I__2417 (
            .O(N__20078),
            .I(N__20024));
    LocalMux I__2416 (
            .O(N__20075),
            .I(N__20024));
    LocalMux I__2415 (
            .O(N__20072),
            .I(N__20024));
    LocalMux I__2414 (
            .O(N__20069),
            .I(N__20024));
    LocalMux I__2413 (
            .O(N__20066),
            .I(N__20024));
    InMux I__2412 (
            .O(N__20065),
            .I(N__20021));
    Span4Mux_s2_v I__2411 (
            .O(N__20062),
            .I(N__20015));
    LocalMux I__2410 (
            .O(N__20059),
            .I(N__20015));
    LocalMux I__2409 (
            .O(N__20056),
            .I(N__20012));
    InMux I__2408 (
            .O(N__20055),
            .I(N__20009));
    LocalMux I__2407 (
            .O(N__20052),
            .I(N__20002));
    LocalMux I__2406 (
            .O(N__20049),
            .I(N__20002));
    LocalMux I__2405 (
            .O(N__20046),
            .I(N__20002));
    LocalMux I__2404 (
            .O(N__20043),
            .I(N__19999));
    InMux I__2403 (
            .O(N__20042),
            .I(N__19996));
    InMux I__2402 (
            .O(N__20041),
            .I(N__19993));
    Span4Mux_v I__2401 (
            .O(N__20038),
            .I(N__19983));
    Span4Mux_v I__2400 (
            .O(N__20035),
            .I(N__19983));
    Span4Mux_v I__2399 (
            .O(N__20024),
            .I(N__19983));
    LocalMux I__2398 (
            .O(N__20021),
            .I(N__19980));
    InMux I__2397 (
            .O(N__20020),
            .I(N__19977));
    Span4Mux_h I__2396 (
            .O(N__20015),
            .I(N__19970));
    Span4Mux_s2_v I__2395 (
            .O(N__20012),
            .I(N__19970));
    LocalMux I__2394 (
            .O(N__20009),
            .I(N__19970));
    Span4Mux_v I__2393 (
            .O(N__20002),
            .I(N__19963));
    Span4Mux_v I__2392 (
            .O(N__19999),
            .I(N__19963));
    LocalMux I__2391 (
            .O(N__19996),
            .I(N__19963));
    LocalMux I__2390 (
            .O(N__19993),
            .I(N__19960));
    InMux I__2389 (
            .O(N__19992),
            .I(N__19957));
    InMux I__2388 (
            .O(N__19991),
            .I(N__19954));
    InMux I__2387 (
            .O(N__19990),
            .I(N__19951));
    Odrv4 I__2386 (
            .O(N__19983),
            .I(\c0.n4_adj_2271 ));
    Odrv4 I__2385 (
            .O(N__19980),
            .I(\c0.n4_adj_2271 ));
    LocalMux I__2384 (
            .O(N__19977),
            .I(\c0.n4_adj_2271 ));
    Odrv4 I__2383 (
            .O(N__19970),
            .I(\c0.n4_adj_2271 ));
    Odrv4 I__2382 (
            .O(N__19963),
            .I(\c0.n4_adj_2271 ));
    Odrv4 I__2381 (
            .O(N__19960),
            .I(\c0.n4_adj_2271 ));
    LocalMux I__2380 (
            .O(N__19957),
            .I(\c0.n4_adj_2271 ));
    LocalMux I__2379 (
            .O(N__19954),
            .I(\c0.n4_adj_2271 ));
    LocalMux I__2378 (
            .O(N__19951),
            .I(\c0.n4_adj_2271 ));
    InMux I__2377 (
            .O(N__19932),
            .I(N__19929));
    LocalMux I__2376 (
            .O(N__19929),
            .I(N__19926));
    Span4Mux_v I__2375 (
            .O(N__19926),
            .I(N__19923));
    Odrv4 I__2374 (
            .O(N__19923),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_22 ));
    InMux I__2373 (
            .O(N__19920),
            .I(N__19916));
    InMux I__2372 (
            .O(N__19919),
            .I(N__19912));
    LocalMux I__2371 (
            .O(N__19916),
            .I(N__19909));
    InMux I__2370 (
            .O(N__19915),
            .I(N__19906));
    LocalMux I__2369 (
            .O(N__19912),
            .I(N__19902));
    Span4Mux_v I__2368 (
            .O(N__19909),
            .I(N__19897));
    LocalMux I__2367 (
            .O(N__19906),
            .I(N__19897));
    InMux I__2366 (
            .O(N__19905),
            .I(N__19894));
    Span4Mux_h I__2365 (
            .O(N__19902),
            .I(N__19891));
    Span4Mux_v I__2364 (
            .O(N__19897),
            .I(N__19888));
    LocalMux I__2363 (
            .O(N__19894),
            .I(N__19885));
    Odrv4 I__2362 (
            .O(N__19891),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__2361 (
            .O(N__19888),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__2360 (
            .O(N__19885),
            .I(\c0.FRAME_MATCHER_i_22 ));
    InMux I__2359 (
            .O(N__19878),
            .I(N__19875));
    LocalMux I__2358 (
            .O(N__19875),
            .I(N__19872));
    Span4Mux_s3_h I__2357 (
            .O(N__19872),
            .I(N__19869));
    Odrv4 I__2356 (
            .O(N__19869),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_22 ));
    InMux I__2355 (
            .O(N__19866),
            .I(\c0.n16507 ));
    InMux I__2354 (
            .O(N__19863),
            .I(N__19860));
    LocalMux I__2353 (
            .O(N__19860),
            .I(N__19857));
    Odrv4 I__2352 (
            .O(N__19857),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_23 ));
    InMux I__2351 (
            .O(N__19854),
            .I(N__19848));
    InMux I__2350 (
            .O(N__19853),
            .I(N__19845));
    InMux I__2349 (
            .O(N__19852),
            .I(N__19842));
    InMux I__2348 (
            .O(N__19851),
            .I(N__19839));
    LocalMux I__2347 (
            .O(N__19848),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__2346 (
            .O(N__19845),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__2345 (
            .O(N__19842),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__2344 (
            .O(N__19839),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__2343 (
            .O(N__19830),
            .I(N__19827));
    LocalMux I__2342 (
            .O(N__19827),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_23 ));
    InMux I__2341 (
            .O(N__19824),
            .I(\c0.n16508 ));
    InMux I__2340 (
            .O(N__19821),
            .I(N__19818));
    LocalMux I__2339 (
            .O(N__19818),
            .I(N__19815));
    Span4Mux_v I__2338 (
            .O(N__19815),
            .I(N__19812));
    Odrv4 I__2337 (
            .O(N__19812),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_24 ));
    InMux I__2336 (
            .O(N__19809),
            .I(N__19806));
    LocalMux I__2335 (
            .O(N__19806),
            .I(N__19801));
    CascadeMux I__2334 (
            .O(N__19805),
            .I(N__19798));
    InMux I__2333 (
            .O(N__19804),
            .I(N__19794));
    Span4Mux_h I__2332 (
            .O(N__19801),
            .I(N__19791));
    InMux I__2331 (
            .O(N__19798),
            .I(N__19786));
    InMux I__2330 (
            .O(N__19797),
            .I(N__19786));
    LocalMux I__2329 (
            .O(N__19794),
            .I(N__19783));
    Span4Mux_v I__2328 (
            .O(N__19791),
            .I(N__19780));
    LocalMux I__2327 (
            .O(N__19786),
            .I(N__19777));
    Odrv4 I__2326 (
            .O(N__19783),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__2325 (
            .O(N__19780),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__2324 (
            .O(N__19777),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__2323 (
            .O(N__19770),
            .I(N__19767));
    LocalMux I__2322 (
            .O(N__19767),
            .I(N__19764));
    Odrv12 I__2321 (
            .O(N__19764),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_24 ));
    InMux I__2320 (
            .O(N__19761),
            .I(bfn_4_14_0_));
    InMux I__2319 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__2318 (
            .O(N__19755),
            .I(N__19752));
    Odrv12 I__2317 (
            .O(N__19752),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_25 ));
    InMux I__2316 (
            .O(N__19749),
            .I(N__19743));
    CascadeMux I__2315 (
            .O(N__19748),
            .I(N__19740));
    InMux I__2314 (
            .O(N__19747),
            .I(N__19737));
    InMux I__2313 (
            .O(N__19746),
            .I(N__19734));
    LocalMux I__2312 (
            .O(N__19743),
            .I(N__19731));
    InMux I__2311 (
            .O(N__19740),
            .I(N__19728));
    LocalMux I__2310 (
            .O(N__19737),
            .I(N__19725));
    LocalMux I__2309 (
            .O(N__19734),
            .I(N__19722));
    Span4Mux_h I__2308 (
            .O(N__19731),
            .I(N__19719));
    LocalMux I__2307 (
            .O(N__19728),
            .I(N__19716));
    Span4Mux_h I__2306 (
            .O(N__19725),
            .I(N__19713));
    Span4Mux_h I__2305 (
            .O(N__19722),
            .I(N__19710));
    Odrv4 I__2304 (
            .O(N__19719),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv12 I__2303 (
            .O(N__19716),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__2302 (
            .O(N__19713),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__2301 (
            .O(N__19710),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__2300 (
            .O(N__19701),
            .I(N__19698));
    LocalMux I__2299 (
            .O(N__19698),
            .I(N__19695));
    Odrv4 I__2298 (
            .O(N__19695),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_25 ));
    InMux I__2297 (
            .O(N__19692),
            .I(\c0.n16510 ));
    InMux I__2296 (
            .O(N__19689),
            .I(N__19686));
    LocalMux I__2295 (
            .O(N__19686),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_26 ));
    InMux I__2294 (
            .O(N__19683),
            .I(\c0.n16511 ));
    InMux I__2293 (
            .O(N__19680),
            .I(\c0.n16512 ));
    InMux I__2292 (
            .O(N__19677),
            .I(\c0.n16513 ));
    InMux I__2291 (
            .O(N__19674),
            .I(N__19671));
    LocalMux I__2290 (
            .O(N__19671),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_29 ));
    InMux I__2289 (
            .O(N__19668),
            .I(\c0.n16514 ));
    InMux I__2288 (
            .O(N__19665),
            .I(N__19662));
    LocalMux I__2287 (
            .O(N__19662),
            .I(N__19659));
    Span4Mux_v I__2286 (
            .O(N__19659),
            .I(N__19656));
    Odrv4 I__2285 (
            .O(N__19656),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_14 ));
    InMux I__2284 (
            .O(N__19653),
            .I(\c0.n16499 ));
    InMux I__2283 (
            .O(N__19650),
            .I(N__19647));
    LocalMux I__2282 (
            .O(N__19647),
            .I(N__19644));
    Span4Mux_v I__2281 (
            .O(N__19644),
            .I(N__19641));
    Odrv4 I__2280 (
            .O(N__19641),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_15 ));
    InMux I__2279 (
            .O(N__19638),
            .I(N__19634));
    CascadeMux I__2278 (
            .O(N__19637),
            .I(N__19631));
    LocalMux I__2277 (
            .O(N__19634),
            .I(N__19627));
    InMux I__2276 (
            .O(N__19631),
            .I(N__19624));
    InMux I__2275 (
            .O(N__19630),
            .I(N__19620));
    Span4Mux_h I__2274 (
            .O(N__19627),
            .I(N__19617));
    LocalMux I__2273 (
            .O(N__19624),
            .I(N__19614));
    InMux I__2272 (
            .O(N__19623),
            .I(N__19611));
    LocalMux I__2271 (
            .O(N__19620),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__2270 (
            .O(N__19617),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__2269 (
            .O(N__19614),
            .I(\c0.FRAME_MATCHER_i_15 ));
    LocalMux I__2268 (
            .O(N__19611),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__2267 (
            .O(N__19602),
            .I(N__19599));
    LocalMux I__2266 (
            .O(N__19599),
            .I(N__19596));
    Odrv4 I__2265 (
            .O(N__19596),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_15 ));
    InMux I__2264 (
            .O(N__19593),
            .I(\c0.n16500 ));
    InMux I__2263 (
            .O(N__19590),
            .I(N__19587));
    LocalMux I__2262 (
            .O(N__19587),
            .I(N__19584));
    Odrv4 I__2261 (
            .O(N__19584),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_16 ));
    CascadeMux I__2260 (
            .O(N__19581),
            .I(N__19578));
    InMux I__2259 (
            .O(N__19578),
            .I(N__19574));
    CascadeMux I__2258 (
            .O(N__19577),
            .I(N__19570));
    LocalMux I__2257 (
            .O(N__19574),
            .I(N__19567));
    InMux I__2256 (
            .O(N__19573),
            .I(N__19561));
    InMux I__2255 (
            .O(N__19570),
            .I(N__19561));
    Span4Mux_v I__2254 (
            .O(N__19567),
            .I(N__19558));
    InMux I__2253 (
            .O(N__19566),
            .I(N__19555));
    LocalMux I__2252 (
            .O(N__19561),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__2251 (
            .O(N__19558),
            .I(\c0.FRAME_MATCHER_i_16 ));
    LocalMux I__2250 (
            .O(N__19555),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__2249 (
            .O(N__19548),
            .I(N__19545));
    LocalMux I__2248 (
            .O(N__19545),
            .I(N__19542));
    Odrv4 I__2247 (
            .O(N__19542),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_16 ));
    InMux I__2246 (
            .O(N__19539),
            .I(bfn_4_13_0_));
    InMux I__2245 (
            .O(N__19536),
            .I(N__19533));
    LocalMux I__2244 (
            .O(N__19533),
            .I(N__19530));
    Span4Mux_v I__2243 (
            .O(N__19530),
            .I(N__19527));
    Odrv4 I__2242 (
            .O(N__19527),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_17 ));
    CascadeMux I__2241 (
            .O(N__19524),
            .I(N__19521));
    InMux I__2240 (
            .O(N__19521),
            .I(N__19517));
    CascadeMux I__2239 (
            .O(N__19520),
            .I(N__19514));
    LocalMux I__2238 (
            .O(N__19517),
            .I(N__19509));
    InMux I__2237 (
            .O(N__19514),
            .I(N__19506));
    InMux I__2236 (
            .O(N__19513),
            .I(N__19503));
    InMux I__2235 (
            .O(N__19512),
            .I(N__19500));
    Span4Mux_h I__2234 (
            .O(N__19509),
            .I(N__19497));
    LocalMux I__2233 (
            .O(N__19506),
            .I(N__19494));
    LocalMux I__2232 (
            .O(N__19503),
            .I(N__19491));
    LocalMux I__2231 (
            .O(N__19500),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__2230 (
            .O(N__19497),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__2229 (
            .O(N__19494),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__2228 (
            .O(N__19491),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__2227 (
            .O(N__19482),
            .I(N__19479));
    LocalMux I__2226 (
            .O(N__19479),
            .I(N__19476));
    Odrv12 I__2225 (
            .O(N__19476),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_17 ));
    InMux I__2224 (
            .O(N__19473),
            .I(\c0.n16502 ));
    InMux I__2223 (
            .O(N__19470),
            .I(\c0.n16503 ));
    InMux I__2222 (
            .O(N__19467),
            .I(N__19464));
    LocalMux I__2221 (
            .O(N__19464),
            .I(N__19461));
    Span4Mux_v I__2220 (
            .O(N__19461),
            .I(N__19458));
    Odrv4 I__2219 (
            .O(N__19458),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_19 ));
    InMux I__2218 (
            .O(N__19455),
            .I(\c0.n16504 ));
    InMux I__2217 (
            .O(N__19452),
            .I(N__19449));
    LocalMux I__2216 (
            .O(N__19449),
            .I(N__19446));
    Span4Mux_v I__2215 (
            .O(N__19446),
            .I(N__19443));
    Odrv4 I__2214 (
            .O(N__19443),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_20 ));
    InMux I__2213 (
            .O(N__19440),
            .I(\c0.n16505 ));
    InMux I__2212 (
            .O(N__19437),
            .I(N__19434));
    LocalMux I__2211 (
            .O(N__19434),
            .I(N__19431));
    Span4Mux_v I__2210 (
            .O(N__19431),
            .I(N__19428));
    Odrv4 I__2209 (
            .O(N__19428),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_21 ));
    InMux I__2208 (
            .O(N__19425),
            .I(N__19422));
    LocalMux I__2207 (
            .O(N__19422),
            .I(N__19418));
    CascadeMux I__2206 (
            .O(N__19421),
            .I(N__19415));
    Span4Mux_v I__2205 (
            .O(N__19418),
            .I(N__19412));
    InMux I__2204 (
            .O(N__19415),
            .I(N__19409));
    Span4Mux_v I__2203 (
            .O(N__19412),
            .I(N__19402));
    LocalMux I__2202 (
            .O(N__19409),
            .I(N__19402));
    InMux I__2201 (
            .O(N__19408),
            .I(N__19397));
    InMux I__2200 (
            .O(N__19407),
            .I(N__19397));
    Odrv4 I__2199 (
            .O(N__19402),
            .I(\c0.FRAME_MATCHER_i_21 ));
    LocalMux I__2198 (
            .O(N__19397),
            .I(\c0.FRAME_MATCHER_i_21 ));
    InMux I__2197 (
            .O(N__19392),
            .I(N__19389));
    LocalMux I__2196 (
            .O(N__19389),
            .I(N__19386));
    Odrv4 I__2195 (
            .O(N__19386),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_21 ));
    InMux I__2194 (
            .O(N__19383),
            .I(\c0.n16506 ));
    InMux I__2193 (
            .O(N__19380),
            .I(\c0.n16491 ));
    InMux I__2192 (
            .O(N__19377),
            .I(N__19374));
    LocalMux I__2191 (
            .O(N__19374),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_7 ));
    InMux I__2190 (
            .O(N__19371),
            .I(N__19368));
    LocalMux I__2189 (
            .O(N__19368),
            .I(N__19362));
    InMux I__2188 (
            .O(N__19367),
            .I(N__19359));
    InMux I__2187 (
            .O(N__19366),
            .I(N__19356));
    InMux I__2186 (
            .O(N__19365),
            .I(N__19353));
    Span4Mux_s3_h I__2185 (
            .O(N__19362),
            .I(N__19350));
    LocalMux I__2184 (
            .O(N__19359),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__2183 (
            .O(N__19356),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__2182 (
            .O(N__19353),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv4 I__2181 (
            .O(N__19350),
            .I(\c0.FRAME_MATCHER_i_7 ));
    InMux I__2180 (
            .O(N__19341),
            .I(N__19338));
    LocalMux I__2179 (
            .O(N__19338),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_7 ));
    InMux I__2178 (
            .O(N__19335),
            .I(\c0.n16492 ));
    InMux I__2177 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__2176 (
            .O(N__19329),
            .I(N__19326));
    Odrv4 I__2175 (
            .O(N__19326),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_8 ));
    InMux I__2174 (
            .O(N__19323),
            .I(N__19319));
    InMux I__2173 (
            .O(N__19322),
            .I(N__19314));
    LocalMux I__2172 (
            .O(N__19319),
            .I(N__19311));
    InMux I__2171 (
            .O(N__19318),
            .I(N__19308));
    InMux I__2170 (
            .O(N__19317),
            .I(N__19305));
    LocalMux I__2169 (
            .O(N__19314),
            .I(N__19302));
    Span4Mux_v I__2168 (
            .O(N__19311),
            .I(N__19297));
    LocalMux I__2167 (
            .O(N__19308),
            .I(N__19297));
    LocalMux I__2166 (
            .O(N__19305),
            .I(N__19294));
    Span4Mux_v I__2165 (
            .O(N__19302),
            .I(N__19291));
    Span4Mux_v I__2164 (
            .O(N__19297),
            .I(N__19288));
    Span4Mux_s2_h I__2163 (
            .O(N__19294),
            .I(N__19285));
    Odrv4 I__2162 (
            .O(N__19291),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv4 I__2161 (
            .O(N__19288),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv4 I__2160 (
            .O(N__19285),
            .I(\c0.FRAME_MATCHER_i_8 ));
    InMux I__2159 (
            .O(N__19278),
            .I(N__19275));
    LocalMux I__2158 (
            .O(N__19275),
            .I(N__19272));
    Span4Mux_v I__2157 (
            .O(N__19272),
            .I(N__19269));
    Odrv4 I__2156 (
            .O(N__19269),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_8 ));
    InMux I__2155 (
            .O(N__19266),
            .I(bfn_4_12_0_));
    InMux I__2154 (
            .O(N__19263),
            .I(N__19260));
    LocalMux I__2153 (
            .O(N__19260),
            .I(N__19257));
    Odrv4 I__2152 (
            .O(N__19257),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_9 ));
    InMux I__2151 (
            .O(N__19254),
            .I(\c0.n16494 ));
    InMux I__2150 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__2149 (
            .O(N__19248),
            .I(N__19245));
    Span4Mux_s3_h I__2148 (
            .O(N__19245),
            .I(N__19242));
    Odrv4 I__2147 (
            .O(N__19242),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_10 ));
    InMux I__2146 (
            .O(N__19239),
            .I(\c0.n16495 ));
    InMux I__2145 (
            .O(N__19236),
            .I(\c0.n16496 ));
    InMux I__2144 (
            .O(N__19233),
            .I(N__19230));
    LocalMux I__2143 (
            .O(N__19230),
            .I(N__19227));
    Span4Mux_s3_h I__2142 (
            .O(N__19227),
            .I(N__19224));
    Odrv4 I__2141 (
            .O(N__19224),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_12 ));
    InMux I__2140 (
            .O(N__19221),
            .I(\c0.n16497 ));
    InMux I__2139 (
            .O(N__19218),
            .I(\c0.n16498 ));
    InMux I__2138 (
            .O(N__19215),
            .I(N__19212));
    LocalMux I__2137 (
            .O(N__19212),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_0 ));
    InMux I__2136 (
            .O(N__19209),
            .I(bfn_4_11_0_));
    InMux I__2135 (
            .O(N__19206),
            .I(N__19203));
    LocalMux I__2134 (
            .O(N__19203),
            .I(N__19200));
    Span4Mux_s3_h I__2133 (
            .O(N__19200),
            .I(N__19197));
    Odrv4 I__2132 (
            .O(N__19197),
            .I(\c0.n27_adj_2426 ));
    InMux I__2131 (
            .O(N__19194),
            .I(\c0.n16486 ));
    InMux I__2130 (
            .O(N__19191),
            .I(N__19188));
    LocalMux I__2129 (
            .O(N__19188),
            .I(N__19185));
    Span4Mux_v I__2128 (
            .O(N__19185),
            .I(N__19182));
    Odrv4 I__2127 (
            .O(N__19182),
            .I(\c0.n115 ));
    InMux I__2126 (
            .O(N__19179),
            .I(N__19176));
    LocalMux I__2125 (
            .O(N__19176),
            .I(N__19173));
    Span4Mux_s3_h I__2124 (
            .O(N__19173),
            .I(N__19170));
    Odrv4 I__2123 (
            .O(N__19170),
            .I(\c0.n29 ));
    InMux I__2122 (
            .O(N__19167),
            .I(\c0.n16487 ));
    InMux I__2121 (
            .O(N__19164),
            .I(\c0.n16488 ));
    InMux I__2120 (
            .O(N__19161),
            .I(N__19158));
    LocalMux I__2119 (
            .O(N__19158),
            .I(N__19155));
    Odrv4 I__2118 (
            .O(N__19155),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_4 ));
    InMux I__2117 (
            .O(N__19152),
            .I(\c0.n16489 ));
    InMux I__2116 (
            .O(N__19149),
            .I(\c0.n16490 ));
    InMux I__2115 (
            .O(N__19146),
            .I(N__19120));
    InMux I__2114 (
            .O(N__19145),
            .I(N__19120));
    InMux I__2113 (
            .O(N__19144),
            .I(N__19120));
    InMux I__2112 (
            .O(N__19143),
            .I(N__19120));
    InMux I__2111 (
            .O(N__19142),
            .I(N__19104));
    InMux I__2110 (
            .O(N__19141),
            .I(N__19104));
    InMux I__2109 (
            .O(N__19140),
            .I(N__19104));
    InMux I__2108 (
            .O(N__19139),
            .I(N__19104));
    InMux I__2107 (
            .O(N__19138),
            .I(N__19104));
    InMux I__2106 (
            .O(N__19137),
            .I(N__19104));
    InMux I__2105 (
            .O(N__19136),
            .I(N__19104));
    InMux I__2104 (
            .O(N__19135),
            .I(N__19089));
    InMux I__2103 (
            .O(N__19134),
            .I(N__19089));
    InMux I__2102 (
            .O(N__19133),
            .I(N__19089));
    InMux I__2101 (
            .O(N__19132),
            .I(N__19089));
    InMux I__2100 (
            .O(N__19131),
            .I(N__19089));
    InMux I__2099 (
            .O(N__19130),
            .I(N__19089));
    InMux I__2098 (
            .O(N__19129),
            .I(N__19089));
    LocalMux I__2097 (
            .O(N__19120),
            .I(N__19083));
    InMux I__2096 (
            .O(N__19119),
            .I(N__19080));
    LocalMux I__2095 (
            .O(N__19104),
            .I(N__19075));
    LocalMux I__2094 (
            .O(N__19089),
            .I(N__19075));
    InMux I__2093 (
            .O(N__19088),
            .I(N__19072));
    InMux I__2092 (
            .O(N__19087),
            .I(N__19067));
    InMux I__2091 (
            .O(N__19086),
            .I(N__19067));
    Span4Mux_s3_h I__2090 (
            .O(N__19083),
            .I(N__19063));
    LocalMux I__2089 (
            .O(N__19080),
            .I(N__19060));
    Span4Mux_s3_h I__2088 (
            .O(N__19075),
            .I(N__19053));
    LocalMux I__2087 (
            .O(N__19072),
            .I(N__19053));
    LocalMux I__2086 (
            .O(N__19067),
            .I(N__19053));
    InMux I__2085 (
            .O(N__19066),
            .I(N__19050));
    Odrv4 I__2084 (
            .O(N__19063),
            .I(\c0.n9575 ));
    Odrv12 I__2083 (
            .O(N__19060),
            .I(\c0.n9575 ));
    Odrv4 I__2082 (
            .O(N__19053),
            .I(\c0.n9575 ));
    LocalMux I__2081 (
            .O(N__19050),
            .I(\c0.n9575 ));
    InMux I__2080 (
            .O(N__19041),
            .I(N__19036));
    InMux I__2079 (
            .O(N__19040),
            .I(N__19033));
    InMux I__2078 (
            .O(N__19039),
            .I(N__19030));
    LocalMux I__2077 (
            .O(N__19036),
            .I(n12966));
    LocalMux I__2076 (
            .O(N__19033),
            .I(n12966));
    LocalMux I__2075 (
            .O(N__19030),
            .I(n12966));
    InMux I__2074 (
            .O(N__19023),
            .I(N__19020));
    LocalMux I__2073 (
            .O(N__19020),
            .I(N__19017));
    Span4Mux_v I__2072 (
            .O(N__19017),
            .I(N__19013));
    InMux I__2071 (
            .O(N__19016),
            .I(N__19010));
    Odrv4 I__2070 (
            .O(N__19013),
            .I(n15118));
    LocalMux I__2069 (
            .O(N__19010),
            .I(n15118));
    InMux I__2068 (
            .O(N__19005),
            .I(N__18997));
    InMux I__2067 (
            .O(N__19004),
            .I(N__18994));
    InMux I__2066 (
            .O(N__19003),
            .I(N__18991));
    InMux I__2065 (
            .O(N__19002),
            .I(N__18986));
    InMux I__2064 (
            .O(N__19001),
            .I(N__18986));
    InMux I__2063 (
            .O(N__19000),
            .I(N__18983));
    LocalMux I__2062 (
            .O(N__18997),
            .I(N__18980));
    LocalMux I__2061 (
            .O(N__18994),
            .I(N__18977));
    LocalMux I__2060 (
            .O(N__18991),
            .I(N__18974));
    LocalMux I__2059 (
            .O(N__18986),
            .I(N__18969));
    LocalMux I__2058 (
            .O(N__18983),
            .I(N__18969));
    Span4Mux_v I__2057 (
            .O(N__18980),
            .I(N__18966));
    Span4Mux_v I__2056 (
            .O(N__18977),
            .I(N__18963));
    Span4Mux_s2_h I__2055 (
            .O(N__18974),
            .I(N__18958));
    Span4Mux_v I__2054 (
            .O(N__18969),
            .I(N__18958));
    Odrv4 I__2053 (
            .O(N__18966),
            .I(FRAME_MATCHER_i_31__N_1273));
    Odrv4 I__2052 (
            .O(N__18963),
            .I(FRAME_MATCHER_i_31__N_1273));
    Odrv4 I__2051 (
            .O(N__18958),
            .I(FRAME_MATCHER_i_31__N_1273));
    CascadeMux I__2050 (
            .O(N__18951),
            .I(\c0.n16685_cascade_ ));
    InMux I__2049 (
            .O(N__18948),
            .I(N__18945));
    LocalMux I__2048 (
            .O(N__18945),
            .I(\c0.n6_adj_2267 ));
    InMux I__2047 (
            .O(N__18942),
            .I(N__18937));
    InMux I__2046 (
            .O(N__18941),
            .I(N__18932));
    InMux I__2045 (
            .O(N__18940),
            .I(N__18932));
    LocalMux I__2044 (
            .O(N__18937),
            .I(N__18929));
    LocalMux I__2043 (
            .O(N__18932),
            .I(N__18926));
    Span4Mux_v I__2042 (
            .O(N__18929),
            .I(N__18921));
    Span4Mux_v I__2041 (
            .O(N__18926),
            .I(N__18918));
    InMux I__2040 (
            .O(N__18925),
            .I(N__18913));
    InMux I__2039 (
            .O(N__18924),
            .I(N__18913));
    Odrv4 I__2038 (
            .O(N__18921),
            .I(FRAME_MATCHER_i_31__N_1270));
    Odrv4 I__2037 (
            .O(N__18918),
            .I(FRAME_MATCHER_i_31__N_1270));
    LocalMux I__2036 (
            .O(N__18913),
            .I(FRAME_MATCHER_i_31__N_1270));
    CascadeMux I__2035 (
            .O(N__18906),
            .I(N__18902));
    CascadeMux I__2034 (
            .O(N__18905),
            .I(N__18899));
    InMux I__2033 (
            .O(N__18902),
            .I(N__18894));
    InMux I__2032 (
            .O(N__18899),
            .I(N__18894));
    LocalMux I__2031 (
            .O(N__18894),
            .I(N__18891));
    Odrv4 I__2030 (
            .O(N__18891),
            .I(\c0.n7528 ));
    InMux I__2029 (
            .O(N__18888),
            .I(N__18884));
    InMux I__2028 (
            .O(N__18887),
            .I(N__18881));
    LocalMux I__2027 (
            .O(N__18884),
            .I(N__18878));
    LocalMux I__2026 (
            .O(N__18881),
            .I(N__18875));
    Span4Mux_s3_h I__2025 (
            .O(N__18878),
            .I(N__18872));
    Span12Mux_s3_v I__2024 (
            .O(N__18875),
            .I(N__18869));
    Odrv4 I__2023 (
            .O(N__18872),
            .I(\c0.n46 ));
    Odrv12 I__2022 (
            .O(N__18869),
            .I(\c0.n46 ));
    SRMux I__2021 (
            .O(N__18864),
            .I(N__18861));
    LocalMux I__2020 (
            .O(N__18861),
            .I(N__18858));
    Span4Mux_h I__2019 (
            .O(N__18858),
            .I(N__18855));
    Odrv4 I__2018 (
            .O(N__18855),
            .I(\c0.n3_adj_2332 ));
    SRMux I__2017 (
            .O(N__18852),
            .I(N__18849));
    LocalMux I__2016 (
            .O(N__18849),
            .I(N__18846));
    Span4Mux_s3_h I__2015 (
            .O(N__18846),
            .I(N__18843));
    Span4Mux_v I__2014 (
            .O(N__18843),
            .I(N__18840));
    Odrv4 I__2013 (
            .O(N__18840),
            .I(\c0.n3_adj_2330 ));
    CascadeMux I__2012 (
            .O(N__18837),
            .I(\c0.n9575_cascade_ ));
    InMux I__2011 (
            .O(N__18834),
            .I(N__18830));
    InMux I__2010 (
            .O(N__18833),
            .I(N__18827));
    LocalMux I__2009 (
            .O(N__18830),
            .I(n12999));
    LocalMux I__2008 (
            .O(N__18827),
            .I(n12999));
    InMux I__2007 (
            .O(N__18822),
            .I(N__18819));
    LocalMux I__2006 (
            .O(N__18819),
            .I(N__18815));
    CascadeMux I__2005 (
            .O(N__18818),
            .I(N__18812));
    Span4Mux_v I__2004 (
            .O(N__18815),
            .I(N__18809));
    InMux I__2003 (
            .O(N__18812),
            .I(N__18806));
    Odrv4 I__2002 (
            .O(N__18809),
            .I(\c0.n232 ));
    LocalMux I__2001 (
            .O(N__18806),
            .I(\c0.n232 ));
    CascadeMux I__2000 (
            .O(N__18801),
            .I(n12999_cascade_));
    InMux I__1999 (
            .O(N__18798),
            .I(N__18795));
    LocalMux I__1998 (
            .O(N__18795),
            .I(N__18792));
    Odrv4 I__1997 (
            .O(N__18792),
            .I(n18));
    InMux I__1996 (
            .O(N__18789),
            .I(N__18786));
    LocalMux I__1995 (
            .O(N__18786),
            .I(N__18783));
    Span4Mux_v I__1994 (
            .O(N__18783),
            .I(N__18780));
    Odrv4 I__1993 (
            .O(N__18780),
            .I(\c0.n10346 ));
    CascadeMux I__1992 (
            .O(N__18777),
            .I(\c0.n17_cascade_ ));
    InMux I__1991 (
            .O(N__18774),
            .I(N__18771));
    LocalMux I__1990 (
            .O(N__18771),
            .I(\c0.n25_adj_2352 ));
    CascadeMux I__1989 (
            .O(N__18768),
            .I(\c0.n17962_cascade_ ));
    SRMux I__1988 (
            .O(N__18765),
            .I(N__18762));
    LocalMux I__1987 (
            .O(N__18762),
            .I(N__18759));
    Span4Mux_h I__1986 (
            .O(N__18759),
            .I(N__18756));
    Odrv4 I__1985 (
            .O(N__18756),
            .I(\c0.n4_adj_2226 ));
    CascadeMux I__1984 (
            .O(N__18753),
            .I(\c0.n2126_cascade_ ));
    InMux I__1983 (
            .O(N__18750),
            .I(N__18747));
    LocalMux I__1982 (
            .O(N__18747),
            .I(\c0.n27 ));
    CascadeMux I__1981 (
            .O(N__18744),
            .I(\c0.n23_cascade_ ));
    CascadeMux I__1980 (
            .O(N__18741),
            .I(\c0.n30_cascade_ ));
    CascadeMux I__1979 (
            .O(N__18738),
            .I(\c0.n50_cascade_ ));
    InMux I__1978 (
            .O(N__18735),
            .I(N__18732));
    LocalMux I__1977 (
            .O(N__18732),
            .I(N__18727));
    InMux I__1976 (
            .O(N__18731),
            .I(N__18722));
    InMux I__1975 (
            .O(N__18730),
            .I(N__18722));
    Span4Mux_s3_h I__1974 (
            .O(N__18727),
            .I(N__18717));
    LocalMux I__1973 (
            .O(N__18722),
            .I(N__18717));
    Odrv4 I__1972 (
            .O(N__18717),
            .I(n13849));
    InMux I__1971 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__1970 (
            .O(N__18711),
            .I(\c0.n19_adj_2351 ));
    CascadeMux I__1969 (
            .O(N__18708),
            .I(\c0.n8_adj_2273_cascade_ ));
    InMux I__1968 (
            .O(N__18705),
            .I(N__18698));
    InMux I__1967 (
            .O(N__18704),
            .I(N__18689));
    InMux I__1966 (
            .O(N__18703),
            .I(N__18689));
    InMux I__1965 (
            .O(N__18702),
            .I(N__18689));
    InMux I__1964 (
            .O(N__18701),
            .I(N__18689));
    LocalMux I__1963 (
            .O(N__18698),
            .I(\c0.n8_adj_2273 ));
    LocalMux I__1962 (
            .O(N__18689),
            .I(\c0.n8_adj_2273 ));
    InMux I__1961 (
            .O(N__18684),
            .I(N__18680));
    InMux I__1960 (
            .O(N__18683),
            .I(N__18676));
    LocalMux I__1959 (
            .O(N__18680),
            .I(N__18673));
    InMux I__1958 (
            .O(N__18679),
            .I(N__18670));
    LocalMux I__1957 (
            .O(N__18676),
            .I(\c0.FRAME_MATCHER_state_22 ));
    Odrv4 I__1956 (
            .O(N__18673),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__1955 (
            .O(N__18670),
            .I(\c0.FRAME_MATCHER_state_22 ));
    SRMux I__1954 (
            .O(N__18663),
            .I(N__18660));
    LocalMux I__1953 (
            .O(N__18660),
            .I(N__18657));
    Odrv12 I__1952 (
            .O(N__18657),
            .I(\c0.n17273 ));
    InMux I__1951 (
            .O(N__18654),
            .I(N__18649));
    InMux I__1950 (
            .O(N__18653),
            .I(N__18646));
    InMux I__1949 (
            .O(N__18652),
            .I(N__18643));
    LocalMux I__1948 (
            .O(N__18649),
            .I(\c0.FRAME_MATCHER_state_28 ));
    LocalMux I__1947 (
            .O(N__18646),
            .I(\c0.FRAME_MATCHER_state_28 ));
    LocalMux I__1946 (
            .O(N__18643),
            .I(\c0.FRAME_MATCHER_state_28 ));
    SRMux I__1945 (
            .O(N__18636),
            .I(N__18633));
    LocalMux I__1944 (
            .O(N__18633),
            .I(\c0.n17299 ));
    InMux I__1943 (
            .O(N__18630),
            .I(N__18627));
    LocalMux I__1942 (
            .O(N__18627),
            .I(N__18624));
    Odrv12 I__1941 (
            .O(N__18624),
            .I(\c0.n45 ));
    CascadeMux I__1940 (
            .O(N__18621),
            .I(N__18618));
    InMux I__1939 (
            .O(N__18618),
            .I(N__18615));
    LocalMux I__1938 (
            .O(N__18615),
            .I(N__18612));
    Odrv4 I__1937 (
            .O(N__18612),
            .I(\c0.n46_adj_2356 ));
    InMux I__1936 (
            .O(N__18609),
            .I(N__18606));
    LocalMux I__1935 (
            .O(N__18606),
            .I(\c0.n56 ));
    CascadeMux I__1934 (
            .O(N__18603),
            .I(\c0.n10513_cascade_ ));
    InMux I__1933 (
            .O(N__18600),
            .I(N__18591));
    InMux I__1932 (
            .O(N__18599),
            .I(N__18591));
    InMux I__1931 (
            .O(N__18598),
            .I(N__18587));
    InMux I__1930 (
            .O(N__18597),
            .I(N__18582));
    InMux I__1929 (
            .O(N__18596),
            .I(N__18582));
    LocalMux I__1928 (
            .O(N__18591),
            .I(N__18579));
    InMux I__1927 (
            .O(N__18590),
            .I(N__18576));
    LocalMux I__1926 (
            .O(N__18587),
            .I(N__18571));
    LocalMux I__1925 (
            .O(N__18582),
            .I(N__18571));
    Span4Mux_v I__1924 (
            .O(N__18579),
            .I(N__18566));
    LocalMux I__1923 (
            .O(N__18576),
            .I(N__18566));
    Odrv4 I__1922 (
            .O(N__18571),
            .I(FRAME_MATCHER_i_31__N_1275));
    Odrv4 I__1921 (
            .O(N__18566),
            .I(FRAME_MATCHER_i_31__N_1275));
    CascadeMux I__1920 (
            .O(N__18561),
            .I(\c0.n6033_cascade_ ));
    IoInMux I__1919 (
            .O(N__18558),
            .I(N__18555));
    LocalMux I__1918 (
            .O(N__18555),
            .I(N__18552));
    Span4Mux_s3_v I__1917 (
            .O(N__18552),
            .I(N__18549));
    Odrv4 I__1916 (
            .O(N__18549),
            .I(PIN_2_c_1));
    InMux I__1915 (
            .O(N__18546),
            .I(N__18541));
    InMux I__1914 (
            .O(N__18545),
            .I(N__18538));
    InMux I__1913 (
            .O(N__18544),
            .I(N__18535));
    LocalMux I__1912 (
            .O(N__18541),
            .I(N__18530));
    LocalMux I__1911 (
            .O(N__18538),
            .I(N__18530));
    LocalMux I__1910 (
            .O(N__18535),
            .I(N__18525));
    Span4Mux_v I__1909 (
            .O(N__18530),
            .I(N__18525));
    Odrv4 I__1908 (
            .O(N__18525),
            .I(\c0.FRAME_MATCHER_state_26 ));
    SRMux I__1907 (
            .O(N__18522),
            .I(N__18519));
    LocalMux I__1906 (
            .O(N__18519),
            .I(N__18516));
    Span4Mux_s1_v I__1905 (
            .O(N__18516),
            .I(N__18513));
    Odrv4 I__1904 (
            .O(N__18513),
            .I(\c0.n8_adj_2245 ));
    CascadeMux I__1903 (
            .O(N__18510),
            .I(N__18507));
    InMux I__1902 (
            .O(N__18507),
            .I(N__18503));
    InMux I__1901 (
            .O(N__18506),
            .I(N__18499));
    LocalMux I__1900 (
            .O(N__18503),
            .I(N__18496));
    InMux I__1899 (
            .O(N__18502),
            .I(N__18493));
    LocalMux I__1898 (
            .O(N__18499),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv12 I__1897 (
            .O(N__18496),
            .I(\c0.FRAME_MATCHER_state_24 ));
    LocalMux I__1896 (
            .O(N__18493),
            .I(\c0.FRAME_MATCHER_state_24 ));
    InMux I__1895 (
            .O(N__18486),
            .I(N__18477));
    InMux I__1894 (
            .O(N__18485),
            .I(N__18477));
    InMux I__1893 (
            .O(N__18484),
            .I(N__18477));
    LocalMux I__1892 (
            .O(N__18477),
            .I(\c0.FRAME_MATCHER_state_18 ));
    SRMux I__1891 (
            .O(N__18474),
            .I(N__18471));
    LocalMux I__1890 (
            .O(N__18471),
            .I(N__18468));
    Odrv4 I__1889 (
            .O(N__18468),
            .I(\c0.n17293 ));
    CascadeMux I__1888 (
            .O(N__18465),
            .I(N__18460));
    InMux I__1887 (
            .O(N__18464),
            .I(N__18457));
    InMux I__1886 (
            .O(N__18463),
            .I(N__18452));
    InMux I__1885 (
            .O(N__18460),
            .I(N__18452));
    LocalMux I__1884 (
            .O(N__18457),
            .I(\c0.FRAME_MATCHER_state_21 ));
    LocalMux I__1883 (
            .O(N__18452),
            .I(\c0.FRAME_MATCHER_state_21 ));
    SRMux I__1882 (
            .O(N__18447),
            .I(N__18444));
    LocalMux I__1881 (
            .O(N__18444),
            .I(N__18441));
    Span4Mux_s1_v I__1880 (
            .O(N__18441),
            .I(N__18438));
    Odrv4 I__1879 (
            .O(N__18438),
            .I(\c0.n8_adj_2247 ));
    InMux I__1878 (
            .O(N__18435),
            .I(N__18406));
    InMux I__1877 (
            .O(N__18434),
            .I(N__18406));
    InMux I__1876 (
            .O(N__18433),
            .I(N__18406));
    InMux I__1875 (
            .O(N__18432),
            .I(N__18406));
    InMux I__1874 (
            .O(N__18431),
            .I(N__18406));
    InMux I__1873 (
            .O(N__18430),
            .I(N__18406));
    InMux I__1872 (
            .O(N__18429),
            .I(N__18406));
    InMux I__1871 (
            .O(N__18428),
            .I(N__18391));
    InMux I__1870 (
            .O(N__18427),
            .I(N__18391));
    InMux I__1869 (
            .O(N__18426),
            .I(N__18391));
    InMux I__1868 (
            .O(N__18425),
            .I(N__18391));
    InMux I__1867 (
            .O(N__18424),
            .I(N__18391));
    InMux I__1866 (
            .O(N__18423),
            .I(N__18391));
    InMux I__1865 (
            .O(N__18422),
            .I(N__18391));
    InMux I__1864 (
            .O(N__18421),
            .I(N__18388));
    LocalMux I__1863 (
            .O(N__18406),
            .I(N__18385));
    LocalMux I__1862 (
            .O(N__18391),
            .I(N__18374));
    LocalMux I__1861 (
            .O(N__18388),
            .I(N__18371));
    Span4Mux_s2_h I__1860 (
            .O(N__18385),
            .I(N__18368));
    InMux I__1859 (
            .O(N__18384),
            .I(N__18353));
    InMux I__1858 (
            .O(N__18383),
            .I(N__18353));
    InMux I__1857 (
            .O(N__18382),
            .I(N__18353));
    InMux I__1856 (
            .O(N__18381),
            .I(N__18353));
    InMux I__1855 (
            .O(N__18380),
            .I(N__18353));
    InMux I__1854 (
            .O(N__18379),
            .I(N__18353));
    InMux I__1853 (
            .O(N__18378),
            .I(N__18353));
    InMux I__1852 (
            .O(N__18377),
            .I(N__18350));
    Span4Mux_v I__1851 (
            .O(N__18374),
            .I(N__18345));
    Span4Mux_v I__1850 (
            .O(N__18371),
            .I(N__18345));
    Odrv4 I__1849 (
            .O(N__18368),
            .I(\c0.n10497 ));
    LocalMux I__1848 (
            .O(N__18353),
            .I(\c0.n10497 ));
    LocalMux I__1847 (
            .O(N__18350),
            .I(\c0.n10497 ));
    Odrv4 I__1846 (
            .O(N__18345),
            .I(\c0.n10497 ));
    CascadeMux I__1845 (
            .O(N__18336),
            .I(N__18333));
    InMux I__1844 (
            .O(N__18333),
            .I(N__18330));
    LocalMux I__1843 (
            .O(N__18330),
            .I(N__18327));
    Span4Mux_v I__1842 (
            .O(N__18327),
            .I(N__18324));
    Odrv4 I__1841 (
            .O(N__18324),
            .I(\c0.n2_adj_2315 ));
    SRMux I__1840 (
            .O(N__18321),
            .I(N__18318));
    LocalMux I__1839 (
            .O(N__18318),
            .I(\c0.n3_adj_2289 ));
    SRMux I__1838 (
            .O(N__18315),
            .I(N__18312));
    LocalMux I__1837 (
            .O(N__18312),
            .I(\c0.n3_adj_2283 ));
    SRMux I__1836 (
            .O(N__18309),
            .I(N__18306));
    LocalMux I__1835 (
            .O(N__18306),
            .I(N__18303));
    Span12Mux_v I__1834 (
            .O(N__18303),
            .I(N__18300));
    Odrv12 I__1833 (
            .O(N__18300),
            .I(\c0.n3_adj_2279 ));
    SRMux I__1832 (
            .O(N__18297),
            .I(N__18294));
    LocalMux I__1831 (
            .O(N__18294),
            .I(N__18291));
    Span4Mux_s3_h I__1830 (
            .O(N__18291),
            .I(N__18288));
    Odrv4 I__1829 (
            .O(N__18288),
            .I(\c0.n3_adj_2303 ));
    CascadeMux I__1828 (
            .O(N__18285),
            .I(\c0.n10353_cascade_ ));
    SRMux I__1827 (
            .O(N__18282),
            .I(N__18279));
    LocalMux I__1826 (
            .O(N__18279),
            .I(N__18276));
    Span4Mux_s2_h I__1825 (
            .O(N__18276),
            .I(N__18273));
    Odrv4 I__1824 (
            .O(N__18273),
            .I(\c0.n3_adj_2345 ));
    SRMux I__1823 (
            .O(N__18270),
            .I(N__18267));
    LocalMux I__1822 (
            .O(N__18267),
            .I(N__18264));
    Span4Mux_v I__1821 (
            .O(N__18264),
            .I(N__18261));
    Odrv4 I__1820 (
            .O(N__18261),
            .I(\c0.n3_adj_2343 ));
    SRMux I__1819 (
            .O(N__18258),
            .I(N__18255));
    LocalMux I__1818 (
            .O(N__18255),
            .I(N__18252));
    Span4Mux_h I__1817 (
            .O(N__18252),
            .I(N__18249));
    Odrv4 I__1816 (
            .O(N__18249),
            .I(\c0.n3 ));
    SRMux I__1815 (
            .O(N__18246),
            .I(N__18243));
    LocalMux I__1814 (
            .O(N__18243),
            .I(N__18240));
    Span4Mux_s3_h I__1813 (
            .O(N__18240),
            .I(N__18237));
    Odrv4 I__1812 (
            .O(N__18237),
            .I(\c0.n3_adj_2295 ));
    SRMux I__1811 (
            .O(N__18234),
            .I(N__18231));
    LocalMux I__1810 (
            .O(N__18231),
            .I(N__18228));
    Span4Mux_v I__1809 (
            .O(N__18228),
            .I(N__18225));
    Span4Mux_s2_h I__1808 (
            .O(N__18225),
            .I(N__18222));
    Odrv4 I__1807 (
            .O(N__18222),
            .I(\c0.n3_adj_2291 ));
    CascadeMux I__1806 (
            .O(N__18219),
            .I(\c0.n232_cascade_ ));
    CascadeMux I__1805 (
            .O(N__18216),
            .I(N__18213));
    InMux I__1804 (
            .O(N__18213),
            .I(N__18210));
    LocalMux I__1803 (
            .O(N__18210),
            .I(N__18207));
    Span4Mux_s2_h I__1802 (
            .O(N__18207),
            .I(N__18204));
    Odrv4 I__1801 (
            .O(N__18204),
            .I(\c0.n6_adj_2364 ));
    CascadeMux I__1800 (
            .O(N__18201),
            .I(N__18198));
    InMux I__1799 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__1798 (
            .O(N__18195),
            .I(n237));
    CascadeMux I__1797 (
            .O(N__18192),
            .I(n237_cascade_));
    InMux I__1796 (
            .O(N__18189),
            .I(N__18186));
    LocalMux I__1795 (
            .O(N__18186),
            .I(n22_adj_2465));
    SRMux I__1794 (
            .O(N__18183),
            .I(N__18180));
    LocalMux I__1793 (
            .O(N__18180),
            .I(N__18177));
    Odrv4 I__1792 (
            .O(N__18177),
            .I(\c0.n3_adj_2309 ));
    InMux I__1791 (
            .O(N__18174),
            .I(N__18168));
    InMux I__1790 (
            .O(N__18173),
            .I(N__18168));
    LocalMux I__1789 (
            .O(N__18168),
            .I(N__18165));
    Odrv4 I__1788 (
            .O(N__18165),
            .I(n1437));
    CascadeMux I__1787 (
            .O(N__18162),
            .I(N__18157));
    InMux I__1786 (
            .O(N__18161),
            .I(N__18153));
    InMux I__1785 (
            .O(N__18160),
            .I(N__18146));
    InMux I__1784 (
            .O(N__18157),
            .I(N__18146));
    InMux I__1783 (
            .O(N__18156),
            .I(N__18146));
    LocalMux I__1782 (
            .O(N__18153),
            .I(N__18143));
    LocalMux I__1781 (
            .O(N__18146),
            .I(N__18140));
    Odrv4 I__1780 (
            .O(N__18143),
            .I(n8_adj_2498));
    Odrv12 I__1779 (
            .O(N__18140),
            .I(n8_adj_2498));
    CascadeMux I__1778 (
            .O(N__18135),
            .I(\c0.n6_adj_2265_cascade_ ));
    SRMux I__1777 (
            .O(N__18132),
            .I(N__18129));
    LocalMux I__1776 (
            .O(N__18129),
            .I(N__18126));
    Span4Mux_s3_h I__1775 (
            .O(N__18126),
            .I(N__18123));
    Odrv4 I__1774 (
            .O(N__18123),
            .I(\c0.n18907 ));
    CascadeMux I__1773 (
            .O(N__18120),
            .I(n13_adj_2469_cascade_));
    InMux I__1772 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__1771 (
            .O(N__18114),
            .I(N__18111));
    Odrv4 I__1770 (
            .O(N__18111),
            .I(n7));
    SRMux I__1769 (
            .O(N__18108),
            .I(N__18105));
    LocalMux I__1768 (
            .O(N__18105),
            .I(N__18102));
    Span4Mux_s2_h I__1767 (
            .O(N__18102),
            .I(N__18099));
    Odrv4 I__1766 (
            .O(N__18099),
            .I(\c0.n3_adj_2301 ));
    CascadeMux I__1765 (
            .O(N__18096),
            .I(n1166_cascade_));
    InMux I__1764 (
            .O(N__18093),
            .I(N__18090));
    LocalMux I__1763 (
            .O(N__18090),
            .I(N__18086));
    InMux I__1762 (
            .O(N__18089),
            .I(N__18083));
    Span4Mux_v I__1761 (
            .O(N__18086),
            .I(N__18077));
    LocalMux I__1760 (
            .O(N__18083),
            .I(N__18077));
    InMux I__1759 (
            .O(N__18082),
            .I(N__18074));
    Span4Mux_h I__1758 (
            .O(N__18077),
            .I(N__18071));
    LocalMux I__1757 (
            .O(N__18074),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__1756 (
            .O(N__18071),
            .I(\c0.FRAME_MATCHER_state_9 ));
    CascadeMux I__1755 (
            .O(N__18066),
            .I(\c0.n10497_cascade_ ));
    CascadeMux I__1754 (
            .O(N__18063),
            .I(N__18052));
    CascadeMux I__1753 (
            .O(N__18062),
            .I(N__18048));
    CascadeMux I__1752 (
            .O(N__18061),
            .I(N__18044));
    CascadeMux I__1751 (
            .O(N__18060),
            .I(N__18037));
    CascadeMux I__1750 (
            .O(N__18059),
            .I(N__18033));
    CascadeMux I__1749 (
            .O(N__18058),
            .I(N__18029));
    CascadeMux I__1748 (
            .O(N__18057),
            .I(N__18024));
    CascadeMux I__1747 (
            .O(N__18056),
            .I(N__18021));
    CascadeMux I__1746 (
            .O(N__18055),
            .I(N__18018));
    InMux I__1745 (
            .O(N__18052),
            .I(N__18000));
    InMux I__1744 (
            .O(N__18051),
            .I(N__18000));
    InMux I__1743 (
            .O(N__18048),
            .I(N__18000));
    InMux I__1742 (
            .O(N__18047),
            .I(N__18000));
    InMux I__1741 (
            .O(N__18044),
            .I(N__18000));
    InMux I__1740 (
            .O(N__18043),
            .I(N__18000));
    InMux I__1739 (
            .O(N__18042),
            .I(N__18000));
    InMux I__1738 (
            .O(N__18041),
            .I(N__17997));
    InMux I__1737 (
            .O(N__18040),
            .I(N__17994));
    InMux I__1736 (
            .O(N__18037),
            .I(N__17979));
    InMux I__1735 (
            .O(N__18036),
            .I(N__17979));
    InMux I__1734 (
            .O(N__18033),
            .I(N__17979));
    InMux I__1733 (
            .O(N__18032),
            .I(N__17979));
    InMux I__1732 (
            .O(N__18029),
            .I(N__17979));
    InMux I__1731 (
            .O(N__18028),
            .I(N__17979));
    InMux I__1730 (
            .O(N__18027),
            .I(N__17979));
    InMux I__1729 (
            .O(N__18024),
            .I(N__17966));
    InMux I__1728 (
            .O(N__18021),
            .I(N__17966));
    InMux I__1727 (
            .O(N__18018),
            .I(N__17966));
    InMux I__1726 (
            .O(N__18017),
            .I(N__17966));
    InMux I__1725 (
            .O(N__18016),
            .I(N__17966));
    InMux I__1724 (
            .O(N__18015),
            .I(N__17966));
    LocalMux I__1723 (
            .O(N__18000),
            .I(\c0.n17713 ));
    LocalMux I__1722 (
            .O(N__17997),
            .I(\c0.n17713 ));
    LocalMux I__1721 (
            .O(N__17994),
            .I(\c0.n17713 ));
    LocalMux I__1720 (
            .O(N__17979),
            .I(\c0.n17713 ));
    LocalMux I__1719 (
            .O(N__17966),
            .I(\c0.n17713 ));
    SRMux I__1718 (
            .O(N__17955),
            .I(N__17952));
    LocalMux I__1717 (
            .O(N__17952),
            .I(N__17949));
    Span4Mux_s2_h I__1716 (
            .O(N__17949),
            .I(N__17946));
    Odrv4 I__1715 (
            .O(N__17946),
            .I(\c0.n17239 ));
    CascadeMux I__1714 (
            .O(N__17943),
            .I(N__17940));
    InMux I__1713 (
            .O(N__17940),
            .I(N__17937));
    LocalMux I__1712 (
            .O(N__17937),
            .I(N__17933));
    InMux I__1711 (
            .O(N__17936),
            .I(N__17929));
    Span4Mux_v I__1710 (
            .O(N__17933),
            .I(N__17926));
    InMux I__1709 (
            .O(N__17932),
            .I(N__17923));
    LocalMux I__1708 (
            .O(N__17929),
            .I(n15));
    Odrv4 I__1707 (
            .O(N__17926),
            .I(n15));
    LocalMux I__1706 (
            .O(N__17923),
            .I(n15));
    CascadeMux I__1705 (
            .O(N__17916),
            .I(n17694_cascade_));
    CascadeMux I__1704 (
            .O(N__17913),
            .I(N__17908));
    InMux I__1703 (
            .O(N__17912),
            .I(N__17905));
    InMux I__1702 (
            .O(N__17911),
            .I(N__17900));
    InMux I__1701 (
            .O(N__17908),
            .I(N__17900));
    LocalMux I__1700 (
            .O(N__17905),
            .I(N__17897));
    LocalMux I__1699 (
            .O(N__17900),
            .I(\c0.FRAME_MATCHER_state_31 ));
    Odrv4 I__1698 (
            .O(N__17897),
            .I(\c0.FRAME_MATCHER_state_31 ));
    SRMux I__1697 (
            .O(N__17892),
            .I(N__17889));
    LocalMux I__1696 (
            .O(N__17889),
            .I(N__17886));
    Span4Mux_s3_h I__1695 (
            .O(N__17886),
            .I(N__17883));
    Odrv4 I__1694 (
            .O(N__17883),
            .I(\c0.n17279 ));
    CascadeMux I__1693 (
            .O(N__17880),
            .I(FRAME_MATCHER_state_31_N_1406_0_cascade_));
    CascadeMux I__1692 (
            .O(N__17877),
            .I(N__17873));
    InMux I__1691 (
            .O(N__17876),
            .I(N__17867));
    InMux I__1690 (
            .O(N__17873),
            .I(N__17867));
    InMux I__1689 (
            .O(N__17872),
            .I(N__17864));
    LocalMux I__1688 (
            .O(N__17867),
            .I(\c0.FRAME_MATCHER_state_17 ));
    LocalMux I__1687 (
            .O(N__17864),
            .I(\c0.FRAME_MATCHER_state_17 ));
    SRMux I__1686 (
            .O(N__17859),
            .I(N__17856));
    LocalMux I__1685 (
            .O(N__17856),
            .I(N__17853));
    Span4Mux_s3_h I__1684 (
            .O(N__17853),
            .I(N__17850));
    Odrv4 I__1683 (
            .O(N__17850),
            .I(\c0.n8_adj_2252 ));
    SRMux I__1682 (
            .O(N__17847),
            .I(N__17844));
    LocalMux I__1681 (
            .O(N__17844),
            .I(N__17841));
    Span4Mux_s1_v I__1680 (
            .O(N__17841),
            .I(N__17838));
    Odrv4 I__1679 (
            .O(N__17838),
            .I(\c0.n8_adj_2246 ));
    CascadeMux I__1678 (
            .O(N__17835),
            .I(N__17831));
    CascadeMux I__1677 (
            .O(N__17834),
            .I(N__17828));
    InMux I__1676 (
            .O(N__17831),
            .I(N__17825));
    InMux I__1675 (
            .O(N__17828),
            .I(N__17822));
    LocalMux I__1674 (
            .O(N__17825),
            .I(N__17816));
    LocalMux I__1673 (
            .O(N__17822),
            .I(N__17816));
    InMux I__1672 (
            .O(N__17821),
            .I(N__17813));
    Span4Mux_v I__1671 (
            .O(N__17816),
            .I(N__17810));
    LocalMux I__1670 (
            .O(N__17813),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv4 I__1669 (
            .O(N__17810),
            .I(\c0.FRAME_MATCHER_state_27 ));
    SRMux I__1668 (
            .O(N__17805),
            .I(N__17802));
    LocalMux I__1667 (
            .O(N__17802),
            .I(N__17799));
    Span4Mux_s2_h I__1666 (
            .O(N__17799),
            .I(N__17796));
    Odrv4 I__1665 (
            .O(N__17796),
            .I(\c0.n17277 ));
    CascadeMux I__1664 (
            .O(N__17793),
            .I(N__17789));
    InMux I__1663 (
            .O(N__17792),
            .I(N__17786));
    InMux I__1662 (
            .O(N__17789),
            .I(N__17783));
    LocalMux I__1661 (
            .O(N__17786),
            .I(N__17779));
    LocalMux I__1660 (
            .O(N__17783),
            .I(N__17776));
    InMux I__1659 (
            .O(N__17782),
            .I(N__17773));
    Span4Mux_v I__1658 (
            .O(N__17779),
            .I(N__17770));
    Span4Mux_v I__1657 (
            .O(N__17776),
            .I(N__17767));
    LocalMux I__1656 (
            .O(N__17773),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__1655 (
            .O(N__17770),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__1654 (
            .O(N__17767),
            .I(\c0.FRAME_MATCHER_state_30 ));
    SRMux I__1653 (
            .O(N__17760),
            .I(N__17757));
    LocalMux I__1652 (
            .O(N__17757),
            .I(N__17754));
    Span4Mux_s3_v I__1651 (
            .O(N__17754),
            .I(N__17751));
    Odrv4 I__1650 (
            .O(N__17751),
            .I(\c0.n17283 ));
    CascadeMux I__1649 (
            .O(N__17748),
            .I(N__17744));
    InMux I__1648 (
            .O(N__17747),
            .I(N__17741));
    InMux I__1647 (
            .O(N__17744),
            .I(N__17737));
    LocalMux I__1646 (
            .O(N__17741),
            .I(N__17734));
    InMux I__1645 (
            .O(N__17740),
            .I(N__17731));
    LocalMux I__1644 (
            .O(N__17737),
            .I(N__17726));
    Span4Mux_v I__1643 (
            .O(N__17734),
            .I(N__17726));
    LocalMux I__1642 (
            .O(N__17731),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__1641 (
            .O(N__17726),
            .I(\c0.FRAME_MATCHER_state_3 ));
    InMux I__1640 (
            .O(N__17721),
            .I(N__17718));
    LocalMux I__1639 (
            .O(N__17718),
            .I(N__17713));
    InMux I__1638 (
            .O(N__17717),
            .I(N__17710));
    InMux I__1637 (
            .O(N__17716),
            .I(N__17707));
    Span4Mux_h I__1636 (
            .O(N__17713),
            .I(N__17704));
    LocalMux I__1635 (
            .O(N__17710),
            .I(\c0.FRAME_MATCHER_state_6 ));
    LocalMux I__1634 (
            .O(N__17707),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv4 I__1633 (
            .O(N__17704),
            .I(\c0.FRAME_MATCHER_state_6 ));
    CascadeMux I__1632 (
            .O(N__17697),
            .I(N__17694));
    InMux I__1631 (
            .O(N__17694),
            .I(N__17691));
    LocalMux I__1630 (
            .O(N__17691),
            .I(N__17686));
    InMux I__1629 (
            .O(N__17690),
            .I(N__17683));
    InMux I__1628 (
            .O(N__17689),
            .I(N__17680));
    Span4Mux_v I__1627 (
            .O(N__17686),
            .I(N__17677));
    LocalMux I__1626 (
            .O(N__17683),
            .I(\c0.FRAME_MATCHER_state_7 ));
    LocalMux I__1625 (
            .O(N__17680),
            .I(\c0.FRAME_MATCHER_state_7 ));
    Odrv4 I__1624 (
            .O(N__17677),
            .I(\c0.FRAME_MATCHER_state_7 ));
    CascadeMux I__1623 (
            .O(N__17670),
            .I(\c0.n49_cascade_ ));
    CascadeMux I__1622 (
            .O(N__17667),
            .I(N__17662));
    InMux I__1621 (
            .O(N__17666),
            .I(N__17659));
    InMux I__1620 (
            .O(N__17665),
            .I(N__17656));
    InMux I__1619 (
            .O(N__17662),
            .I(N__17653));
    LocalMux I__1618 (
            .O(N__17659),
            .I(N__17650));
    LocalMux I__1617 (
            .O(N__17656),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__1616 (
            .O(N__17653),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__1615 (
            .O(N__17650),
            .I(\c0.FRAME_MATCHER_state_15 ));
    CascadeMux I__1614 (
            .O(N__17643),
            .I(N__17640));
    InMux I__1613 (
            .O(N__17640),
            .I(N__17637));
    LocalMux I__1612 (
            .O(N__17637),
            .I(N__17633));
    InMux I__1611 (
            .O(N__17636),
            .I(N__17629));
    Span4Mux_h I__1610 (
            .O(N__17633),
            .I(N__17626));
    InMux I__1609 (
            .O(N__17632),
            .I(N__17623));
    LocalMux I__1608 (
            .O(N__17629),
            .I(N__17620));
    Span4Mux_s1_h I__1607 (
            .O(N__17626),
            .I(N__17617));
    LocalMux I__1606 (
            .O(N__17623),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv12 I__1605 (
            .O(N__17620),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__1604 (
            .O(N__17617),
            .I(\c0.FRAME_MATCHER_state_14 ));
    InMux I__1603 (
            .O(N__17610),
            .I(N__17607));
    LocalMux I__1602 (
            .O(N__17607),
            .I(\c0.n50_adj_2353 ));
    CascadeMux I__1601 (
            .O(N__17604),
            .I(N__17600));
    InMux I__1600 (
            .O(N__17603),
            .I(N__17594));
    InMux I__1599 (
            .O(N__17600),
            .I(N__17594));
    InMux I__1598 (
            .O(N__17599),
            .I(N__17591));
    LocalMux I__1597 (
            .O(N__17594),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__1596 (
            .O(N__17591),
            .I(\c0.FRAME_MATCHER_state_10 ));
    InMux I__1595 (
            .O(N__17586),
            .I(N__17583));
    LocalMux I__1594 (
            .O(N__17583),
            .I(\c0.n47 ));
    CascadeMux I__1593 (
            .O(N__17580),
            .I(N__17577));
    InMux I__1592 (
            .O(N__17577),
            .I(N__17572));
    CascadeMux I__1591 (
            .O(N__17576),
            .I(N__17569));
    InMux I__1590 (
            .O(N__17575),
            .I(N__17566));
    LocalMux I__1589 (
            .O(N__17572),
            .I(N__17563));
    InMux I__1588 (
            .O(N__17569),
            .I(N__17560));
    LocalMux I__1587 (
            .O(N__17566),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv4 I__1586 (
            .O(N__17563),
            .I(\c0.FRAME_MATCHER_state_13 ));
    LocalMux I__1585 (
            .O(N__17560),
            .I(\c0.FRAME_MATCHER_state_13 ));
    CascadeMux I__1584 (
            .O(N__17553),
            .I(N__17550));
    InMux I__1583 (
            .O(N__17550),
            .I(N__17546));
    InMux I__1582 (
            .O(N__17549),
            .I(N__17542));
    LocalMux I__1581 (
            .O(N__17546),
            .I(N__17539));
    InMux I__1580 (
            .O(N__17545),
            .I(N__17536));
    LocalMux I__1579 (
            .O(N__17542),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv12 I__1578 (
            .O(N__17539),
            .I(\c0.FRAME_MATCHER_state_25 ));
    LocalMux I__1577 (
            .O(N__17536),
            .I(\c0.FRAME_MATCHER_state_25 ));
    InMux I__1576 (
            .O(N__17529),
            .I(N__17526));
    LocalMux I__1575 (
            .O(N__17526),
            .I(\c0.n48 ));
    InMux I__1574 (
            .O(N__17523),
            .I(N__17514));
    InMux I__1573 (
            .O(N__17522),
            .I(N__17514));
    InMux I__1572 (
            .O(N__17521),
            .I(N__17514));
    LocalMux I__1571 (
            .O(N__17514),
            .I(\c0.FRAME_MATCHER_state_23 ));
    SRMux I__1570 (
            .O(N__17511),
            .I(N__17508));
    LocalMux I__1569 (
            .O(N__17508),
            .I(N__17505));
    Odrv4 I__1568 (
            .O(N__17505),
            .I(\c0.n17275 ));
    SRMux I__1567 (
            .O(N__17502),
            .I(N__17499));
    LocalMux I__1566 (
            .O(N__17499),
            .I(N__17496));
    Sp12to4 I__1565 (
            .O(N__17496),
            .I(N__17493));
    Odrv12 I__1564 (
            .O(N__17493),
            .I(\c0.n3_adj_2293 ));
    SRMux I__1563 (
            .O(N__17490),
            .I(N__17487));
    LocalMux I__1562 (
            .O(N__17487),
            .I(N__17484));
    Span4Mux_s1_h I__1561 (
            .O(N__17484),
            .I(N__17481));
    Odrv4 I__1560 (
            .O(N__17481),
            .I(\c0.n3_adj_2297 ));
    SRMux I__1559 (
            .O(N__17478),
            .I(N__17475));
    LocalMux I__1558 (
            .O(N__17475),
            .I(N__17472));
    Odrv4 I__1557 (
            .O(N__17472),
            .I(\c0.n3_adj_2326 ));
    SRMux I__1556 (
            .O(N__17469),
            .I(N__17466));
    LocalMux I__1555 (
            .O(N__17466),
            .I(N__17463));
    Span4Mux_v I__1554 (
            .O(N__17463),
            .I(N__17460));
    Odrv4 I__1553 (
            .O(N__17460),
            .I(\c0.n3_adj_2313 ));
    SRMux I__1552 (
            .O(N__17457),
            .I(N__17454));
    LocalMux I__1551 (
            .O(N__17454),
            .I(N__17451));
    Odrv4 I__1550 (
            .O(N__17451),
            .I(\c0.n3_adj_2281 ));
    SRMux I__1549 (
            .O(N__17448),
            .I(N__17445));
    LocalMux I__1548 (
            .O(N__17445),
            .I(N__17442));
    Span4Mux_s1_h I__1547 (
            .O(N__17442),
            .I(N__17439));
    Odrv4 I__1546 (
            .O(N__17439),
            .I(\c0.n3_adj_2322 ));
    SRMux I__1545 (
            .O(N__17436),
            .I(N__17433));
    LocalMux I__1544 (
            .O(N__17433),
            .I(N__17430));
    Odrv4 I__1543 (
            .O(N__17430),
            .I(\c0.n3_adj_2311 ));
    SRMux I__1542 (
            .O(N__17427),
            .I(N__17424));
    LocalMux I__1541 (
            .O(N__17424),
            .I(N__17421));
    Span4Mux_s1_h I__1540 (
            .O(N__17421),
            .I(N__17418));
    Odrv4 I__1539 (
            .O(N__17418),
            .I(\c0.n3_adj_2307 ));
    InMux I__1538 (
            .O(N__17415),
            .I(N__17412));
    LocalMux I__1537 (
            .O(N__17412),
            .I(N__17409));
    Odrv4 I__1536 (
            .O(N__17409),
            .I(\c0.n42 ));
    SRMux I__1535 (
            .O(N__17406),
            .I(N__17403));
    LocalMux I__1534 (
            .O(N__17403),
            .I(N__17400));
    Odrv4 I__1533 (
            .O(N__17400),
            .I(\c0.n3_adj_2299 ));
    SRMux I__1532 (
            .O(N__17397),
            .I(N__17394));
    LocalMux I__1531 (
            .O(N__17394),
            .I(N__17391));
    Odrv12 I__1530 (
            .O(N__17391),
            .I(\c0.n8_adj_2258 ));
    CascadeMux I__1529 (
            .O(N__17388),
            .I(\c0.n39_cascade_ ));
    CascadeMux I__1528 (
            .O(N__17385),
            .I(\c0.n48_adj_2383_cascade_ ));
    InMux I__1527 (
            .O(N__17382),
            .I(N__17379));
    LocalMux I__1526 (
            .O(N__17379),
            .I(\c0.n40 ));
    InMux I__1525 (
            .O(N__17376),
            .I(N__17373));
    LocalMux I__1524 (
            .O(N__17373),
            .I(\c0.n41 ));
    InMux I__1523 (
            .O(N__17370),
            .I(N__17367));
    LocalMux I__1522 (
            .O(N__17367),
            .I(\c0.n43_adj_2384 ));
    CascadeMux I__1521 (
            .O(N__17364),
            .I(\c0.n17713_cascade_ ));
    SRMux I__1520 (
            .O(N__17361),
            .I(N__17358));
    LocalMux I__1519 (
            .O(N__17358),
            .I(N__17355));
    Span4Mux_s3_v I__1518 (
            .O(N__17355),
            .I(N__17352));
    Odrv4 I__1517 (
            .O(N__17352),
            .I(\c0.n8_adj_2234 ));
    SRMux I__1516 (
            .O(N__17349),
            .I(N__17346));
    LocalMux I__1515 (
            .O(N__17346),
            .I(N__17343));
    Odrv4 I__1514 (
            .O(N__17343),
            .I(\c0.n17281 ));
    SRMux I__1513 (
            .O(N__17340),
            .I(N__17337));
    LocalMux I__1512 (
            .O(N__17337),
            .I(N__17334));
    Span4Mux_s1_h I__1511 (
            .O(N__17334),
            .I(N__17331));
    Odrv4 I__1510 (
            .O(N__17331),
            .I(\c0.n17259 ));
    SRMux I__1509 (
            .O(N__17328),
            .I(N__17325));
    LocalMux I__1508 (
            .O(N__17325),
            .I(\c0.n17261 ));
    SRMux I__1507 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__1506 (
            .O(N__17319),
            .I(N__17316));
    Span4Mux_s2_h I__1505 (
            .O(N__17316),
            .I(N__17313));
    Odrv4 I__1504 (
            .O(N__17313),
            .I(\c0.n13900 ));
    InMux I__1503 (
            .O(N__17310),
            .I(N__17305));
    InMux I__1502 (
            .O(N__17309),
            .I(N__17300));
    InMux I__1501 (
            .O(N__17308),
            .I(N__17300));
    LocalMux I__1500 (
            .O(N__17305),
            .I(\c0.FRAME_MATCHER_state_8 ));
    LocalMux I__1499 (
            .O(N__17300),
            .I(\c0.FRAME_MATCHER_state_8 ));
    SRMux I__1498 (
            .O(N__17295),
            .I(N__17292));
    LocalMux I__1497 (
            .O(N__17292),
            .I(N__17289));
    Span4Mux_v I__1496 (
            .O(N__17289),
            .I(N__17286));
    Odrv4 I__1495 (
            .O(N__17286),
            .I(\c0.n8_adj_2257 ));
    SRMux I__1494 (
            .O(N__17283),
            .I(N__17280));
    LocalMux I__1493 (
            .O(N__17280),
            .I(N__17277));
    Span4Mux_s2_h I__1492 (
            .O(N__17277),
            .I(N__17274));
    Odrv4 I__1491 (
            .O(N__17274),
            .I(\c0.n17263 ));
    CascadeMux I__1490 (
            .O(N__17271),
            .I(N__17268));
    InMux I__1489 (
            .O(N__17268),
            .I(N__17265));
    LocalMux I__1488 (
            .O(N__17265),
            .I(N__17260));
    InMux I__1487 (
            .O(N__17264),
            .I(N__17257));
    InMux I__1486 (
            .O(N__17263),
            .I(N__17254));
    Span4Mux_v I__1485 (
            .O(N__17260),
            .I(N__17251));
    LocalMux I__1484 (
            .O(N__17257),
            .I(N__17248));
    LocalMux I__1483 (
            .O(N__17254),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv4 I__1482 (
            .O(N__17251),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv12 I__1481 (
            .O(N__17248),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__1480 (
            .O(N__17241),
            .I(N__17238));
    LocalMux I__1479 (
            .O(N__17238),
            .I(N__17235));
    Span4Mux_s1_h I__1478 (
            .O(N__17235),
            .I(N__17232));
    Odrv4 I__1477 (
            .O(N__17232),
            .I(\c0.n17265 ));
    InMux I__1476 (
            .O(N__17229),
            .I(N__17226));
    LocalMux I__1475 (
            .O(N__17226),
            .I(N__17221));
    InMux I__1474 (
            .O(N__17225),
            .I(N__17218));
    InMux I__1473 (
            .O(N__17224),
            .I(N__17215));
    Span4Mux_h I__1472 (
            .O(N__17221),
            .I(N__17210));
    LocalMux I__1471 (
            .O(N__17218),
            .I(N__17210));
    LocalMux I__1470 (
            .O(N__17215),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__1469 (
            .O(N__17210),
            .I(\c0.FRAME_MATCHER_state_12 ));
    SRMux I__1468 (
            .O(N__17205),
            .I(N__17202));
    LocalMux I__1467 (
            .O(N__17202),
            .I(N__17199));
    Sp12to4 I__1466 (
            .O(N__17199),
            .I(N__17196));
    Odrv12 I__1465 (
            .O(N__17196),
            .I(\c0.n17267 ));
    SRMux I__1464 (
            .O(N__17193),
            .I(N__17190));
    LocalMux I__1463 (
            .O(N__17190),
            .I(\c0.n17269 ));
    SRMux I__1462 (
            .O(N__17187),
            .I(N__17184));
    LocalMux I__1461 (
            .O(N__17184),
            .I(N__17181));
    Sp12to4 I__1460 (
            .O(N__17181),
            .I(N__17178));
    Odrv12 I__1459 (
            .O(N__17178),
            .I(\c0.n17303 ));
    SRMux I__1458 (
            .O(N__17175),
            .I(N__17172));
    LocalMux I__1457 (
            .O(N__17172),
            .I(N__17169));
    Span4Mux_s1_h I__1456 (
            .O(N__17169),
            .I(N__17166));
    Odrv4 I__1455 (
            .O(N__17166),
            .I(\c0.n17271 ));
    CascadeMux I__1454 (
            .O(N__17163),
            .I(n10429_cascade_));
    InMux I__1453 (
            .O(N__17160),
            .I(N__17157));
    LocalMux I__1452 (
            .O(N__17157),
            .I(n12965));
    InMux I__1451 (
            .O(N__17154),
            .I(N__17151));
    LocalMux I__1450 (
            .O(N__17151),
            .I(n242));
    CascadeMux I__1449 (
            .O(N__17148),
            .I(n12965_cascade_));
    InMux I__1448 (
            .O(N__17145),
            .I(N__17142));
    LocalMux I__1447 (
            .O(N__17142),
            .I(n10429));
    InMux I__1446 (
            .O(N__17139),
            .I(N__17136));
    LocalMux I__1445 (
            .O(N__17136),
            .I(N__17133));
    Odrv12 I__1444 (
            .O(N__17133),
            .I(n8_adj_2541));
    InMux I__1443 (
            .O(N__17130),
            .I(N__17127));
    LocalMux I__1442 (
            .O(N__17127),
            .I(n18_adj_2539));
    CascadeMux I__1441 (
            .O(N__17124),
            .I(n21_adj_2538_cascade_));
    InMux I__1440 (
            .O(N__17121),
            .I(N__17118));
    LocalMux I__1439 (
            .O(N__17118),
            .I(n15_adj_2540));
    CascadeMux I__1438 (
            .O(N__17115),
            .I(\c0.n4_adj_2271_cascade_ ));
    InMux I__1437 (
            .O(N__17112),
            .I(N__17109));
    LocalMux I__1436 (
            .O(N__17109),
            .I(\c0.n2_adj_2341 ));
    CascadeMux I__1435 (
            .O(N__17106),
            .I(\c0.n2_adj_2341_cascade_ ));
    InMux I__1434 (
            .O(N__17103),
            .I(N__17100));
    LocalMux I__1433 (
            .O(N__17100),
            .I(\c0.n10425 ));
    CascadeMux I__1432 (
            .O(N__17097),
            .I(N__17094));
    InMux I__1431 (
            .O(N__17094),
            .I(N__17091));
    LocalMux I__1430 (
            .O(N__17091),
            .I(\c0.n10465 ));
    IoInMux I__1429 (
            .O(N__17088),
            .I(N__17085));
    LocalMux I__1428 (
            .O(N__17085),
            .I(N__17082));
    IoSpan4Mux I__1427 (
            .O(N__17082),
            .I(N__17079));
    IoSpan4Mux I__1426 (
            .O(N__17079),
            .I(N__17076));
    IoSpan4Mux I__1425 (
            .O(N__17076),
            .I(N__17073));
    Odrv4 I__1424 (
            .O(N__17073),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(n16585),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(n16593),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(n16601),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(n16554),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(n16562),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(n16570),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\control.n16654 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\c0.tx2.n16546 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\c0.tx.n16531 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\c0.n16641 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(\c0.n16493 ),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\c0.n16501 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\c0.n16509 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(n16616),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(n16624),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(n16632),
            .carryinitout(bfn_6_24_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__17088),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i4_LC_1_1_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_1_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_1_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__20308),
            .in2(_gnd_net_),
            .in3(N__20091),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49785),
            .ce(),
            .sr(N__17361));
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_2_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_1_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__17263),
            .in2(_gnd_net_),
            .in3(N__20065),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49769),
            .ce(),
            .sr(N__17241));
    defparam \c0.FRAME_MATCHER_state_i12_LC_1_3_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_1_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_1_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__17224),
            .in2(_gnd_net_),
            .in3(N__20041),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49756),
            .ce(),
            .sr(N__17205));
    defparam \c0.FRAME_MATCHER_state_i15_LC_1_4_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_1_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_1_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__17665),
            .in2(_gnd_net_),
            .in3(N__19991),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49743),
            .ce(),
            .sr(N__17175));
    defparam \c0.i1_4_lut_adj_507_LC_1_5_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_507_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_507_LC_1_5_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.i1_4_lut_adj_507_LC_1_5_0  (
            .in0(N__18596),
            .in1(N__17112),
            .in2(N__17097),
            .in3(N__21297),
            .lcout(\c0.n4_adj_2271 ),
            .ltout(\c0.n4_adj_2271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_5_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_5_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_1_5_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_1_5_1  (
            .in0(N__17309),
            .in1(_gnd_net_),
            .in2(N__17115),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49731),
            .ce(),
            .sr(N__17295));
    defparam \c0.i16_4_lut_LC_1_5_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_1_5_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_LC_1_5_2  (
            .in0(N__17225),
            .in1(N__17264),
            .in2(N__17793),
            .in3(N__17308),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_620_LC_1_5_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_620_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_620_LC_1_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_620_LC_1_5_3  (
            .in0(N__30517),
            .in1(N__21915),
            .in2(N__28712),
            .in3(N__21505),
            .lcout(\c0.n2_adj_2341 ),
            .ltout(\c0.n2_adj_2341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_553_LC_1_5_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_553_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_553_LC_1_5_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.i1_4_lut_adj_553_LC_1_5_4  (
            .in0(N__21916),
            .in1(N__18598),
            .in2(N__17106),
            .in3(N__17103),
            .lcout(\c0.n4_adj_2349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_550_LC_1_5_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_550_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_550_LC_1_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_550_LC_1_5_5  (
            .in0(N__18156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21504),
            .lcout(\c0.n10425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_1_5_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_1_5_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_708_LC_1_5_6  (
            .in0(N__21503),
            .in1(N__18160),
            .in2(_gnd_net_),
            .in3(N__21203),
            .lcout(\c0.n10465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_1_5_7.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_1_5_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 i2_3_lut_4_lut_LC_1_5_7 (
            .in0(N__21204),
            .in1(N__18597),
            .in2(N__18162),
            .in3(N__21506),
            .lcout(n8_adj_2541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_1_6_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_1_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_1_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__17740),
            .in2(_gnd_net_),
            .in3(N__19992),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49720),
            .ce(),
            .sr(N__17349));
    defparam \c0.FRAME_MATCHER_state_i6_LC_1_7_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_1_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_1_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__17717),
            .in2(_gnd_net_),
            .in3(N__20055),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49707),
            .ce(),
            .sr(N__17328));
    defparam \c0.FRAME_MATCHER_state_i5_LC_1_8_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_1_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_1_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__20371),
            .in2(_gnd_net_),
            .in3(N__20087),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(N__17340));
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_1_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_686_LC_1_9_0 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_686_LC_1_9_0  (
            .in0(N__23338),
            .in1(_gnd_net_),
            .in2(N__25626),
            .in3(N__23445),
            .lcout(n242),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_1_9_1.C_ON=1'b0;
    defparam i1_3_lut_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_1_9_1.LUT_INIT=16'b1100110010001000;
    LogicCell40 i1_3_lut_LC_1_9_1 (
            .in0(N__19023),
            .in1(N__19005),
            .in2(_gnd_net_),
            .in3(N__17160),
            .lcout(n18_adj_2539),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_597_LC_1_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_597_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_597_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_597_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__21195),
            .in2(_gnd_net_),
            .in3(N__21453),
            .lcout(n10429),
            .ltout(n10429_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_450_LC_1_9_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_450_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_450_LC_1_9_3 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_450_LC_1_9_3  (
            .in0(N__20982),
            .in1(N__18173),
            .in2(N__17163),
            .in3(N__20815),
            .lcout(n12965),
            .ltout(n12965_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_827_LC_1_9_4.C_ON=1'b0;
    defparam i1_4_lut_adj_827_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_827_LC_1_9_4.LUT_INIT=16'b1010000010101000;
    LogicCell40 i1_4_lut_adj_827_LC_1_9_4 (
            .in0(N__18942),
            .in1(N__17154),
            .in2(N__17148),
            .in3(N__20983),
            .lcout(n15_adj_2540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_1_9_5.C_ON=1'b0;
    defparam i1_4_lut_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_1_9_5.LUT_INIT=16'b1100110010000000;
    LogicCell40 i1_4_lut_LC_1_9_5 (
            .in0(N__17145),
            .in1(N__18174),
            .in2(N__17943),
            .in3(N__17139),
            .lcout(),
            .ltout(n21_adj_2538_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_1_9_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i1_LC_1_9_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_1_9_6  (
            .in0(N__17130),
            .in1(N__18735),
            .in2(N__17124),
            .in3(N__17121),
            .lcout(\c0.FRAME_MATCHER_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_779_LC_1_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_779_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_779_LC_1_9_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_779_LC_1_9_7  (
            .in0(N__20981),
            .in1(N__23337),
            .in2(_gnd_net_),
            .in3(N__20814),
            .lcout(n8_adj_2498),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_1_10_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i12_LC_1_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_1_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__24565),
            .in2(_gnd_net_),
            .in3(N__19233),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49685),
            .ce(),
            .sr(N__17448));
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_11_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_11_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__24586),
            .in2(_gnd_net_),
            .in3(N__19161),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49680),
            .ce(),
            .sr(N__21552));
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_12_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__24626),
            .in2(_gnd_net_),
            .in3(N__19602),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49675),
            .ce(),
            .sr(N__17436));
    defparam \c0.FRAME_MATCHER_i_i17_LC_1_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i17_LC_1_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_1_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__24627),
            .in2(_gnd_net_),
            .in3(N__19482),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49671),
            .ce(),
            .sr(N__17427));
    defparam \c0.FRAME_MATCHER_i_i24_LC_1_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i24_LC_1_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_1_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__24628),
            .in2(_gnd_net_),
            .in3(N__19770),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49668),
            .ce(),
            .sr(N__17502));
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_1_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__24629),
            .in2(_gnd_net_),
            .in3(N__19878),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(N__17490));
    defparam \c0.FRAME_MATCHER_state_i27_LC_2_1_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_2_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_2_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_2_1_0  (
            .in0(_gnd_net_),
            .in1(N__17821),
            .in2(_gnd_net_),
            .in3(N__20495),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49798),
            .ce(),
            .sr(N__17805));
    defparam \c0.FRAME_MATCHER_state_i14_LC_2_2_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_2_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_2_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__17632),
            .in2(_gnd_net_),
            .in3(N__20098),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49786),
            .ce(),
            .sr(N__17187));
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_3_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__17549),
            .in2(_gnd_net_),
            .in3(N__20097),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49770),
            .ce(),
            .sr(N__17322));
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_4_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__17575),
            .in2(_gnd_net_),
            .in3(N__20020),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49757),
            .ce(),
            .sr(N__17193));
    defparam \c0.i1_2_lut_4_lut_adj_647_LC_2_5_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_647_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_647_LC_2_5_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_647_LC_2_5_0  (
            .in0(N__18429),
            .in1(N__18027),
            .in2(N__17604),
            .in3(N__19136),
            .lcout(\c0.n17263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i10_LC_2_5_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_2_5_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_2_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__19990),
            .in2(_gnd_net_),
            .in3(N__17603),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49744),
            .ce(),
            .sr(N__17283));
    defparam \c0.i1_2_lut_4_lut_adj_650_LC_2_5_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_650_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_650_LC_2_5_2 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_650_LC_2_5_2  (
            .in0(N__18430),
            .in1(N__18028),
            .in2(N__17271),
            .in3(N__19137),
            .lcout(\c0.n17265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_657_LC_2_5_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_657_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_657_LC_2_5_3 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_657_LC_2_5_3  (
            .in0(N__19138),
            .in1(N__17229),
            .in2(N__18058),
            .in3(N__18431),
            .lcout(\c0.n17267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_659_LC_2_5_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_659_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_659_LC_2_5_4 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_659_LC_2_5_4  (
            .in0(N__18432),
            .in1(N__18032),
            .in2(N__17580),
            .in3(N__19139),
            .lcout(\c0.n17269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_663_LC_2_5_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_663_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_663_LC_2_5_5 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_663_LC_2_5_5  (
            .in0(N__19140),
            .in1(N__17636),
            .in2(N__18059),
            .in3(N__18433),
            .lcout(\c0.n17303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_669_LC_2_5_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_669_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_669_LC_2_5_6 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_669_LC_2_5_6  (
            .in0(N__18434),
            .in1(N__18036),
            .in2(N__17667),
            .in3(N__19141),
            .lcout(\c0.n17271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_673_LC_2_5_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_673_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_673_LC_2_5_7 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_673_LC_2_5_7  (
            .in0(N__19142),
            .in1(N__20349),
            .in2(N__18060),
            .in3(N__18435),
            .lcout(\c0.n8_adj_2254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_548_LC_2_6_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_548_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_548_LC_2_6_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.i1_4_lut_adj_548_LC_2_6_0  (
            .in0(N__19003),
            .in1(N__18888),
            .in2(N__18216),
            .in3(N__22567),
            .lcout(\c0.n17713 ),
            .ltout(\c0.n17713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_442_LC_2_6_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_442_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_442_LC_2_6_1 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_442_LC_2_6_1  (
            .in0(N__22569),
            .in1(N__20318),
            .in2(N__17364),
            .in3(N__18380),
            .lcout(\c0.n8_adj_2234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_2_6_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_2_6_2 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_2_6_2  (
            .in0(N__18379),
            .in1(N__18016),
            .in2(N__17748),
            .in3(N__22568),
            .lcout(\c0.n17281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_639_LC_2_6_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_639_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_639_LC_2_6_3 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_639_LC_2_6_3  (
            .in0(N__19145),
            .in1(N__17689),
            .in2(N__18056),
            .in3(N__18383),
            .lcout(\c0.n8_adj_2258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_446_LC_2_6_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_446_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_446_LC_2_6_4 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_446_LC_2_6_4  (
            .in0(N__18381),
            .in1(N__18017),
            .in2(N__20382),
            .in3(N__22570),
            .lcout(\c0.n17259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_638_LC_2_6_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_638_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_638_LC_2_6_5 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_638_LC_2_6_5  (
            .in0(N__19144),
            .in1(N__17716),
            .in2(N__18055),
            .in3(N__18382),
            .lcout(\c0.n17261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11136_2_lut_4_lut_LC_2_6_6 .C_ON=1'b0;
    defparam \c0.i11136_2_lut_4_lut_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11136_2_lut_4_lut_LC_2_6_6 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i11136_2_lut_4_lut_LC_2_6_6  (
            .in0(N__18378),
            .in1(N__18015),
            .in2(N__17553),
            .in3(N__19143),
            .lcout(\c0.n13900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_640_LC_2_6_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_640_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_640_LC_2_6_7 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_640_LC_2_6_7  (
            .in0(N__19146),
            .in1(N__17310),
            .in2(N__18057),
            .in3(N__18384),
            .lcout(\c0.n8_adj_2257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_7_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_2_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__17690),
            .in2(_gnd_net_),
            .in3(N__20101),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49721),
            .ce(),
            .sr(N__17397));
    defparam \c0.FRAME_MATCHER_state_i9_LC_2_8_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_2_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_2_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_2_8_0  (
            .in0(N__20102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18082),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49708),
            .ce(),
            .sr(N__17955));
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_9_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__24502),
            .in2(_gnd_net_),
            .in3(N__19206),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(N__18282));
    defparam \c0.FRAME_MATCHER_i_i20_LC_2_10_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i20_LC_2_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_2_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_2_10_0  (
            .in0(N__24503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19452),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49692),
            .ce(),
            .sr(N__18108));
    defparam \c0.i14_4_lut_adj_607_LC_2_11_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_607_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_607_LC_2_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_607_LC_2_11_0  (
            .in0(N__20229),
            .in1(N__22222),
            .in2(N__21046),
            .in3(N__19371),
            .lcout(),
            .ltout(\c0.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_2_11_1 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_2_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i23_4_lut_LC_2_11_1  (
            .in0(N__17415),
            .in1(N__17382),
            .in2(N__17388),
            .in3(N__17376),
            .lcout(),
            .ltout(\c0.n48_adj_2383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_612_LC_2_11_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_612_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_612_LC_2_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_612_LC_2_11_2  (
            .in0(N__21947),
            .in1(N__17370),
            .in2(N__17385),
            .in3(N__22083),
            .lcout(\c0.n10522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_605_LC_2_11_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_605_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_605_LC_2_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_605_LC_2_11_3  (
            .in0(N__19746),
            .in1(N__22439),
            .in2(N__22179),
            .in3(N__19851),
            .lcout(\c0.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_606_LC_2_11_4 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_606_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_606_LC_2_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_606_LC_2_11_4  (
            .in0(N__19623),
            .in1(N__19513),
            .in2(N__24704),
            .in3(N__19317),
            .lcout(\c0.n41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_611_LC_2_12_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_611_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_611_LC_2_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_611_LC_2_12_0  (
            .in0(N__21093),
            .in1(N__19566),
            .in2(N__24380),
            .in3(N__20751),
            .lcout(\c0.n43_adj_2384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i30_LC_2_12_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i30_LC_2_12_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_2_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__24567),
            .in2(_gnd_net_),
            .in3(N__20271),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49681),
            .ce(),
            .sr(N__17457));
    defparam \c0.select_284_Select_30_i3_2_lut_3_lut_4_lut_LC_2_12_2 .C_ON=1'b0;
    defparam \c0.select_284_Select_30_i3_2_lut_3_lut_4_lut_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_30_i3_2_lut_3_lut_4_lut_LC_2_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.select_284_Select_30_i3_2_lut_3_lut_4_lut_LC_2_12_2  (
            .in0(N__21520),
            .in1(N__20752),
            .in2(N__21924),
            .in3(N__21670),
            .lcout(\c0.n3_adj_2281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_14_i3_2_lut_3_lut_4_lut_LC_2_12_3 .C_ON=1'b0;
    defparam \c0.select_284_Select_14_i3_2_lut_3_lut_4_lut_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_14_i3_2_lut_3_lut_4_lut_LC_2_12_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_14_i3_2_lut_3_lut_4_lut_LC_2_12_3  (
            .in0(N__21664),
            .in1(N__21902),
            .in2(N__21108),
            .in3(N__21516),
            .lcout(\c0.n3_adj_2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_13_i3_2_lut_3_lut_4_lut_LC_2_12_4 .C_ON=1'b0;
    defparam \c0.select_284_Select_13_i3_2_lut_3_lut_4_lut_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_13_i3_2_lut_3_lut_4_lut_LC_2_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.select_284_Select_13_i3_2_lut_3_lut_4_lut_LC_2_12_4  (
            .in0(N__21515),
            .in1(N__24379),
            .in2(N__21922),
            .in3(N__21663),
            .lcout(\c0.n3_adj_2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_12_i3_2_lut_3_lut_4_lut_LC_2_12_5 .C_ON=1'b0;
    defparam \c0.select_284_Select_12_i3_2_lut_3_lut_4_lut_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_12_i3_2_lut_3_lut_4_lut_LC_2_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_12_i3_2_lut_3_lut_4_lut_LC_2_12_5  (
            .in0(N__21665),
            .in1(N__21903),
            .in2(N__22626),
            .in3(N__21517),
            .lcout(\c0.n3_adj_2322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_15_i3_2_lut_3_lut_4_lut_LC_2_12_6 .C_ON=1'b0;
    defparam \c0.select_284_Select_15_i3_2_lut_3_lut_4_lut_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_15_i3_2_lut_3_lut_4_lut_LC_2_12_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_15_i3_2_lut_3_lut_4_lut_LC_2_12_6  (
            .in0(N__21519),
            .in1(N__21669),
            .in2(N__21923),
            .in3(N__19630),
            .lcout(\c0.n3_adj_2311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_17_i3_2_lut_3_lut_4_lut_LC_2_12_7 .C_ON=1'b0;
    defparam \c0.select_284_Select_17_i3_2_lut_3_lut_4_lut_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_17_i3_2_lut_3_lut_4_lut_LC_2_12_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_17_i3_2_lut_3_lut_4_lut_LC_2_12_7  (
            .in0(N__19512),
            .in1(N__21904),
            .in2(N__21708),
            .in3(N__21518),
            .lcout(\c0.n3_adj_2307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_602_LC_2_13_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_602_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_602_LC_2_13_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_602_LC_2_13_0  (
            .in0(N__19905),
            .in1(N__19797),
            .in2(N__20717),
            .in3(N__19407),
            .lcout(\c0.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i21_LC_2_13_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i21_LC_2_13_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_2_13_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_2_13_1  (
            .in0(N__24569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19392),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49676),
            .ce(),
            .sr(N__17406));
    defparam \c0.select_284_Select_21_i3_2_lut_3_lut_4_lut_LC_2_13_2 .C_ON=1'b0;
    defparam \c0.select_284_Select_21_i3_2_lut_3_lut_4_lut_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_21_i3_2_lut_3_lut_4_lut_LC_2_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_21_i3_2_lut_3_lut_4_lut_LC_2_13_2  (
            .in0(N__21531),
            .in1(N__19408),
            .in2(N__21715),
            .in3(N__21885),
            .lcout(\c0.n3_adj_2299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_24_i3_2_lut_3_lut_4_lut_LC_2_13_3 .C_ON=1'b0;
    defparam \c0.select_284_Select_24_i3_2_lut_3_lut_4_lut_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_24_i3_2_lut_3_lut_4_lut_LC_2_13_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_24_i3_2_lut_3_lut_4_lut_LC_2_13_3  (
            .in0(N__21881),
            .in1(N__21684),
            .in2(N__19805),
            .in3(N__21527),
            .lcout(\c0.n3_adj_2293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_22_i3_2_lut_3_lut_4_lut_LC_2_13_4 .C_ON=1'b0;
    defparam \c0.select_284_Select_22_i3_2_lut_3_lut_4_lut_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_22_i3_2_lut_3_lut_4_lut_LC_2_13_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_22_i3_2_lut_3_lut_4_lut_LC_2_13_4  (
            .in0(N__21528),
            .in1(N__19919),
            .in2(N__21713),
            .in3(N__21883),
            .lcout(\c0.n3_adj_2297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_29_i3_2_lut_3_lut_4_lut_LC_2_13_5 .C_ON=1'b0;
    defparam \c0.select_284_Select_29_i3_2_lut_3_lut_4_lut_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_29_i3_2_lut_3_lut_4_lut_LC_2_13_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.select_284_Select_29_i3_2_lut_3_lut_4_lut_LC_2_13_5  (
            .in0(N__21886),
            .in1(N__20712),
            .in2(N__21543),
            .in3(N__21695),
            .lcout(\c0.n3_adj_2283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_10_i3_2_lut_3_lut_4_lut_LC_2_13_6 .C_ON=1'b0;
    defparam \c0.select_284_Select_10_i3_2_lut_3_lut_4_lut_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_10_i3_2_lut_3_lut_4_lut_LC_2_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_10_i3_2_lut_3_lut_4_lut_LC_2_13_6  (
            .in0(N__21530),
            .in1(N__22221),
            .in2(N__21714),
            .in3(N__21884),
            .lcout(\c0.n3_adj_2326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_11_i3_2_lut_3_lut_4_lut_LC_2_13_7 .C_ON=1'b0;
    defparam \c0.select_284_Select_11_i3_2_lut_3_lut_4_lut_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_11_i3_2_lut_3_lut_4_lut_LC_2_13_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_11_i3_2_lut_3_lut_4_lut_LC_2_13_7  (
            .in0(N__21882),
            .in1(N__21685),
            .in2(N__22071),
            .in3(N__21529),
            .lcout(\c0.n3_adj_2324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_2_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i25_LC_2_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_2_14_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_2_14_0  (
            .in0(N__24585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19701),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(N__18234));
    defparam \c0.FRAME_MATCHER_i_i10_LC_2_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i10_LC_2_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_2_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_2_15_0  (
            .in0(N__24623),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19251),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49669),
            .ce(),
            .sr(N__17478));
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_2_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__24625),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49667),
            .ce(),
            .sr(N__17469));
    defparam \c0.FRAME_MATCHER_state_i30_LC_3_1_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_3_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_3_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_3_1_0  (
            .in0(_gnd_net_),
            .in1(N__17782),
            .in2(_gnd_net_),
            .in3(N__20496),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49810),
            .ce(),
            .sr(N__17760));
    defparam \c0.FRAME_MATCHER_state_i24_LC_3_2_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_3_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_3_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_3_2_0  (
            .in0(_gnd_net_),
            .in1(N__18506),
            .in2(_gnd_net_),
            .in3(N__20100),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49799),
            .ce(),
            .sr(N__17847));
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_3_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_3_3_0  (
            .in0(_gnd_net_),
            .in1(N__18683),
            .in2(_gnd_net_),
            .in3(N__20099),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49787),
            .ce(),
            .sr(N__18663));
    defparam \c0.i20_4_lut_LC_3_4_0 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_3_4_0 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_3_4_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20_4_lut_LC_3_4_0  (
            .in0(N__17747),
            .in1(N__17721),
            .in2(N__17697),
            .in3(N__20132),
            .lcout(),
            .ltout(\c0.n49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_3_4_1 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_3_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_3_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i27_4_lut_LC_3_4_1  (
            .in0(N__17610),
            .in1(N__17529),
            .in2(N__17670),
            .in3(N__17586),
            .lcout(\c0.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_3_4_2 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_3_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_3_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i21_4_lut_LC_3_4_2  (
            .in0(N__17666),
            .in1(N__18089),
            .in2(N__17643),
            .in3(N__18545),
            .lcout(\c0.n50_adj_2353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_3_4_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_3_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_3_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_LC_3_4_3  (
            .in0(N__17912),
            .in1(N__17599),
            .in2(N__17834),
            .in3(N__17521),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_3_4_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_3_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_3_4_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_LC_3_4_4  (
            .in0(N__17872),
            .in1(N__18679),
            .in2(N__17576),
            .in3(N__17545),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i23_LC_3_4_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_3_4_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_3_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_3_4_5  (
            .in0(_gnd_net_),
            .in1(N__17523),
            .in2(_gnd_net_),
            .in3(N__20096),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49771),
            .ce(),
            .sr(N__17511));
    defparam \c0.i1_2_lut_adj_497_LC_3_4_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_497_LC_3_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_497_LC_3_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_497_LC_3_4_6  (
            .in0(N__17522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18705),
            .lcout(\c0.n17275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_697_LC_3_5_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_697_LC_3_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_697_LC_3_5_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_697_LC_3_5_0  (
            .in0(N__18422),
            .in1(N__18042),
            .in2(N__17877),
            .in3(N__19129),
            .lcout(\c0.n8_adj_2252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i17_LC_3_5_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_3_5_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_3_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_3_5_1  (
            .in0(_gnd_net_),
            .in1(N__17876),
            .in2(_gnd_net_),
            .in3(N__20042),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49759),
            .ce(),
            .sr(N__17859));
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_3_5_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_3_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_698_LC_3_5_2 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_698_LC_3_5_2  (
            .in0(N__18423),
            .in1(N__18043),
            .in2(N__18510),
            .in3(N__19130),
            .lcout(\c0.n8_adj_2246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_5_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_5_3 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_720_LC_3_5_3  (
            .in0(N__19131),
            .in1(N__18546),
            .in2(N__18061),
            .in3(N__18424),
            .lcout(\c0.n8_adj_2245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_3_5_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_3_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_3_5_4 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_732_LC_3_5_4  (
            .in0(N__18425),
            .in1(N__18047),
            .in2(N__17835),
            .in3(N__19132),
            .lcout(\c0.n17277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_736_LC_3_5_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_736_LC_3_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_736_LC_3_5_5 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_736_LC_3_5_5  (
            .in0(N__19133),
            .in1(N__18653),
            .in2(N__18062),
            .in3(N__18426),
            .lcout(\c0.n17299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_742_LC_3_5_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_742_LC_3_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_742_LC_3_5_6 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_742_LC_3_5_6  (
            .in0(N__18427),
            .in1(N__18051),
            .in2(N__20406),
            .in3(N__19134),
            .lcout(\c0.n8_adj_2244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_745_LC_3_5_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_745_LC_3_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_745_LC_3_5_7 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_745_LC_3_5_7  (
            .in0(N__19135),
            .in1(N__17792),
            .in2(N__18063),
            .in3(N__18428),
            .lcout(\c0.n17283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_749_LC_3_6_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_749_LC_3_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_749_LC_3_6_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_749_LC_3_6_0  (
            .in0(N__18377),
            .in1(N__18040),
            .in2(N__17913),
            .in3(N__19088),
            .lcout(\c0.n17279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_451_LC_3_6_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_451_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_451_LC_3_6_1 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \c0.i1_4_lut_adj_451_LC_3_6_1  (
            .in0(N__30492),
            .in1(N__25052),
            .in2(N__29943),
            .in3(N__30114),
            .lcout(n17694),
            .ltout(n17694_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_3_6_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_3_6_2 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_755_LC_3_6_2  (
            .in0(N__25053),
            .in1(N__46151),
            .in2(N__17916),
            .in3(N__33057),
            .lcout(\c0.n4_adj_2231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_3_6_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_3_6_3 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_765_LC_3_6_3  (
            .in0(N__33060),
            .in1(N__25056),
            .in2(N__25114),
            .in3(N__49107),
            .lcout(\c0.n4_adj_2216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_3_6_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_3_6_4 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_760_LC_3_6_4  (
            .in0(N__25054),
            .in1(N__25100),
            .in2(N__48570),
            .in3(N__33058),
            .lcout(\c0.n4_adj_2226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_3_6_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_3_6_5 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_761_LC_3_6_5  (
            .in0(N__33059),
            .in1(N__25055),
            .in2(N__25113),
            .in3(N__48017),
            .lcout(\c0.n4_adj_2225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i31_LC_3_6_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_3_6_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_3_6_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_3_6_6  (
            .in0(N__17911),
            .in1(_gnd_net_),
            .in2(N__20498),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49745),
            .ce(),
            .sr(N__17892));
    defparam \c0.i1_2_lut_4_lut_adj_768_LC_3_6_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_768_LC_3_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_768_LC_3_6_7 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_768_LC_3_6_7  (
            .in0(N__33061),
            .in1(N__25057),
            .in2(N__25115),
            .in3(N__48928),
            .lcout(\c0.n4_adj_2204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10973_2_lut_LC_3_7_0 .C_ON=1'b0;
    defparam \c0.i10973_2_lut_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10973_2_lut_LC_3_7_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i10973_2_lut_LC_3_7_0  (
            .in0(_gnd_net_),
            .in1(N__30011),
            .in2(_gnd_net_),
            .in3(N__19086),
            .lcout(),
            .ltout(FRAME_MATCHER_state_31_N_1406_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_829_LC_3_7_1.C_ON=1'b0;
    defparam i2_4_lut_adj_829_LC_3_7_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_829_LC_3_7_1.LUT_INIT=16'b1110110010100000;
    LogicCell40 i2_4_lut_adj_829_LC_3_7_1 (
            .in0(N__17932),
            .in1(N__18925),
            .in2(N__17880),
            .in3(N__18798),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_3_7_2.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_3_7_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_3_7_2.LUT_INIT=16'b1111010001000100;
    LogicCell40 i1_3_lut_4_lut_LC_3_7_2 (
            .in0(N__24446),
            .in1(N__25099),
            .in2(N__28713),
            .in3(N__30518),
            .lcout(n15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_3_7_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i2_LC_3_7_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_3_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_3_7_3  (
            .in0(_gnd_net_),
            .in1(N__24447),
            .in2(_gnd_net_),
            .in3(N__19179),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49732),
            .ce(),
            .sr(N__18270));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_625_LC_3_7_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_625_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_625_LC_3_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_625_LC_3_7_4  (
            .in0(N__21197),
            .in1(N__21295),
            .in2(N__23342),
            .in3(N__21507),
            .lcout(\c0.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_718_LC_3_7_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_718_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_718_LC_3_7_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_718_LC_3_7_5  (
            .in0(N__19000),
            .in1(N__18924),
            .in2(_gnd_net_),
            .in3(N__18590),
            .lcout(n1166),
            .ltout(n1166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_588_LC_3_7_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_588_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_588_LC_3_7_6 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \c0.i1_2_lut_adj_588_LC_3_7_6  (
            .in0(_gnd_net_),
            .in1(N__25098),
            .in2(N__18096),
            .in3(_gnd_net_),
            .lcout(\c0.n10497 ),
            .ltout(\c0.n10497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_644_LC_3_7_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_644_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_644_LC_3_7_7 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_644_LC_3_7_7  (
            .in0(N__19087),
            .in1(N__18093),
            .in2(N__18066),
            .in3(N__18041),
            .lcout(\c0.n17239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_3_8_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_3_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_3_8_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_3_8_0  (
            .in0(N__17936),
            .in1(N__20847),
            .in2(_gnd_net_),
            .in3(N__21535),
            .lcout(\c0.FRAME_MATCHER_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49722),
            .ce(),
            .sr(N__18132));
    defparam \c0.rx.i1_2_lut_adj_398_LC_3_8_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_398_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_398_LC_3_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_398_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(N__27999),
            .in2(_gnd_net_),
            .in3(N__27939),
            .lcout(\c0.rx.n57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15583_2_lut_LC_3_8_3 .C_ON=1'b0;
    defparam \c0.rx.i15583_2_lut_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15583_2_lut_LC_3_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i15583_2_lut_LC_3_8_3  (
            .in0(N__27942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26975),
            .lcout(\c0.rx.n18304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_397_LC_3_8_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_397_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_397_LC_3_8_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_397_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__27430),
            .in2(_gnd_net_),
            .in3(N__27940),
            .lcout(\c0.rx.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_421_LC_3_8_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_421_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_421_LC_3_8_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \c0.rx.i1_2_lut_adj_421_LC_3_8_5  (
            .in0(N__27941),
            .in1(_gnd_net_),
            .in2(N__27449),
            .in3(_gnd_net_),
            .lcout(\c0.rx.n167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_adj_413_LC_3_8_6 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_adj_413_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_adj_413_LC_3_8_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.rx.i1_3_lut_adj_413_LC_3_8_6  (
            .in0(N__34220),
            .in1(N__21951),
            .in2(_gnd_net_),
            .in3(N__24448),
            .lcout(\c0.rx.n12963 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_510_LC_3_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_510_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_510_LC_3_9_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.i1_2_lut_adj_510_LC_3_9_0  (
            .in0(N__33237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21291),
            .lcout(n1437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_452_LC_3_9_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_452_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_452_LC_3_9_1 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \c0.i1_3_lut_adj_452_LC_3_9_1  (
            .in0(N__20843),
            .in1(N__18161),
            .in2(_gnd_net_),
            .in3(N__21454),
            .lcout(),
            .ltout(\c0.n6_adj_2265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_455_LC_3_9_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_455_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_455_LC_3_9_2 .LUT_INIT=16'b1111111101011101;
    LogicCell40 \c0.i3_4_lut_adj_455_LC_3_9_2  (
            .in0(N__18730),
            .in1(N__18599),
            .in2(N__18135),
            .in3(N__18948),
            .lcout(\c0.n18907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_593_LC_3_9_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_593_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_593_LC_3_9_3 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_593_LC_3_9_3  (
            .in0(N__18600),
            .in1(N__18834),
            .in2(N__23336),
            .in3(N__19041),
            .lcout(),
            .ltout(n13_adj_2469_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_3_9_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_3_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i0_LC_3_9_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_3_9_4  (
            .in0(N__18731),
            .in1(N__18189),
            .in2(N__18120),
            .in3(N__18117),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_31_i3_2_lut_3_lut_4_lut_LC_3_9_5 .C_ON=1'b0;
    defparam \c0.select_284_Select_31_i3_2_lut_3_lut_4_lut_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_31_i3_2_lut_3_lut_4_lut_LC_3_9_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_31_i3_2_lut_3_lut_4_lut_LC_3_9_5  (
            .in0(N__21711),
            .in1(N__21917),
            .in2(N__20985),
            .in3(N__21455),
            .lcout(\c0.n3_adj_2279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_20_i3_2_lut_3_lut_4_lut_LC_3_9_7 .C_ON=1'b0;
    defparam \c0.select_284_Select_20_i3_2_lut_3_lut_4_lut_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_20_i3_2_lut_3_lut_4_lut_LC_3_9_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_20_i3_2_lut_3_lut_4_lut_LC_3_9_7  (
            .in0(N__21712),
            .in1(N__21918),
            .in2(N__22026),
            .in3(N__21456),
            .lcout(\c0.n3_adj_2301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_716_LC_3_10_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_716_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_716_LC_3_10_0 .LUT_INIT=16'b1100110100000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_716_LC_3_10_0  (
            .in0(N__20797),
            .in1(N__20952),
            .in2(N__18201),
            .in3(N__19001),
            .lcout(\c0.n2_adj_2315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_746_LC_3_10_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_746_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_746_LC_3_10_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_746_LC_3_10_1  (
            .in0(N__23404),
            .in1(N__23295),
            .in2(N__20975),
            .in3(N__25598),
            .lcout(n15118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_614_LC_3_10_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_614_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_614_LC_3_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_614_LC_3_10_2  (
            .in0(N__25596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23402),
            .lcout(\c0.n232 ),
            .ltout(\c0.n232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_777_LC_3_10_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_777_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_777_LC_3_10_3 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_777_LC_3_10_3  (
            .in0(N__20950),
            .in1(N__23290),
            .in2(N__18219),
            .in3(N__20795),
            .lcout(\c0.n7528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i0_LC_3_10_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i0_LC_3_10_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_3_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(N__24500),
            .in2(_gnd_net_),
            .in3(N__19215),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(N__18258));
    defparam \c0.i1_3_lut_4_lut_adj_634_LC_3_10_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_634_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_634_LC_3_10_5 .LUT_INIT=16'b1010101010111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_634_LC_3_10_5  (
            .in0(N__20951),
            .in1(N__23294),
            .in2(N__18818),
            .in3(N__20796),
            .lcout(\c0.n6_adj_2364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_3_10_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_578_LC_3_10_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_578_LC_3_10_6  (
            .in0(N__25597),
            .in1(_gnd_net_),
            .in2(N__23331),
            .in3(N__23403),
            .lcout(n237),
            .ltout(n237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_828_LC_3_10_7.C_ON=1'b0;
    defparam i1_4_lut_adj_828_LC_3_10_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_828_LC_3_10_7.LUT_INIT=16'b1010101000001000;
    LogicCell40 i1_4_lut_adj_828_LC_3_10_7 (
            .in0(N__19002),
            .in1(N__18833),
            .in2(N__18192),
            .in3(N__19040),
            .lcout(n22_adj_2465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10991_2_lut_3_lut_4_lut_LC_3_11_0 .C_ON=1'b0;
    defparam \c0.i10991_2_lut_3_lut_4_lut_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10991_2_lut_3_lut_4_lut_LC_3_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10991_2_lut_3_lut_4_lut_LC_3_11_0  (
            .in0(N__21196),
            .in1(N__21296),
            .in2(N__19577),
            .in3(N__21508),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_3_11_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i16_LC_3_11_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_3_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__19548),
            .in2(_gnd_net_),
            .in3(N__24499),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49693),
            .ce(),
            .sr(N__18183));
    defparam \c0.select_284_Select_16_i3_2_lut_3_lut_LC_3_11_2 .C_ON=1'b0;
    defparam \c0.select_284_Select_16_i3_2_lut_3_lut_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_16_i3_2_lut_3_lut_LC_3_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_284_Select_16_i3_2_lut_3_lut_LC_3_11_2  (
            .in0(N__19573),
            .in1(N__21678),
            .in2(_gnd_net_),
            .in3(N__22571),
            .lcout(\c0.n3_adj_2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_556_LC_3_11_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_556_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_556_LC_3_11_3 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_556_LC_3_11_3  (
            .in0(N__33142),
            .in1(N__18789),
            .in2(N__30043),
            .in3(N__24498),
            .lcout(\c0.n10353 ),
            .ltout(\c0.n10353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_18_i3_2_lut_3_lut_LC_3_11_4 .C_ON=1'b0;
    defparam \c0.select_284_Select_18_i3_2_lut_3_lut_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_18_i3_2_lut_3_lut_LC_3_11_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.select_284_Select_18_i3_2_lut_3_lut_LC_3_11_4  (
            .in0(N__24699),
            .in1(_gnd_net_),
            .in2(N__18285),
            .in3(N__22572),
            .lcout(\c0.n3_adj_2305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_596_LC_3_11_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_596_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_596_LC_3_11_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_596_LC_3_11_5  (
            .in0(N__21511),
            .in1(N__25659),
            .in2(N__21710),
            .in3(N__21914),
            .lcout(\c0.n3_adj_2345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_598_LC_3_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_598_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_598_LC_3_11_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_598_LC_3_11_6  (
            .in0(N__21912),
            .in1(N__21671),
            .in2(N__23335),
            .in3(N__21510),
            .lcout(\c0.n3_adj_2343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_627_LC_3_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_627_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_627_LC_3_11_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_627_LC_3_11_7  (
            .in0(N__21509),
            .in1(N__23427),
            .in2(N__21709),
            .in3(N__21913),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_23_i3_2_lut_3_lut_4_lut_LC_3_12_0 .C_ON=1'b0;
    defparam \c0.select_284_Select_23_i3_2_lut_3_lut_4_lut_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_23_i3_2_lut_3_lut_4_lut_LC_3_12_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_23_i3_2_lut_3_lut_4_lut_LC_3_12_0  (
            .in0(N__19854),
            .in1(N__21897),
            .in2(N__21699),
            .in3(N__21525),
            .lcout(\c0.n3_adj_2295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i23_LC_3_12_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i23_LC_3_12_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_3_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__24501),
            .in2(_gnd_net_),
            .in3(N__19830),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(N__18246));
    defparam \c0.i10982_2_lut_LC_3_12_2 .C_ON=1'b0;
    defparam \c0.i10982_2_lut_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10982_2_lut_LC_3_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10982_2_lut_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__19853),
            .in2(_gnd_net_),
            .in3(N__22566),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_25_i3_2_lut_3_lut_4_lut_LC_3_12_3 .C_ON=1'b0;
    defparam \c0.select_284_Select_25_i3_2_lut_3_lut_4_lut_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_25_i3_2_lut_3_lut_4_lut_LC_3_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_25_i3_2_lut_3_lut_4_lut_LC_3_12_3  (
            .in0(N__21521),
            .in1(N__21647),
            .in2(N__21919),
            .in3(N__19749),
            .lcout(\c0.n3_adj_2291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_26_i3_2_lut_3_lut_4_lut_LC_3_12_4 .C_ON=1'b0;
    defparam \c0.select_284_Select_26_i3_2_lut_3_lut_4_lut_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_26_i3_2_lut_3_lut_4_lut_LC_3_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_26_i3_2_lut_3_lut_4_lut_LC_3_12_4  (
            .in0(N__22438),
            .in1(N__21898),
            .in2(N__21700),
            .in3(N__21526),
            .lcout(\c0.n3_adj_2289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_27_i3_2_lut_3_lut_4_lut_LC_3_12_5 .C_ON=1'b0;
    defparam \c0.select_284_Select_27_i3_2_lut_3_lut_4_lut_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_27_i3_2_lut_3_lut_4_lut_LC_3_12_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.select_284_Select_27_i3_2_lut_3_lut_4_lut_LC_3_12_5  (
            .in0(N__21524),
            .in1(N__22397),
            .in2(N__21921),
            .in3(N__21649),
            .lcout(\c0.n3_adj_2287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_28_i3_2_lut_3_lut_4_lut_LC_3_12_6 .C_ON=1'b0;
    defparam \c0.select_284_Select_28_i3_2_lut_3_lut_4_lut_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_28_i3_2_lut_3_lut_4_lut_LC_3_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_28_i3_2_lut_3_lut_4_lut_LC_3_12_6  (
            .in0(N__21646),
            .in1(N__21887),
            .in2(N__22287),
            .in3(N__21522),
            .lcout(\c0.n3_adj_2285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_6_i3_2_lut_3_lut_4_lut_LC_3_12_7 .C_ON=1'b0;
    defparam \c0.select_284_Select_6_i3_2_lut_3_lut_4_lut_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_6_i3_2_lut_3_lut_4_lut_LC_3_12_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.select_284_Select_6_i3_2_lut_3_lut_4_lut_LC_3_12_7  (
            .in0(N__21523),
            .in1(N__22178),
            .in2(N__21920),
            .in3(N__21648),
            .lcout(\c0.n3_adj_2334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i26_LC_3_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i26_LC_3_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_3_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__24566),
            .in2(_gnd_net_),
            .in3(N__19689),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49682),
            .ce(),
            .sr(N__18321));
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__24568),
            .in2(_gnd_net_),
            .in3(N__19674),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49677),
            .ce(),
            .sr(N__18315));
    defparam \c0.FRAME_MATCHER_i_i8_LC_3_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i8_LC_3_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_3_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__24621),
            .in2(_gnd_net_),
            .in3(N__19278),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(N__18852));
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__24622),
            .in2(_gnd_net_),
            .in3(N__20253),
            .lcout(FRAME_MATCHER_i_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49670),
            .ce(),
            .sr(N__18309));
    defparam \c0.FRAME_MATCHER_i_i19_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i19_LC_3_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_3_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__24624),
            .in2(_gnd_net_),
            .in3(N__19467),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(N__18297));
    defparam \c0.select_284_Select_19_i3_2_lut_3_lut_4_lut_LC_3_18_3 .C_ON=1'b0;
    defparam \c0.select_284_Select_19_i3_2_lut_3_lut_4_lut_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_19_i3_2_lut_3_lut_4_lut_LC_3_18_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.select_284_Select_19_i3_2_lut_3_lut_4_lut_LC_3_18_3  (
            .in0(N__21698),
            .in1(N__21911),
            .in2(N__21036),
            .in3(N__21542),
            .lcout(\c0.n3_adj_2303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.PHASES_i2_LC_3_29_7 .C_ON=1'b0;
    defparam \control.PHASES_i2_LC_3_29_7 .SEQ_MODE=4'b1000;
    defparam \control.PHASES_i2_LC_3_29_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \control.PHASES_i2_LC_3_29_7  (
            .in0(N__35639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35411),
            .lcout(PIN_2_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49758),
            .ce(N__20163),
            .sr(N__35352));
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_1_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(N__18544),
            .in2(_gnd_net_),
            .in3(N__20497),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49823),
            .ce(),
            .sr(N__18522));
    defparam \c0.FRAME_MATCHER_state_i21_LC_4_2_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_4_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_4_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_4_2_0  (
            .in0(_gnd_net_),
            .in1(N__18464),
            .in2(_gnd_net_),
            .in3(N__20089),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49811),
            .ce(),
            .sr(N__18447));
    defparam \c0.i17_4_lut_LC_4_3_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_4_3_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_LC_4_3_0  (
            .in0(N__18502),
            .in1(N__18652),
            .in2(N__18465),
            .in3(N__18484),
            .lcout(\c0.n46_adj_2356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i18_LC_4_3_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_4_3_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_4_3_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_4_3_1  (
            .in0(N__18486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20092),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49800),
            .ce(),
            .sr(N__18474));
    defparam \c0.i1_2_lut_adj_473_LC_4_3_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_473_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_473_LC_4_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_473_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__18485),
            .in2(_gnd_net_),
            .in3(N__18703),
            .lcout(\c0.n17293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_480_LC_4_3_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_480_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_480_LC_4_3_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i1_2_lut_adj_480_LC_4_3_3  (
            .in0(N__18702),
            .in1(N__18463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n8_adj_2247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_475_LC_4_3_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_475_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_475_LC_4_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_475_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__20136),
            .in2(_gnd_net_),
            .in3(N__18701),
            .lcout(\c0.n8_adj_2250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_491_LC_4_3_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_491_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_491_LC_4_3_5 .LUT_INIT=16'b1111110111001100;
    LogicCell40 \c0.i1_4_lut_adj_491_LC_4_3_5  (
            .in0(N__18421),
            .in1(N__18887),
            .in2(N__18336),
            .in3(N__19119),
            .lcout(\c0.n8_adj_2273 ),
            .ltout(\c0.n8_adj_2273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_477_LC_4_3_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_477_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_477_LC_4_3_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_477_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18708),
            .in3(N__20423),
            .lcout(\c0.n8_adj_2249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_488_LC_4_3_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_488_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_488_LC_4_3_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_488_LC_4_3_7  (
            .in0(N__18704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18684),
            .lcout(\c0.n17273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_4_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__18654),
            .in2(_gnd_net_),
            .in3(N__20491),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49788),
            .ce(),
            .sr(N__18636));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_791_LC_4_5_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_791_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_791_LC_4_5_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_791_LC_4_5_0  (
            .in0(N__33180),
            .in1(N__33263),
            .in2(N__30044),
            .in3(N__30108),
            .lcout(\c0.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_4_5_1 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_4_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i28_4_lut_LC_4_5_1  (
            .in0(N__18630),
            .in1(N__20286),
            .in2(N__18621),
            .in3(N__18609),
            .lcout(\c0.n10513 ),
            .ltout(\c0.n10513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_804_LC_4_5_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_804_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_804_LC_4_5_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_804_LC_4_5_2  (
            .in0(N__33179),
            .in1(N__30034),
            .in2(N__18603),
            .in3(N__33264),
            .lcout(FRAME_MATCHER_i_31__N_1275),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_547_LC_4_5_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_547_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_547_LC_4_5_3 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_547_LC_4_5_3  (
            .in0(N__30110),
            .in1(N__30022),
            .in2(N__33282),
            .in3(N__33182),
            .lcout(\c0.n6033 ),
            .ltout(\c0.n6033_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i7_LC_4_5_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i7_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i7_LC_4_5_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.data_out_frame2_0___i7_LC_4_5_4  (
            .in0(N__28814),
            .in1(N__28935),
            .in2(N__18561),
            .in3(N__28836),
            .lcout(\c0.data_out_frame2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49772),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_799_LC_4_5_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_799_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_799_LC_4_5_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_799_LC_4_5_5  (
            .in0(N__30109),
            .in1(N__30021),
            .in2(N__33281),
            .in3(N__33181),
            .lcout(FRAME_MATCHER_i_31__N_1272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1014_2_lut_LC_4_5_6 .C_ON=1'b0;
    defparam \c0.i1014_2_lut_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1014_2_lut_LC_4_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1014_2_lut_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__23132),
            .in2(_gnd_net_),
            .in3(N__25914),
            .lcout(\c0.n2126 ),
            .ltout(\c0.n2126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_509_LC_4_5_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_509_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_509_LC_4_5_7 .LUT_INIT=16'b1111111101111011;
    LogicCell40 \c0.i11_4_lut_adj_509_LC_4_5_7  (
            .in0(N__23679),
            .in1(N__22931),
            .in2(N__18753),
            .in3(N__20277),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_4_6_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_4_6_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_4_6_0  (
            .in0(N__30112),
            .in1(N__33170),
            .in2(N__33277),
            .in3(N__30007),
            .lcout(FRAME_MATCHER_i_31__N_1273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_616_LC_4_6_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_616_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_616_LC_4_6_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_616_LC_4_6_1  (
            .in0(N__33169),
            .in1(N__33255),
            .in2(N__30035),
            .in3(N__30111),
            .lcout(FRAME_MATCHER_i_31__N_1270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_469_LC_4_6_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_469_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_469_LC_4_6_2 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i7_4_lut_adj_469_LC_4_6_2  (
            .in0(N__26008),
            .in1(N__23083),
            .in2(N__23520),
            .in3(N__26043),
            .lcout(),
            .ltout(\c0.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_4_6_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_4_6_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i14_4_lut_LC_4_6_3  (
            .in0(N__18750),
            .in1(N__26307),
            .in2(N__18744),
            .in3(N__25952),
            .lcout(),
            .ltout(\c0.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_4_6_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_4_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_LC_4_6_4  (
            .in0(N__26262),
            .in1(N__18714),
            .in2(N__18741),
            .in3(N__18774),
            .lcout(\c0.n50 ),
            .ltout(\c0.n50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11086_2_lut_LC_4_6_5 .C_ON=1'b0;
    defparam \c0.i11086_2_lut_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11086_2_lut_LC_4_6_5 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \c0.i11086_2_lut_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__25058),
            .in2(N__18738),
            .in3(_gnd_net_),
            .lcout(n13849),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_519_LC_4_6_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_519_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_519_LC_4_6_6 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i3_4_lut_adj_519_LC_4_6_6  (
            .in0(N__20574),
            .in1(N__25443),
            .in2(N__22652),
            .in3(N__20607),
            .lcout(\c0.n19_adj_2351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_714_LC_4_6_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_714_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_714_LC_4_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_714_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(N__33259),
            .in2(_gnd_net_),
            .in3(N__30113),
            .lcout(\c0.n10346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_7_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_4_7_0  (
            .in0(N__22747),
            .in1(N__30724),
            .in2(_gnd_net_),
            .in3(N__30306),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_4_7_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_4_7_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_4_7_1  (
            .in0(N__26002),
            .in1(N__23591),
            .in2(_gnd_net_),
            .in3(N__24155),
            .lcout(data_in_frame_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_4_7_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_4_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i47_LC_4_7_2  (
            .in0(N__27621),
            .in1(N__20546),
            .in2(_gnd_net_),
            .in3(N__23635),
            .lcout(data_in_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_514_LC_4_7_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_514_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_514_LC_4_7_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i1_4_lut_adj_514_LC_4_7_3  (
            .in0(N__26133),
            .in1(N__23107),
            .in2(N__20592),
            .in3(N__23082),
            .lcout(),
            .ltout(\c0.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_521_LC_4_7_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_521_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_521_LC_4_7_4 .LUT_INIT=16'b1111011011111111;
    LogicCell40 \c0.i9_4_lut_adj_521_LC_4_7_4  (
            .in0(N__23556),
            .in1(N__23180),
            .in2(N__18777),
            .in3(N__22989),
            .lcout(\c0.n25_adj_2352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15103_3_lut_4_lut_LC_4_7_5 .C_ON=1'b0;
    defparam \c0.i15103_3_lut_4_lut_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15103_3_lut_4_lut_LC_4_7_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \c0.i15103_3_lut_4_lut_LC_4_7_5  (
            .in0(N__20590),
            .in1(N__25998),
            .in2(N__20573),
            .in3(N__25913),
            .lcout(),
            .ltout(\c0.n17962_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_695_LC_4_7_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_695_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_695_LC_4_7_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i10_4_lut_adj_695_LC_4_7_6  (
            .in0(N__26394),
            .in1(N__23181),
            .in2(N__18768),
            .in3(N__26079),
            .lcout(\c0.n24_adj_2418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i1_LC_4_8_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i1_LC_4_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i1_LC_4_8_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i1_LC_4_8_0  (
            .in0(N__25011),
            .in1(N__48286),
            .in2(N__30663),
            .in3(N__30519),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49733),
            .ce(),
            .sr(N__18765));
    defparam \c0.tx2.i15302_3_lut_LC_4_8_1 .C_ON=1'b0;
    defparam \c0.tx2.i15302_3_lut_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15302_3_lut_LC_4_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.i15302_3_lut_LC_4_8_1  (
            .in0(N__33941),
            .in1(N__28512),
            .in2(_gnd_net_),
            .in3(N__48840),
            .lcout(\c0.tx2.n18163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15303_3_lut_LC_4_8_2 .C_ON=1'b0;
    defparam \c0.tx2.i15303_3_lut_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15303_3_lut_LC_4_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx2.i15303_3_lut_LC_4_8_2  (
            .in0(N__28548),
            .in1(N__33942),
            .in2(_gnd_net_),
            .in3(N__42993),
            .lcout(\c0.tx2.n18164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_LC_4_8_3 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_LC_4_8_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.tx2.i2_3_lut_LC_4_8_3  (
            .in0(N__29094),
            .in1(N__29070),
            .in2(_gnd_net_),
            .in3(N__29043),
            .lcout(\c0.tx2.n12769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10981_2_lut_LC_4_8_4 .C_ON=1'b0;
    defparam \c0.i10981_2_lut_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10981_2_lut_LC_4_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10981_2_lut_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__19809),
            .in2(_gnd_net_),
            .in3(N__22501),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10983_2_lut_LC_4_8_5 .C_ON=1'b0;
    defparam \c0.i10983_2_lut_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10983_2_lut_LC_4_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10983_2_lut_LC_4_8_5  (
            .in0(N__22502),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19920),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10984_2_lut_LC_4_8_6 .C_ON=1'b0;
    defparam \c0.i10984_2_lut_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10984_2_lut_LC_4_8_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10984_2_lut_LC_4_8_6  (
            .in0(N__19425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22503),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10992_2_lut_LC_4_8_7 .C_ON=1'b0;
    defparam \c0.i10992_2_lut_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10992_2_lut_LC_4_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10992_2_lut_LC_4_8_7  (
            .in0(N__22504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19638),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_576_LC_4_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_576_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_576_LC_4_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_576_LC_4_9_0  (
            .in0(N__21163),
            .in1(N__21254),
            .in2(_gnd_net_),
            .in3(N__21373),
            .lcout(\c0.n9575 ),
            .ltout(\c0.n9575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_575_LC_4_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_575_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_575_LC_4_9_1 .LUT_INIT=16'b0000000011001111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_575_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__29982),
            .in2(N__18837),
            .in3(N__20816),
            .lcout(n12999),
            .ltout(n12999_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_591_LC_4_9_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_591_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_591_LC_4_9_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_591_LC_4_9_2  (
            .in0(N__18822),
            .in1(N__23356),
            .in2(N__18801),
            .in3(N__19039),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_571_LC_4_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_571_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_571_LC_4_9_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_571_LC_4_9_3  (
            .in0(N__20976),
            .in1(N__29983),
            .in2(_gnd_net_),
            .in3(N__19066),
            .lcout(n12966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10989_2_lut_3_lut_4_lut_LC_4_9_4 .C_ON=1'b0;
    defparam \c0.i10989_2_lut_3_lut_4_lut_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10989_2_lut_3_lut_4_lut_LC_4_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10989_2_lut_3_lut_4_lut_LC_4_9_4  (
            .in0(N__21164),
            .in1(N__21255),
            .in2(N__19524),
            .in3(N__21374),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_449_LC_4_9_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_449_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_449_LC_4_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i3_4_lut_adj_449_LC_4_9_5  (
            .in0(N__21375),
            .in1(N__18941),
            .in2(N__18906),
            .in3(N__20836),
            .lcout(),
            .ltout(\c0.n16685_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_453_LC_4_9_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_453_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_453_LC_4_9_6 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \c0.i2_4_lut_adj_453_LC_4_9_6  (
            .in0(N__19016),
            .in1(N__19004),
            .in2(N__18951),
            .in3(N__20775),
            .lcout(\c0.n6_adj_2267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i57_3_lut_4_lut_LC_4_9_7 .C_ON=1'b0;
    defparam \c0.i57_3_lut_4_lut_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i57_3_lut_4_lut_LC_4_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i57_3_lut_4_lut_LC_4_9_7  (
            .in0(N__21372),
            .in1(N__18940),
            .in2(N__18905),
            .in3(N__21788),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_7_i3_2_lut_3_lut_4_lut_LC_4_10_0 .C_ON=1'b0;
    defparam \c0.select_284_Select_7_i3_2_lut_3_lut_4_lut_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_7_i3_2_lut_3_lut_4_lut_LC_4_10_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_7_i3_2_lut_3_lut_4_lut_LC_4_10_0  (
            .in0(N__19367),
            .in1(N__21811),
            .in2(N__21697),
            .in3(N__21423),
            .lcout(\c0.n3_adj_2332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_4_10_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i7_LC_4_10_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_4_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__24533),
            .in2(_gnd_net_),
            .in3(N__19341),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(N__18864));
    defparam \c0.i11000_2_lut_LC_4_10_2 .C_ON=1'b0;
    defparam \c0.i11000_2_lut_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11000_2_lut_LC_4_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i11000_2_lut_LC_4_10_2  (
            .in0(N__22500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19366),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_8_i3_2_lut_3_lut_4_lut_LC_4_10_3 .C_ON=1'b0;
    defparam \c0.select_284_Select_8_i3_2_lut_3_lut_4_lut_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_8_i3_2_lut_3_lut_4_lut_LC_4_10_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_8_i3_2_lut_3_lut_4_lut_LC_4_10_3  (
            .in0(N__21421),
            .in1(N__21639),
            .in2(N__21870),
            .in3(N__19322),
            .lcout(\c0.n3_adj_2330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_9_i3_2_lut_3_lut_4_lut_LC_4_10_4 .C_ON=1'b0;
    defparam \c0.select_284_Select_9_i3_2_lut_3_lut_4_lut_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_9_i3_2_lut_3_lut_4_lut_LC_4_10_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_9_i3_2_lut_3_lut_4_lut_LC_4_10_4  (
            .in0(N__20234),
            .in1(N__21810),
            .in2(N__21696),
            .in3(N__21422),
            .lcout(\c0.n3_adj_2328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10998_2_lut_LC_4_10_5 .C_ON=1'b0;
    defparam \c0.i10998_2_lut_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10998_2_lut_LC_4_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10998_2_lut_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(N__20233),
            .in2(_gnd_net_),
            .in3(N__22498),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10999_2_lut_LC_4_10_6 .C_ON=1'b0;
    defparam \c0.i10999_2_lut_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10999_2_lut_LC_4_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10999_2_lut_LC_4_10_6  (
            .in0(N__22499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19323),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10980_2_lut_LC_4_10_7 .C_ON=1'b0;
    defparam \c0.i10980_2_lut_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10980_2_lut_LC_4_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10980_2_lut_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(N__19747),
            .in2(_gnd_net_),
            .in3(N__22497),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_2_lut_LC_4_11_0 .C_ON=1'b1;
    defparam \c0.add_977_2_lut_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_2_lut_LC_4_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_2_lut_LC_4_11_0  (
            .in0(N__22116),
            .in1(N__23401),
            .in2(N__23853),
            .in3(N__19209),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_0 ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\c0.n16486 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_3_lut_LC_4_11_1 .C_ON=1'b1;
    defparam \c0.add_977_3_lut_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_3_lut_LC_4_11_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_3_lut_LC_4_11_1  (
            .in0(N__21117),
            .in1(N__25647),
            .in2(N__23856),
            .in3(N__19194),
            .lcout(\c0.n27_adj_2426 ),
            .ltout(),
            .carryin(\c0.n16486 ),
            .carryout(\c0.n16487 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_4_lut_LC_4_11_2 .C_ON=1'b1;
    defparam \c0.add_977_4_lut_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_4_lut_LC_4_11_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_4_lut_LC_4_11_2  (
            .in0(N__19191),
            .in1(N__23790),
            .in2(N__23366),
            .in3(N__19167),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(\c0.n16487 ),
            .carryout(\c0.n16488 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_5_lut_LC_4_11_3 .C_ON=1'b1;
    defparam \c0.add_977_5_lut_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_5_lut_LC_4_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_5_lut_LC_4_11_3  (
            .in0(N__20859),
            .in1(N__22344),
            .in2(N__23857),
            .in3(N__19164),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_3 ),
            .ltout(),
            .carryin(\c0.n16488 ),
            .carryout(\c0.n16489 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_6_lut_LC_4_11_4 .C_ON=1'b1;
    defparam \c0.add_977_6_lut_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_6_lut_LC_4_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_6_lut_LC_4_11_4  (
            .in0(N__21930),
            .in1(N__21746),
            .in2(N__23854),
            .in3(N__19152),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_4 ),
            .ltout(),
            .carryin(\c0.n16489 ),
            .carryout(\c0.n16490 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_7_lut_LC_4_11_5 .C_ON=1'b1;
    defparam \c0.add_977_7_lut_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_7_lut_LC_4_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_7_lut_LC_4_11_5  (
            .in0(N__20868),
            .in1(N__21971),
            .in2(N__23858),
            .in3(N__19149),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_5 ),
            .ltout(),
            .carryin(\c0.n16490 ),
            .carryout(\c0.n16491 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_8_lut_LC_4_11_6 .C_ON=1'b1;
    defparam \c0.add_977_8_lut_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_8_lut_LC_4_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_8_lut_LC_4_11_6  (
            .in0(N__22128),
            .in1(N__22158),
            .in2(N__23855),
            .in3(N__19380),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_6 ),
            .ltout(),
            .carryin(\c0.n16491 ),
            .carryout(\c0.n16492 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_9_lut_LC_4_11_7 .C_ON=1'b1;
    defparam \c0.add_977_9_lut_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_9_lut_LC_4_11_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_9_lut_LC_4_11_7  (
            .in0(N__19377),
            .in1(N__19365),
            .in2(N__23859),
            .in3(N__19335),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_7 ),
            .ltout(),
            .carryin(\c0.n16492 ),
            .carryout(\c0.n16493 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_10_lut_LC_4_12_0 .C_ON=1'b1;
    defparam \c0.add_977_10_lut_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_10_lut_LC_4_12_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_10_lut_LC_4_12_0  (
            .in0(N__19332),
            .in1(N__19318),
            .in2(N__23906),
            .in3(N__19266),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_8 ),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\c0.n16494 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_11_lut_LC_4_12_1 .C_ON=1'b1;
    defparam \c0.add_977_11_lut_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_11_lut_LC_4_12_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_11_lut_LC_4_12_1  (
            .in0(N__19263),
            .in1(N__23863),
            .in2(N__20235),
            .in3(N__19254),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_9 ),
            .ltout(),
            .carryin(\c0.n16494 ),
            .carryout(\c0.n16495 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_12_lut_LC_4_12_2 .C_ON=1'b1;
    defparam \c0.add_977_12_lut_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_12_lut_LC_4_12_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_12_lut_LC_4_12_2  (
            .in0(N__22188),
            .in1(N__22223),
            .in2(N__23907),
            .in3(N__19239),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_10 ),
            .ltout(),
            .carryin(\c0.n16495 ),
            .carryout(\c0.n16496 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_13_lut_LC_4_12_3 .C_ON=1'b1;
    defparam \c0.add_977_13_lut_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_13_lut_LC_4_12_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_13_lut_LC_4_12_3  (
            .in0(N__22038),
            .in1(N__23867),
            .in2(N__22070),
            .in3(N__19236),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_11 ),
            .ltout(),
            .carryin(\c0.n16496 ),
            .carryout(\c0.n16497 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_14_lut_LC_4_12_4 .C_ON=1'b1;
    defparam \c0.add_977_14_lut_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_14_lut_LC_4_12_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_14_lut_LC_4_12_4  (
            .in0(N__22584),
            .in1(N__22618),
            .in2(N__23908),
            .in3(N__19221),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_12 ),
            .ltout(),
            .carryin(\c0.n16497 ),
            .carryout(\c0.n16498 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_15_lut_LC_4_12_5 .C_ON=1'b1;
    defparam \c0.add_977_15_lut_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_15_lut_LC_4_12_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_15_lut_LC_4_12_5  (
            .in0(N__22233),
            .in1(N__23871),
            .in2(N__24381),
            .in3(N__19218),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_13 ),
            .ltout(),
            .carryin(\c0.n16498 ),
            .carryout(\c0.n16499 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_16_lut_LC_4_12_6 .C_ON=1'b1;
    defparam \c0.add_977_16_lut_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_16_lut_LC_4_12_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_16_lut_LC_4_12_6  (
            .in0(N__21069),
            .in1(N__21103),
            .in2(N__23909),
            .in3(N__19653),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_14 ),
            .ltout(),
            .carryin(\c0.n16499 ),
            .carryout(\c0.n16500 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_17_lut_LC_4_12_7 .C_ON=1'b1;
    defparam \c0.add_977_17_lut_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_17_lut_LC_4_12_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_17_lut_LC_4_12_7  (
            .in0(N__19650),
            .in1(N__23875),
            .in2(N__19637),
            .in3(N__19593),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_15 ),
            .ltout(),
            .carryin(\c0.n16500 ),
            .carryout(\c0.n16501 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_18_lut_LC_4_13_0 .C_ON=1'b1;
    defparam \c0.add_977_18_lut_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_18_lut_LC_4_13_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_18_lut_LC_4_13_0  (
            .in0(N__19590),
            .in1(N__23877),
            .in2(N__19581),
            .in3(N__19539),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_16 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\c0.n16502 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_19_lut_LC_4_13_1 .C_ON=1'b1;
    defparam \c0.add_977_19_lut_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_19_lut_LC_4_13_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_19_lut_LC_4_13_1  (
            .in0(N__19536),
            .in1(N__23881),
            .in2(N__19520),
            .in3(N__19473),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_17 ),
            .ltout(),
            .carryin(\c0.n16502 ),
            .carryout(\c0.n16503 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_20_lut_LC_4_13_2 .C_ON=1'b1;
    defparam \c0.add_977_20_lut_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_20_lut_LC_4_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_20_lut_LC_4_13_2  (
            .in0(N__20880),
            .in1(N__24703),
            .in2(N__23911),
            .in3(N__19470),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_18 ),
            .ltout(),
            .carryin(\c0.n16503 ),
            .carryout(\c0.n16504 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_21_lut_LC_4_13_3 .C_ON=1'b1;
    defparam \c0.add_977_21_lut_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_21_lut_LC_4_13_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_21_lut_LC_4_13_3  (
            .in0(N__20997),
            .in1(N__23885),
            .in2(N__21048),
            .in3(N__19455),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_19 ),
            .ltout(),
            .carryin(\c0.n16504 ),
            .carryout(\c0.n16505 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_22_lut_LC_4_13_4 .C_ON=1'b1;
    defparam \c0.add_977_22_lut_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_22_lut_LC_4_13_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_22_lut_LC_4_13_4  (
            .in0(N__21999),
            .in1(N__23876),
            .in2(N__22032),
            .in3(N__19440),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_20 ),
            .ltout(),
            .carryin(\c0.n16505 ),
            .carryout(\c0.n16506 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_23_lut_LC_4_13_5 .C_ON=1'b1;
    defparam \c0.add_977_23_lut_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_23_lut_LC_4_13_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_23_lut_LC_4_13_5  (
            .in0(N__19437),
            .in1(N__23886),
            .in2(N__19421),
            .in3(N__19383),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_21 ),
            .ltout(),
            .carryin(\c0.n16506 ),
            .carryout(\c0.n16507 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_24_lut_LC_4_13_6 .C_ON=1'b1;
    defparam \c0.add_977_24_lut_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_24_lut_LC_4_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_24_lut_LC_4_13_6  (
            .in0(N__19932),
            .in1(N__19915),
            .in2(N__23912),
            .in3(N__19866),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_22 ),
            .ltout(),
            .carryin(\c0.n16507 ),
            .carryout(\c0.n16508 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_25_lut_LC_4_13_7 .C_ON=1'b1;
    defparam \c0.add_977_25_lut_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_25_lut_LC_4_13_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_25_lut_LC_4_13_7  (
            .in0(N__19863),
            .in1(N__19852),
            .in2(N__23910),
            .in3(N__19824),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_23 ),
            .ltout(),
            .carryin(\c0.n16508 ),
            .carryout(\c0.n16509 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_26_lut_LC_4_14_0 .C_ON=1'b1;
    defparam \c0.add_977_26_lut_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_26_lut_LC_4_14_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_26_lut_LC_4_14_0  (
            .in0(N__19821),
            .in1(N__19804),
            .in2(N__23913),
            .in3(N__19761),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_24 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\c0.n16510 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_27_lut_LC_4_14_1 .C_ON=1'b1;
    defparam \c0.add_977_27_lut_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_27_lut_LC_4_14_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_27_lut_LC_4_14_1  (
            .in0(N__19758),
            .in1(N__23893),
            .in2(N__19748),
            .in3(N__19692),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_25 ),
            .ltout(),
            .carryin(\c0.n16510 ),
            .carryout(\c0.n16511 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_28_lut_LC_4_14_2 .C_ON=1'b1;
    defparam \c0.add_977_28_lut_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_28_lut_LC_4_14_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_28_lut_LC_4_14_2  (
            .in0(N__22410),
            .in1(N__22434),
            .in2(N__23914),
            .in3(N__19683),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_26 ),
            .ltout(),
            .carryin(\c0.n16511 ),
            .carryout(\c0.n16512 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_29_lut_LC_4_14_3 .C_ON=1'b1;
    defparam \c0.add_977_29_lut_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_29_lut_LC_4_14_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_29_lut_LC_4_14_3  (
            .in0(N__22578),
            .in1(N__23897),
            .in2(N__22398),
            .in3(N__19680),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_27 ),
            .ltout(),
            .carryin(\c0.n16512 ),
            .carryout(\c0.n16513 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_30_lut_LC_4_14_4 .C_ON=1'b1;
    defparam \c0.add_977_30_lut_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_30_lut_LC_4_14_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_30_lut_LC_4_14_4  (
            .in0(N__21060),
            .in1(N__23901),
            .in2(N__22283),
            .in3(N__19677),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_28 ),
            .ltout(),
            .carryin(\c0.n16513 ),
            .carryout(\c0.n16514 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_31_lut_LC_4_14_5 .C_ON=1'b1;
    defparam \c0.add_977_31_lut_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_31_lut_LC_4_14_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_31_lut_LC_4_14_5  (
            .in0(N__20682),
            .in1(N__20716),
            .in2(N__23916),
            .in3(N__19668),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_29 ),
            .ltout(),
            .carryin(\c0.n16514 ),
            .carryout(\c0.n16515 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_32_lut_LC_4_14_6 .C_ON=1'b1;
    defparam \c0.add_977_32_lut_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_32_lut_LC_4_14_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_32_lut_LC_4_14_6  (
            .in0(N__20733),
            .in1(N__20766),
            .in2(N__23915),
            .in3(N__20259),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_30 ),
            .ltout(),
            .carryin(\c0.n16515 ),
            .carryout(\c0.n16516 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_33_lut_LC_4_14_7 .C_ON=1'b0;
    defparam \c0.add_977_33_lut_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_33_lut_LC_4_14_7 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \c0.add_977_33_lut_LC_4_14_7  (
            .in0(N__23905),
            .in1(N__20949),
            .in2(N__20898),
            .in3(N__20256),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_4_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i9_LC_4_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_4_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_4_15_0  (
            .in0(N__24632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20244),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49678),
            .ce(),
            .sr(N__20199));
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_4_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_4_16_0  (
            .in0(N__24643),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20184),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(N__20175));
    defparam \control.i3_4_lut_4_lut_LC_4_29_0 .C_ON=1'b0;
    defparam \control.i3_4_lut_4_lut_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \control.i3_4_lut_4_lut_LC_4_29_0 .LUT_INIT=16'b1111111101111110;
    LogicCell40 \control.i3_4_lut_4_lut_LC_4_29_0  (
            .in0(N__35675),
            .in1(N__35546),
            .in2(N__35454),
            .in3(N__35351),
            .lcout(\control.n18909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i16_LC_5_1_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_5_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_5_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(N__20341),
            .in2(_gnd_net_),
            .in3(N__20103),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49833),
            .ce(),
            .sr(N__20151));
    defparam \c0.FRAME_MATCHER_state_i19_LC_5_2_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_5_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_5_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__20125),
            .in2(_gnd_net_),
            .in3(N__20090),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(),
            .sr(N__20109));
    defparam \c0.FRAME_MATCHER_state_i20_LC_5_3_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_5_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_5_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__20424),
            .in2(_gnd_net_),
            .in3(N__20088),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49812),
            .ce(),
            .sr(N__20508));
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_4_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_5_4_0  (
            .in0(N__20396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20499),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(),
            .sr(N__20436));
    defparam \c0.i1_2_lut_adj_525_LC_5_4_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_525_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_525_LC_5_4_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_525_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__20422),
            .in2(_gnd_net_),
            .in3(N__20395),
            .lcout(),
            .ltout(\c0.n30_adj_2355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_5_4_2 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_5_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i22_4_lut_LC_5_4_2  (
            .in0(N__20378),
            .in1(N__20342),
            .in2(N__20322),
            .in3(N__20319),
            .lcout(\c0.n51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_554_LC_5_4_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_554_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_554_LC_5_4_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_554_LC_5_4_3  (
            .in0(N__20664),
            .in1(N__25335),
            .in2(N__22932),
            .in3(N__23022),
            .lcout(\c0.n16863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_447_LC_5_4_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_447_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_447_LC_5_4_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_447_LC_5_4_4  (
            .in0(N__23021),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20663),
            .lcout(),
            .ltout(\c0.n10613_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_701_LC_5_4_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_701_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_701_LC_5_4_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i7_4_lut_adj_701_LC_5_4_5  (
            .in0(N__25392),
            .in1(N__22869),
            .in2(N__20280),
            .in3(N__25435),
            .lcout(\c0.n21_adj_2421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_5_4_6 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_5_4_6 .LUT_INIT=16'b1011011101111011;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_5_4_6  (
            .in0(N__23020),
            .in1(N__25479),
            .in2(N__22691),
            .in3(N__20662),
            .lcout(\c0.n22_adj_2346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1010_2_lut_LC_5_4_7 .C_ON=1'b0;
    defparam \c0.i1010_2_lut_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1010_2_lut_LC_5_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1010_2_lut_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__23163),
            .in2(_gnd_net_),
            .in3(N__26175),
            .lcout(\c0.n2122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_5_5_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_5_5_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_in_frame_0__i25_LC_5_5_0  (
            .in0(N__25671),
            .in1(N__20531),
            .in2(N__26642),
            .in3(N__25548),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_655_LC_5_5_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_655_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_655_LC_5_5_1 .LUT_INIT=16'b1001011011111111;
    LogicCell40 \c0.i3_4_lut_adj_655_LC_5_5_1  (
            .in0(N__22981),
            .in1(N__25953),
            .in2(N__20550),
            .in3(N__22938),
            .lcout(\c0.n19_adj_2400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_5_5_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_5_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i49_LC_5_5_2  (
            .in0(N__26633),
            .in1(N__22950),
            .in2(_gnd_net_),
            .in3(N__25864),
            .lcout(data_in_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_5_5_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_5_5_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_5_5_3  (
            .in0(N__25549),
            .in1(N__25673),
            .in2(N__20625),
            .in3(N__27096),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_5_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_5_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_5_5_4  (
            .in0(N__28011),
            .in1(N__27372),
            .in2(N__26474),
            .in3(N__26823),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_5_5_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_5_5_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i16_LC_5_5_5  (
            .in0(N__25547),
            .in1(N__25672),
            .in2(N__24180),
            .in3(N__23519),
            .lcout(\c0.data_in_frame_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_5_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_5_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_5_5_6  (
            .in0(N__28010),
            .in1(N__27371),
            .in2(N__27110),
            .in3(N__25802),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_692_LC_5_5_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_692_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_692_LC_5_5_7 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i4_4_lut_adj_692_LC_5_5_7  (
            .in0(N__20519),
            .in1(N__22851),
            .in2(N__20532),
            .in3(N__23084),
            .lcout(\c0.n18_adj_2417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_5_6_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_5_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i46_LC_5_6_0  (
            .in0(N__27217),
            .in1(N__26321),
            .in2(_gnd_net_),
            .in3(N__23637),
            .lcout(data_in_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_653_LC_5_6_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_653_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_653_LC_5_6_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i2_4_lut_adj_653_LC_5_6_1  (
            .in0(N__20520),
            .in1(N__23051),
            .in2(N__25377),
            .in3(N__26132),
            .lcout(\c0.n18_adj_2398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_5_6_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_5_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i1_LC_5_6_2  (
            .in0(N__26638),
            .in1(N__23012),
            .in2(_gnd_net_),
            .in3(N__23587),
            .lcout(data_in_frame_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_5_6_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_5_6_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \c0.data_in_frame_0__i6_LC_5_6_3  (
            .in0(N__23588),
            .in1(N__27218),
            .in2(N__23139),
            .in3(_gnd_net_),
            .lcout(data_in_frame_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_691_LC_5_6_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_691_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_691_LC_5_6_4 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i1_4_lut_adj_691_LC_5_6_4  (
            .in0(N__22707),
            .in1(N__23555),
            .in2(N__20624),
            .in3(N__20606),
            .lcout(\c0.n15_adj_2416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_748_LC_5_6_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_748_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_748_LC_5_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_748_LC_5_6_5  (
            .in0(N__25994),
            .in1(N__25902),
            .in2(_gnd_net_),
            .in3(N__23040),
            .lcout(\c0.n2137_adj_2237 ),
            .ltout(\c0.n2137_adj_2237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1026_2_lut_LC_5_6_6 .C_ON=1'b0;
    defparam \c0.i1026_2_lut_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1026_2_lut_LC_5_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1026_2_lut_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20595),
            .in3(N__23011),
            .lcout(\c0.n2138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_5_6_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_5_6_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_5_6_7  (
            .in0(N__31910),
            .in1(N__46065),
            .in2(_gnd_net_),
            .in3(N__44057),
            .lcout(\c0.n5_adj_2197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_5_7_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_5_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i17_LC_5_7_0  (
            .in0(N__26624),
            .in1(N__20591),
            .in2(_gnd_net_),
            .in3(N__26421),
            .lcout(data_in_frame_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_5_7_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_5_7_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i22_LC_5_7_1  (
            .in0(N__26422),
            .in1(_gnd_net_),
            .in2(N__27205),
            .in3(N__20572),
            .lcout(data_in_frame_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_5_7_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_5_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i23_LC_5_7_2  (
            .in0(N__27620),
            .in1(N__23109),
            .in2(_gnd_net_),
            .in3(N__26423),
            .lcout(data_in_frame_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_adj_405_LC_5_7_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_adj_405_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_adj_405_LC_5_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_adj_405_LC_5_7_3  (
            .in0(N__23221),
            .in1(N__25670),
            .in2(N__23349),
            .in3(N__23462),
            .lcout(n16802),
            .ltout(n16802_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_5_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_5_7_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0__i5_LC_5_7_4  (
            .in0(N__23158),
            .in1(_gnd_net_),
            .in2(N__20670),
            .in3(N__26495),
            .lcout(data_in_frame_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_444_LC_5_7_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_444_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_444_LC_5_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_444_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__26191),
            .in2(_gnd_net_),
            .in3(N__20653),
            .lcout(\c0.n10569 ),
            .ltout(\c0.n10569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_445_LC_5_7_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_445_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_445_LC_5_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_445_LC_5_7_6  (
            .in0(N__23157),
            .in1(N__26163),
            .in2(N__20667),
            .in3(N__23130),
            .lcout(\c0.n17813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_5_7_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_5_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i2_LC_5_7_7  (
            .in0(N__27111),
            .in1(N__23586),
            .in2(_gnd_net_),
            .in3(N__20654),
            .lcout(data_in_frame_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_5_8_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_5_8_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_5_8_0  (
            .in0(N__26343),
            .in1(N__27993),
            .in2(N__24165),
            .in3(N__26358),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_5_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_5_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i18_LC_5_8_1  (
            .in0(N__27112),
            .in1(N__22645),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(data_in_frame_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_5_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_5_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i45_LC_5_8_2  (
            .in0(N__26496),
            .in1(N__25826),
            .in2(_gnd_net_),
            .in3(N__23625),
            .lcout(data_in_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_5_8_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_5_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_5_8_3  (
            .in0(N__20640),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_410_LC_5_8_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_410_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_410_LC_5_8_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_410_LC_5_8_4  (
            .in0(N__27853),
            .in1(N__26870),
            .in2(_gnd_net_),
            .in3(N__26976),
            .lcout(n12600),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_adj_406_LC_5_8_5 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_adj_406_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_adj_406_LC_5_8_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_adj_406_LC_5_8_5  (
            .in0(N__25678),
            .in1(N__23453),
            .in2(N__23362),
            .in3(N__23210),
            .lcout(n11058),
            .ltout(n11058_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_5_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_5_8_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0__i41_LC_5_8_6  (
            .in0(N__26628),
            .in1(_gnd_net_),
            .in2(N__20862),
            .in3(N__26222),
            .lcout(data_in_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_5_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_5_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i19_LC_5_8_7  (
            .in0(N__26725),
            .in1(N__22684),
            .in2(_gnd_net_),
            .in3(N__26427),
            .lcout(data_in_frame_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_623_LC_5_9_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_623_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_623_LC_5_9_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i8_4_lut_adj_623_LC_5_9_0  (
            .in0(N__26550),
            .in1(N__23922),
            .in2(N__23976),
            .in3(N__23982),
            .lcout(n63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_809_LC_5_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_809_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_809_LC_5_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_809_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__22336),
            .in2(_gnd_net_),
            .in3(N__22493),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_5_9_2 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \c0.i1_3_lut_LC_5_9_2  (
            .in0(N__33178),
            .in1(N__21165),
            .in2(_gnd_net_),
            .in3(N__21253),
            .lcout(\c0.n1502 ),
            .ltout(\c0.n1502_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_454_LC_5_9_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_454_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_454_LC_5_9_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_454_LC_5_9_3  (
            .in0(N__21371),
            .in1(N__20977),
            .in2(N__20820),
            .in3(N__20817),
            .lcout(\c0.n4_adj_2266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_561_LC_5_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_561_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_561_LC_5_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_561_LC_5_9_4  (
            .in0(N__21169),
            .in1(N__21252),
            .in2(_gnd_net_),
            .in3(N__21370),
            .lcout(\c0.n13033 ),
            .ltout(\c0.n13033_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10975_2_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \c0.i10975_2_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10975_2_lut_LC_5_9_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i10975_2_lut_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20769),
            .in3(N__20765),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10976_2_lut_LC_5_9_6 .C_ON=1'b0;
    defparam \c0.i10976_2_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10976_2_lut_LC_5_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10976_2_lut_LC_5_9_6  (
            .in0(N__22494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20721),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10977_2_lut_LC_5_9_7 .C_ON=1'b0;
    defparam \c0.i10977_2_lut_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10977_2_lut_LC_5_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10977_2_lut_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__22282),
            .in2(_gnd_net_),
            .in3(N__22495),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10986_2_lut_3_lut_4_lut_LC_5_10_0 .C_ON=1'b0;
    defparam \c0.i10986_2_lut_3_lut_4_lut_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10986_2_lut_3_lut_4_lut_LC_5_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10986_2_lut_3_lut_4_lut_LC_5_10_0  (
            .in0(N__21396),
            .in1(N__21047),
            .in2(N__21289),
            .in3(N__21168),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_763_LC_5_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_763_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_763_LC_5_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_763_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__20984),
            .in2(_gnd_net_),
            .in3(N__22496),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_5_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_5_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i42_LC_5_10_2  (
            .in0(N__27121),
            .in1(N__25349),
            .in2(_gnd_net_),
            .in3(N__23636),
            .lcout(data_in_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49723),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_609_LC_5_10_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_609_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_609_LC_5_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_609_LC_5_10_3  (
            .in0(N__23715),
            .in1(N__24027),
            .in2(N__24054),
            .in3(N__24006),
            .lcout(n63_adj_2534),
            .ltout(n63_adj_2534_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10988_2_lut_3_lut_4_lut_LC_5_10_4 .C_ON=1'b0;
    defparam \c0.i10988_2_lut_3_lut_4_lut_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10988_2_lut_3_lut_4_lut_LC_5_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10988_2_lut_3_lut_4_lut_LC_5_10_4  (
            .in0(N__21397),
            .in1(N__21272),
            .in2(N__20883),
            .in3(N__24705),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_LC_5_10_5 .C_ON=1'b0;
    defparam \c0.i4_3_lut_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_LC_5_10_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i4_3_lut_LC_5_10_5  (
            .in0(N__23714),
            .in1(N__24015),
            .in2(_gnd_net_),
            .in3(N__26919),
            .lcout(\c0.n63_adj_2262 ),
            .ltout(\c0.n63_adj_2262_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4650_2_lut_LC_5_10_6 .C_ON=1'b0;
    defparam \c0.i4650_2_lut_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4650_2_lut_LC_5_10_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i4650_2_lut_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20871),
            .in3(N__21166),
            .lcout(\c0.n7199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_515_LC_5_10_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_515_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_515_LC_5_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_515_LC_5_10_7  (
            .in0(N__21167),
            .in1(N__21398),
            .in2(N__21978),
            .in3(N__21271),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_5_11_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i5_LC_5_11_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_5_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__24599),
            .in2(_gnd_net_),
            .in3(N__21993),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49711),
            .ce(),
            .sr(N__21987));
    defparam \c0.select_284_Select_5_i3_2_lut_3_lut_4_lut_LC_5_11_2 .C_ON=1'b0;
    defparam \c0.select_284_Select_5_i3_2_lut_3_lut_4_lut_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_5_i3_2_lut_3_lut_4_lut_LC_5_11_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_5_i3_2_lut_3_lut_4_lut_LC_5_11_2  (
            .in0(N__21814),
            .in1(N__21970),
            .in2(N__21717),
            .in3(N__21452),
            .lcout(\c0.n3_adj_2336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_599_LC_5_11_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_599_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_599_LC_5_11_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_599_LC_5_11_3  (
            .in0(N__21969),
            .in1(N__21735),
            .in2(_gnd_net_),
            .in3(N__22335),
            .lcout(\c0.n10_adj_2378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_524_LC_5_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_524_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_524_LC_5_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_524_LC_5_11_4  (
            .in0(N__21173),
            .in1(N__21276),
            .in2(N__21745),
            .in3(N__21449),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_3_i3_2_lut_3_lut_4_lut_LC_5_11_5 .C_ON=1'b0;
    defparam \c0.select_284_Select_3_i3_2_lut_3_lut_4_lut_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_3_i3_2_lut_3_lut_4_lut_LC_5_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.select_284_Select_3_i3_2_lut_3_lut_4_lut_LC_5_11_5  (
            .in0(N__21450),
            .in1(N__21701),
            .in2(N__22343),
            .in3(N__21812),
            .lcout(\c0.n3_adj_2340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_284_Select_4_i3_2_lut_3_lut_4_lut_LC_5_11_6 .C_ON=1'b0;
    defparam \c0.select_284_Select_4_i3_2_lut_3_lut_4_lut_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_284_Select_4_i3_2_lut_3_lut_4_lut_LC_5_11_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.select_284_Select_4_i3_2_lut_3_lut_4_lut_LC_5_11_6  (
            .in0(N__21813),
            .in1(N__21747),
            .in2(N__21716),
            .in3(N__21451),
            .lcout(\c0.n3_adj_2338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_560_LC_5_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_560_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_560_LC_5_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_560_LC_5_11_7  (
            .in0(N__21448),
            .in1(N__25648),
            .in2(N__21290),
            .in3(N__21174),
            .lcout(\c0.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__0__2184_LC_5_12_0 .C_ON=1'b0;
    defparam \c0.data_out_9__0__2184_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__0__2184_LC_5_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_9__0__2184_LC_5_12_0  (
            .in0(N__32412),
            .in1(N__36993),
            .in2(_gnd_net_),
            .in3(N__37407),
            .lcout(\c0.data_out_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49701),
            .ce(N__46845),
            .sr(_gnd_net_));
    defparam \c0.i10993_2_lut_LC_5_12_1 .C_ON=1'b0;
    defparam \c0.i10993_2_lut_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10993_2_lut_LC_5_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10993_2_lut_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__21104),
            .in2(_gnd_net_),
            .in3(N__22528),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10994_2_lut_LC_5_12_2 .C_ON=1'b0;
    defparam \c0.i10994_2_lut_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10994_2_lut_LC_5_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10994_2_lut_LC_5_12_2  (
            .in0(N__22529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10997_2_lut_LC_5_12_3 .C_ON=1'b0;
    defparam \c0.i10997_2_lut_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10997_2_lut_LC_5_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10997_2_lut_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__22224),
            .in2(_gnd_net_),
            .in3(N__22530),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11001_2_lut_LC_5_12_4 .C_ON=1'b0;
    defparam \c0.i11001_2_lut_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11001_2_lut_LC_5_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i11001_2_lut_LC_5_12_4  (
            .in0(N__22531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22168),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_724_LC_5_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_724_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_724_LC_5_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_724_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__23446),
            .in2(_gnd_net_),
            .in3(N__22532),
            .lcout(\c0.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_5_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__24630),
            .in2(_gnd_net_),
            .in3(N__22104),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49694),
            .ce(),
            .sr(N__22098));
    defparam \c0.i1_2_lut_adj_600_LC_5_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_600_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_600_LC_5_13_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i1_2_lut_adj_600_LC_5_13_1  (
            .in0(N__22383),
            .in1(N__22056),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n26_adj_2379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_608_LC_5_13_2 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_608_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_608_LC_5_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_adj_608_LC_5_13_2  (
            .in0(N__22275),
            .in1(N__22617),
            .in2(N__22086),
            .in3(N__22027),
            .lcout(\c0.n44_adj_2382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10996_2_lut_LC_5_13_3 .C_ON=1'b0;
    defparam \c0.i10996_2_lut_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10996_2_lut_LC_5_13_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i10996_2_lut_LC_5_13_3  (
            .in0(N__22565),
            .in1(N__22057),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10985_2_lut_LC_5_13_4 .C_ON=1'b0;
    defparam \c0.i10985_2_lut_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10985_2_lut_LC_5_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10985_2_lut_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__22028),
            .in2(_gnd_net_),
            .in3(N__22563),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10995_2_lut_LC_5_13_5 .C_ON=1'b0;
    defparam \c0.i10995_2_lut_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10995_2_lut_LC_5_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10995_2_lut_LC_5_13_5  (
            .in0(N__22564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22619),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10978_2_lut_LC_5_13_6 .C_ON=1'b0;
    defparam \c0.i10978_2_lut_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10978_2_lut_LC_5_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10978_2_lut_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__22384),
            .in2(_gnd_net_),
            .in3(N__22561),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10979_2_lut_LC_5_13_7 .C_ON=1'b0;
    defparam \c0.i10979_2_lut_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10979_2_lut_LC_5_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10979_2_lut_LC_5_13_7  (
            .in0(N__22562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22440),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i27_LC_5_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i27_LC_5_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_5_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__24631),
            .in2(_gnd_net_),
            .in3(N__22404),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(N__22368));
    defparam \c0.FRAME_MATCHER_i_i3_LC_5_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i3_LC_5_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_5_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__24633),
            .in2(_gnd_net_),
            .in3(N__22356),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49683),
            .ce(),
            .sr(N__22308));
    defparam \c0.FRAME_MATCHER_i_i28_LC_5_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i28_LC_5_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_5_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__22296),
            .in2(_gnd_net_),
            .in3(N__24644),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49679),
            .ce(),
            .sr(N__22248));
    defparam i15182_4_lut_LC_5_23_2.C_ON=1'b0;
    defparam i15182_4_lut_LC_5_23_2.SEQ_MODE=4'b0000;
    defparam i15182_4_lut_LC_5_23_2.LUT_INIT=16'b1011101100100000;
    LogicCell40 i15182_4_lut_LC_5_23_2 (
            .in0(N__24983),
            .in1(N__24944),
            .in2(N__24966),
            .in3(N__24824),
            .lcout(n18043),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15183_4_lut_LC_5_23_3.C_ON=1'b0;
    defparam i15183_4_lut_LC_5_23_3.SEQ_MODE=4'b0000;
    defparam i15183_4_lut_LC_5_23_3.LUT_INIT=16'b1111100011101100;
    LogicCell40 i15183_4_lut_LC_5_23_3 (
            .in0(N__24945),
            .in1(N__24965),
            .in2(N__24828),
            .in3(N__24984),
            .lcout(n18044),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15184_3_lut_LC_5_24_4.C_ON=1'b0;
    defparam i15184_3_lut_LC_5_24_4.SEQ_MODE=4'b0000;
    defparam i15184_3_lut_LC_5_24_4.LUT_INIT=16'b0011001101010101;
    LogicCell40 i15184_3_lut_LC_5_24_4 (
            .in0(N__22821),
            .in1(N__22815),
            .in2(_gnd_net_),
            .in3(N__24924),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.PHASES_i3_LC_5_28_0 .C_ON=1'b0;
    defparam \control.PHASES_i3_LC_5_28_0 .SEQ_MODE=4'b1000;
    defparam \control.PHASES_i3_LC_5_28_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \control.PHASES_i3_LC_5_28_0  (
            .in0(N__35656),
            .in1(N__35461),
            .in2(_gnd_net_),
            .in3(N__35511),
            .lcout(PIN_3_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49773),
            .ce(N__24912),
            .sr(N__35347));
    defparam \c0.byte_transmit_counter2_i7_LC_6_1_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i7_LC_6_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i7_LC_6_1_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i7_LC_6_1_0  (
            .in0(N__25164),
            .in1(N__25225),
            .in2(N__30658),
            .in3(N__30555),
            .lcout(\c0.byte_transmit_counter2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49842),
            .ce(),
            .sr(N__25026));
    defparam \c0.byte_transmit_counter2_i2_LC_6_2_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i2_LC_6_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i2_LC_6_2_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i2_LC_6_2_0  (
            .in0(N__24993),
            .in1(N__47981),
            .in2(N__30657),
            .in3(N__30547),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(N__22785));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_6_2_2 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_6_2_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_6_2_2  (
            .in0(N__22770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i3_LC_6_3_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i3_LC_6_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i3_LC_6_3_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i3_LC_6_3_0  (
            .in0(N__25317),
            .in1(N__49027),
            .in2(N__30643),
            .in3(N__30546),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49825),
            .ce(),
            .sr(N__22722));
    defparam \c0.data_in_frame_0__i50_LC_6_4_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_6_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_6_4_0  (
            .in0(N__27106),
            .in1(N__22835),
            .in2(_gnd_net_),
            .in3(N__25860),
            .lcout(data_in_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_6_4_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_6_4_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_in_frame_0__i28_LC_6_4_1  (
            .in0(N__22706),
            .in1(N__25706),
            .in2(N__25785),
            .in3(N__25550),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_700_LC_6_4_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_700_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_700_LC_6_4_2 .LUT_INIT=16'b1101111111111101;
    LogicCell40 \c0.i9_4_lut_adj_700_LC_6_4_2  (
            .in0(N__22692),
            .in1(N__22662),
            .in2(N__22656),
            .in3(N__26013),
            .lcout(),
            .ltout(\c0.n23_adj_2420_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_703_LC_6_4_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_703_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_703_LC_6_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i13_4_lut_adj_703_LC_6_4_3  (
            .in0(N__22893),
            .in1(N__22887),
            .in2(N__22875),
            .in3(N__23061),
            .lcout(\c0.n4494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_adj_412_LC_6_4_4 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_adj_412_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_adj_412_LC_6_4_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_adj_412_LC_6_4_4  (
            .in0(N__25705),
            .in1(N__23466),
            .in2(N__23367),
            .in3(N__23226),
            .lcout(n16797),
            .ltout(n16797_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_6_4_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_6_4_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0__i54_LC_6_4_5  (
            .in0(N__27211),
            .in1(_gnd_net_),
            .in2(N__22872),
            .in3(N__25416),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_6_4_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_6_4_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_in_frame_0__i30_LC_6_4_6  (
            .in0(N__25551),
            .in1(N__27212),
            .in2(N__25716),
            .in3(N__22868),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_6_4_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_6_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i52_LC_6_4_7  (
            .in0(N__25861),
            .in1(N__25784),
            .in2(_gnd_net_),
            .in3(N__23537),
            .lcout(data_in_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_6_5_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_6_5_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i15_LC_6_5_0  (
            .in0(N__25546),
            .in1(N__25713),
            .in2(N__27627),
            .in3(N__22927),
            .lcout(\c0.data_in_frame_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_LC_6_5_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_LC_6_5_1  (
            .in0(N__23461),
            .in1(N__23360),
            .in2(_gnd_net_),
            .in3(N__23220),
            .lcout(\c0.rx.n129 ),
            .ltout(\c0.rx.n129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_6_5_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_6_5_2 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \c0.data_in_frame_0__i32_LC_6_5_2  (
            .in0(N__22850),
            .in1(N__25715),
            .in2(N__22854),
            .in3(N__24178),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_6_5_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_6_5_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i12_LC_6_5_3  (
            .in0(N__25712),
            .in1(N__26303),
            .in2(N__25782),
            .in3(N__25544),
            .lcout(\c0.data_in_frame_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_642_LC_6_5_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_642_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_642_LC_6_5_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_642_LC_6_5_4  (
            .in0(N__22977),
            .in1(N__22926),
            .in2(N__22836),
            .in3(N__23028),
            .lcout(\c0.n16994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_6_5_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_6_5_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i11_LC_6_5_5  (
            .in0(N__25711),
            .in1(N__25477),
            .in2(N__26727),
            .in3(N__25543),
            .lcout(\c0.data_in_frame_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_6_5_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_6_5_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i14_LC_6_5_6  (
            .in0(N__25545),
            .in1(N__27216),
            .in2(N__22985),
            .in3(N__25714),
            .lcout(\c0.data_in_frame_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_6_5_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_6_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i56_LC_6_5_7  (
            .in0(N__24177),
            .in1(N__23052),
            .in2(_gnd_net_),
            .in3(N__25863),
            .lcout(data_in_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_628_LC_6_6_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_628_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_628_LC_6_6_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_628_LC_6_6_0  (
            .in0(N__23039),
            .in1(N__26297),
            .in2(N__25478),
            .in3(N__25872),
            .lcout(\c0.n10761 ),
            .ltout(\c0.n10761_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_629_LC_6_6_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_629_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_629_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_629_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__23010),
            .in2(N__22992),
            .in3(N__23514),
            .lcout(\c0.n17733 ),
            .ltout(\c0.n17733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_632_LC_6_6_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_632_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_632_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_632_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__22976),
            .in2(N__22953),
            .in3(N__22949),
            .lcout(\c0.n17735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_641_LC_6_6_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_641_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_641_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_641_LC_6_6_3  (
            .in0(N__23481),
            .in1(N__26068),
            .in2(_gnd_net_),
            .in3(N__26042),
            .lcout(\c0.n17722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_645_LC_6_6_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_645_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_645_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_645_LC_6_6_4  (
            .in0(N__23690),
            .in1(N__22922),
            .in2(_gnd_net_),
            .in3(N__22899),
            .lcout(),
            .ltout(\c0.n17734_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15141_4_lut_LC_6_6_5 .C_ON=1'b0;
    defparam \c0.i15141_4_lut_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15141_4_lut_LC_6_6_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \c0.i15141_4_lut_LC_6_6_5  (
            .in0(N__23554),
            .in1(N__23538),
            .in2(N__23523),
            .in3(N__23515),
            .lcout(),
            .ltout(\c0.n18000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_672_LC_6_6_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_672_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_672_LC_6_6_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i13_4_lut_adj_672_LC_6_6_6  (
            .in0(N__23496),
            .in1(N__23490),
            .in2(N__23484),
            .in3(N__26268),
            .lcout(\c0.n29_adj_2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_6_7_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_6_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i43_LC_6_7_0  (
            .in0(N__23480),
            .in1(N__26704),
            .in2(_gnd_net_),
            .in3(N__23633),
            .lcout(data_in_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_407_LC_6_7_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_407_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_407_LC_6_7_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_4_lut_adj_407_LC_6_7_1  (
            .in0(N__23460),
            .in1(N__25710),
            .in2(N__23361),
            .in3(N__23222),
            .lcout(n120),
            .ltout(n120_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_6_7_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_6_7_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0__i20_LC_6_7_2  (
            .in0(N__25763),
            .in1(_gnd_net_),
            .in2(N__23184),
            .in3(N__23179),
            .lcout(data_in_frame_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1012_2_lut_LC_6_7_3 .C_ON=1'b0;
    defparam \c0.i1012_2_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1012_2_lut_LC_6_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1012_2_lut_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__23159),
            .in2(_gnd_net_),
            .in3(N__23131),
            .lcout(\c0.n2124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_6_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_6_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i3_LC_6_7_4  (
            .in0(N__26196),
            .in1(N__23589),
            .in2(_gnd_net_),
            .in3(N__26703),
            .lcout(data_in_frame_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_699_LC_6_7_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_699_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_699_LC_6_7_5 .LUT_INIT=16'b1111110111011111;
    LogicCell40 \c0.i8_4_lut_adj_699_LC_6_7_5  (
            .in0(N__23108),
            .in1(N__23091),
            .in2(N__23678),
            .in3(N__23085),
            .lcout(\c0.n22_adj_2419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_6_7_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_6_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i7_LC_6_7_6  (
            .in0(N__27604),
            .in1(N__23590),
            .in2(_gnd_net_),
            .in3(N__25909),
            .lcout(data_in_frame_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_6_7_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_6_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_frame_0__i48_LC_6_7_7  (
            .in0(N__23634),
            .in1(N__24154),
            .in2(_gnd_net_),
            .in3(N__23691),
            .lcout(data_in_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_6_8_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_6_8_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_6_8_0  (
            .in0(N__27429),
            .in1(N__27938),
            .in2(N__28135),
            .in3(N__26967),
            .lcout(\c0.rx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_6_8_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_6_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i24_LC_6_8_1  (
            .in0(N__24153),
            .in1(N__23674),
            .in2(_gnd_net_),
            .in3(N__26425),
            .lcout(data_in_frame_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_423_LC_6_8_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_423_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_423_LC_6_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_423_LC_6_8_2  (
            .in0(N__28102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27981),
            .lcout(\c0.rx.n17702 ),
            .ltout(\c0.rx.n17702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_6_8_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_6_8_3 .LUT_INIT=16'b1101100011011100;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_6_8_3  (
            .in0(N__26733),
            .in1(N__26629),
            .in2(N__23652),
            .in3(N__28106),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_adj_400_LC_6_8_4 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_adj_400_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_adj_400_LC_6_8_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.rx.i3_4_lut_adj_400_LC_6_8_4  (
            .in0(N__27539),
            .in1(N__27796),
            .in2(N__23649),
            .in3(N__26661),
            .lcout(),
            .ltout(\c0.rx.n17704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_8_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_8_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__27187),
            .in2(N__23640),
            .in3(N__26367),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_6_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_6_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i44_LC_6_8_6  (
            .in0(N__25779),
            .in1(N__25493),
            .in2(_gnd_net_),
            .in3(N__23626),
            .lcout(data_in_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_6_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_6_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i4_LC_6_8_7  (
            .in0(N__26170),
            .in1(N__23592),
            .in2(_gnd_net_),
            .in3(N__25780),
            .lcout(data_in_frame_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15143_4_lut_LC_6_9_0 .C_ON=1'b0;
    defparam \c0.i15143_4_lut_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15143_4_lut_LC_6_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15143_4_lut_LC_6_9_0  (
            .in0(N__23937),
            .in1(N__27060),
            .in2(N__26574),
            .in3(N__23998),
            .lcout(),
            .ltout(\c0.n18002_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_582_LC_6_9_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_582_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_582_LC_6_9_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i3_4_lut_adj_582_LC_6_9_1  (
            .in0(N__23967),
            .in1(N__26545),
            .in2(N__23718),
            .in3(N__34048),
            .lcout(\c0.n10498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4__2265_LC_6_9_2 .C_ON=1'b0;
    defparam \c0.data_in_3__4__2265_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4__2265_LC_6_9_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_3__4__2265_LC_6_9_2  (
            .in0(N__23938),
            .in1(_gnd_net_),
            .in2(N__34221),
            .in3(N__26501),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4__2281_LC_6_9_3 .C_ON=1'b0;
    defparam \c0.data_in_1__4__2281_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4__2281_LC_6_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_1__4__2281_LC_6_9_3  (
            .in0(N__23968),
            .in1(N__34198),
            .in2(_gnd_net_),
            .in3(N__24080),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_6_9_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_6_9_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.rx.i1_4_lut_LC_6_9_4  (
            .in0(N__27410),
            .in1(N__27920),
            .in2(N__28154),
            .in3(N__26958),
            .lcout(\c0.rx.n10988 ),
            .ltout(\c0.rx.n10988_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i9849_3_lut_4_lut_LC_6_9_5 .C_ON=1'b0;
    defparam \c0.rx.i9849_3_lut_4_lut_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i9849_3_lut_4_lut_LC_6_9_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \c0.rx.i9849_3_lut_4_lut_LC_6_9_5  (
            .in0(N__27854),
            .in1(N__27528),
            .in2(N__23706),
            .in3(N__26863),
            .lcout(),
            .ltout(\c0.rx.n12624_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_6_9_6 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_6_9_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_6_9_6  (
            .in0(N__28148),
            .in1(N__24041),
            .in2(N__23703),
            .in3(N__27855),
            .lcout(\c0.rx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5__2288_LC_6_9_7 .C_ON=1'b0;
    defparam \c0.data_in_0__5__2288_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5__2288_LC_6_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0__5__2288_LC_6_9_7  (
            .in0(N__23999),
            .in1(N__34197),
            .in2(_gnd_net_),
            .in3(N__24102),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2__2291_LC_6_10_0 .C_ON=1'b0;
    defparam \c0.data_in_0__2__2291_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2__2291_LC_6_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__2__2291_LC_6_10_0  (
            .in0(N__26902),
            .in1(N__34212),
            .in2(_gnd_net_),
            .in3(N__23700),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_570_LC_6_10_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_570_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_570_LC_6_10_1 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.i9_4_lut_adj_570_LC_6_10_1  (
            .in0(N__23699),
            .in1(N__23948),
            .in2(N__26886),
            .in3(N__24060),
            .lcout(),
            .ltout(\c0.n20_adj_2371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_580_LC_6_10_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_580_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_580_LC_6_10_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i10_4_lut_adj_580_LC_6_10_2  (
            .in0(N__26749),
            .in1(N__34280),
            .in2(N__24018),
            .in3(N__26910),
            .lcout(\c0.n10516 ),
            .ltout(\c0.n10516_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_581_LC_6_10_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_581_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_581_LC_6_10_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i3_4_lut_adj_581_LC_6_10_3  (
            .in0(N__26523),
            .in1(N__29278),
            .in2(N__24009),
            .in3(N__26901),
            .lcout(\c0.n10367 ),
            .ltout(\c0.n10367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_622_LC_6_10_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_622_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_622_LC_6_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_622_LC_6_10_4  (
            .in0(N__24000),
            .in1(N__23939),
            .in2(N__23985),
            .in3(N__27061),
            .lcout(\c0.n15_adj_2389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4__2289_LC_6_10_5 .C_ON=1'b0;
    defparam \c0.data_in_0__4__2289_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4__2289_LC_6_10_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0__4__2289_LC_6_10_5  (
            .in0(N__23972),
            .in1(_gnd_net_),
            .in2(N__34228),
            .in3(N__23949),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4__2273_LC_6_10_6 .C_ON=1'b0;
    defparam \c0.data_in_2__4__2273_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4__2273_LC_6_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__4__2273_LC_6_10_6  (
            .in0(N__24079),
            .in1(N__23940),
            .in2(_gnd_net_),
            .in3(N__34216),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_619_LC_6_10_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_619_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_619_LC_6_10_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.i5_3_lut_adj_619_LC_6_10_7  (
            .in0(N__34049),
            .in1(N__26571),
            .in2(_gnd_net_),
            .in3(N__26769),
            .lcout(\c0.n14_adj_2388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3__2282_LC_6_11_0 .C_ON=1'b0;
    defparam \c0.data_in_1__3__2282_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3__2282_LC_6_11_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__3__2282_LC_6_11_0  (
            .in0(N__34050),
            .in1(N__34127),
            .in2(_gnd_net_),
            .in3(N__27689),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5__2280_LC_6_11_1 .C_ON=1'b0;
    defparam \c0.data_in_1__5__2280_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5__2280_LC_6_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_1__5__2280_LC_6_11_1  (
            .in0(N__24101),
            .in1(N__34186),
            .in2(_gnd_net_),
            .in3(N__24197),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15770_1_lut_LC_6_11_2 .C_ON=1'b0;
    defparam \c0.rx.i15770_1_lut_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15770_1_lut_LC_6_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.rx.i15770_1_lut_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34126),
            .lcout(\c0.n18631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15148_3_lut_LC_6_11_3 .C_ON=1'b0;
    defparam \c0.i15148_3_lut_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15148_3_lut_LC_6_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i15148_3_lut_LC_6_11_3  (
            .in0(N__24213),
            .in1(N__24195),
            .in2(_gnd_net_),
            .in3(N__27658),
            .lcout(\c0.n18008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_569_LC_6_11_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_569_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_569_LC_6_11_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i7_4_lut_adj_569_LC_6_11_4  (
            .in0(N__24097),
            .in1(N__34297),
            .in2(N__24081),
            .in3(N__27688),
            .lcout(\c0.n18_adj_2370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_604_LC_6_11_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_604_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_604_LC_6_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_604_LC_6_11_5  (
            .in0(N__24214),
            .in1(N__24196),
            .in2(N__26808),
            .in3(N__27659),
            .lcout(\c0.n13_adj_2380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3__2266_LC_6_11_6 .C_ON=1'b0;
    defparam \c0.data_in_3__3__2266_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3__2266_LC_6_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_3__3__2266_LC_6_11_6  (
            .in0(N__34250),
            .in1(N__25783),
            .in2(_gnd_net_),
            .in3(N__34128),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6__2263_LC_6_11_7 .C_ON=1'b0;
    defparam \c0.data_in_3__6__2263_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6__2263_LC_6_11_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__6__2263_LC_6_11_7  (
            .in0(N__27587),
            .in1(N__34187),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_6_12_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_6_12_0 .LUT_INIT=16'b0100100011110000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_6_12_0  (
            .in0(N__26871),
            .in1(N__28082),
            .in2(N__27540),
            .in3(N__24045),
            .lcout(\c0.rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7__2270_LC_6_12_1 .C_ON=1'b0;
    defparam \c0.data_in_2__7__2270_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7__2270_LC_6_12_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_2__7__2270_LC_6_12_1  (
            .in0(N__27714),
            .in1(N__34185),
            .in2(_gnd_net_),
            .in3(N__24215),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15146_4_lut_LC_6_12_2 .C_ON=1'b0;
    defparam \c0.i15146_4_lut_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15146_4_lut_LC_6_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15146_4_lut_LC_6_12_2  (
            .in0(N__27254),
            .in1(N__27728),
            .in2(N__27156),
            .in3(N__27712),
            .lcout(),
            .ltout(\c0.n18006_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_589_LC_6_12_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_589_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_589_LC_6_12_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i6_4_lut_adj_589_LC_6_12_3  (
            .in0(N__27031),
            .in1(N__27001),
            .in2(N__24030),
            .in3(N__27675),
            .lcout(\c0.n14_adj_2375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7__2278_LC_6_12_4 .C_ON=1'b0;
    defparam \c0.data_in_1__7__2278_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7__2278_LC_6_12_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_1__7__2278_LC_6_12_4  (
            .in0(N__24216),
            .in1(_gnd_net_),
            .in2(N__27008),
            .in3(N__34183),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5__2272_LC_6_12_5 .C_ON=1'b0;
    defparam \c0.data_in_2__5__2272_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5__2272_LC_6_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__5__2272_LC_6_12_5  (
            .in0(N__34181),
            .in1(N__27155),
            .in2(_gnd_net_),
            .in3(N__24198),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7__2262_LC_6_12_6 .C_ON=1'b0;
    defparam \c0.data_in_3__7__2262_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7__2262_LC_6_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__7__2262_LC_6_12_6  (
            .in0(N__24179),
            .in1(N__34182),
            .in2(_gnd_net_),
            .in3(N__27713),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__0__2293_LC_6_12_7 .C_ON=1'b0;
    defparam \c0.data_in_0__0__2293_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0__2293_LC_6_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0__0__2293_LC_6_12_7  (
            .in0(N__27729),
            .in1(N__34184),
            .in2(_gnd_net_),
            .in3(N__26757),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_6_13_0 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__28199),
            .in2(_gnd_net_),
            .in3(N__24117),
            .lcout(\c0.rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\c0.rx.n16532 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i1_LC_6_13_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__27354),
            .in2(_gnd_net_),
            .in3(N__24114),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.rx.n16532 ),
            .carryout(\c0.rx.n16533 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i2_LC_6_13_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i2_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_6_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__27336),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.rx.n16533 ),
            .carryout(\c0.rx.n16534 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i3_LC_6_13_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__27317),
            .in2(_gnd_net_),
            .in3(N__24108),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.rx.n16534 ),
            .carryout(\c0.rx.n16535 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i4_LC_6_13_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i4_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_6_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__27294),
            .in2(_gnd_net_),
            .in3(N__24105),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.rx.n16535 ),
            .carryout(\c0.rx.n16536 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i5_LC_6_13_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__28253),
            .in2(_gnd_net_),
            .in3(N__24279),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.rx.n16536 ),
            .carryout(\c0.rx.n16537 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i6_LC_6_13_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i6_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_6_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__29177),
            .in2(_gnd_net_),
            .in3(N__24276),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.rx.n16537 ),
            .carryout(\c0.rx.n16538 ),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.r_Clock_Count__i7_LC_6_13_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__29204),
            .in2(_gnd_net_),
            .in3(N__24273),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49702),
            .ce(N__24729),
            .sr(N__24270));
    defparam \c0.rx.i1_2_lut_adj_399_LC_6_14_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_399_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_399_LC_6_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_399_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__27447),
            .in2(_gnd_net_),
            .in3(N__24222),
            .lcout(\c0.rx.n12819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15562_2_lut_LC_6_14_1 .C_ON=1'b0;
    defparam \c0.i15562_2_lut_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15562_2_lut_LC_6_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15562_2_lut_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__39036),
            .in2(_gnd_net_),
            .in3(N__47412),
            .lcout(),
            .ltout(\c0.n18225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1__2207_LC_6_14_2 .C_ON=1'b0;
    defparam \c0.data_out_6__1__2207_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1__2207_LC_6_14_2 .LUT_INIT=16'b1111001111010001;
    LogicCell40 \c0.data_out_6__1__2207_LC_6_14_2  (
            .in0(N__47689),
            .in1(N__47122),
            .in2(N__24261),
            .in3(N__42498),
            .lcout(\c0.data_out_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49695),
            .ce(N__43423),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_408_LC_6_14_3 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_408_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_408_LC_6_14_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_4_lut_adj_408_LC_6_14_3  (
            .in0(N__29200),
            .in1(N__29173),
            .in2(N__28196),
            .in3(N__28224),
            .lcout(),
            .ltout(\c0.rx.n15905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i21_4_lut_LC_6_14_4 .C_ON=1'b0;
    defparam \c0.rx.i21_4_lut_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i21_4_lut_LC_6_14_4 .LUT_INIT=16'b1010101000111010;
    LogicCell40 \c0.rx.i21_4_lut_LC_6_14_4  (
            .in0(N__24258),
            .in1(N__24243),
            .in2(N__24228),
            .in3(N__28250),
            .lcout(),
            .ltout(\c0.rx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13229_4_lut_LC_6_14_5 .C_ON=1'b0;
    defparam \c0.rx.i13229_4_lut_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13229_4_lut_LC_6_14_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \c0.rx.i13229_4_lut_LC_6_14_5  (
            .in0(N__28119),
            .in1(N__28161),
            .in2(N__24225),
            .in3(N__29154),
            .lcout(\c0.rx.n12 ),
            .ltout(\c0.rx.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15076_4_lut_LC_6_14_6 .C_ON=1'b0;
    defparam \c0.rx.i15076_4_lut_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15076_4_lut_LC_6_14_6 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \c0.rx.i15076_4_lut_LC_6_14_6  (
            .in0(N__28286),
            .in1(N__27876),
            .in2(N__24732),
            .in3(N__27448),
            .lcout(\c0.rx.n11082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__24645),
            .in2(_gnd_net_),
            .in3(N__24717),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(N__24660));
    defparam \c0.FRAME_MATCHER_i_i13_LC_6_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i13_LC_6_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_6_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__24620),
            .in2(_gnd_net_),
            .in3(N__24393),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49684),
            .ce(),
            .sr(N__24345));
    defparam blink_counter_2483__i0_LC_6_21_0.C_ON=1'b1;
    defparam blink_counter_2483__i0_LC_6_21_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i0_LC_6_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i0_LC_6_21_0 (
            .in0(_gnd_net_),
            .in1(N__24330),
            .in2(_gnd_net_),
            .in3(N__24324),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(n16609),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i1_LC_6_21_1.C_ON=1'b1;
    defparam blink_counter_2483__i1_LC_6_21_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i1_LC_6_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i1_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__24321),
            .in2(_gnd_net_),
            .in3(N__24315),
            .lcout(n25),
            .ltout(),
            .carryin(n16609),
            .carryout(n16610),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i2_LC_6_21_2.C_ON=1'b1;
    defparam blink_counter_2483__i2_LC_6_21_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i2_LC_6_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i2_LC_6_21_2 (
            .in0(_gnd_net_),
            .in1(N__24312),
            .in2(_gnd_net_),
            .in3(N__24306),
            .lcout(n24),
            .ltout(),
            .carryin(n16610),
            .carryout(n16611),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i3_LC_6_21_3.C_ON=1'b1;
    defparam blink_counter_2483__i3_LC_6_21_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i3_LC_6_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i3_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__24303),
            .in2(_gnd_net_),
            .in3(N__24297),
            .lcout(n23),
            .ltout(),
            .carryin(n16611),
            .carryout(n16612),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i4_LC_6_21_4.C_ON=1'b1;
    defparam blink_counter_2483__i4_LC_6_21_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i4_LC_6_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i4_LC_6_21_4 (
            .in0(_gnd_net_),
            .in1(N__24294),
            .in2(_gnd_net_),
            .in3(N__24288),
            .lcout(n22_adj_2481),
            .ltout(),
            .carryin(n16612),
            .carryout(n16613),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i5_LC_6_21_5.C_ON=1'b1;
    defparam blink_counter_2483__i5_LC_6_21_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i5_LC_6_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i5_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(N__24285),
            .in2(_gnd_net_),
            .in3(N__24807),
            .lcout(n21),
            .ltout(),
            .carryin(n16613),
            .carryout(n16614),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i6_LC_6_21_6.C_ON=1'b1;
    defparam blink_counter_2483__i6_LC_6_21_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i6_LC_6_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i6_LC_6_21_6 (
            .in0(_gnd_net_),
            .in1(N__24804),
            .in2(_gnd_net_),
            .in3(N__24798),
            .lcout(n20),
            .ltout(),
            .carryin(n16614),
            .carryout(n16615),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i7_LC_6_21_7.C_ON=1'b1;
    defparam blink_counter_2483__i7_LC_6_21_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i7_LC_6_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i7_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__24795),
            .in2(_gnd_net_),
            .in3(N__24789),
            .lcout(n19),
            .ltout(),
            .carryin(n16615),
            .carryout(n16616),
            .clk(N__49703),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i8_LC_6_22_0.C_ON=1'b1;
    defparam blink_counter_2483__i8_LC_6_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i8_LC_6_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i8_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__24786),
            .in2(_gnd_net_),
            .in3(N__24780),
            .lcout(n18_adj_2480),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(n16617),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i9_LC_6_22_1.C_ON=1'b1;
    defparam blink_counter_2483__i9_LC_6_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i9_LC_6_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i9_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(N__24777),
            .in2(_gnd_net_),
            .in3(N__24771),
            .lcout(n17),
            .ltout(),
            .carryin(n16617),
            .carryout(n16618),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i10_LC_6_22_2.C_ON=1'b1;
    defparam blink_counter_2483__i10_LC_6_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i10_LC_6_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i10_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(N__24768),
            .in2(_gnd_net_),
            .in3(N__24762),
            .lcout(n16),
            .ltout(),
            .carryin(n16618),
            .carryout(n16619),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i11_LC_6_22_3.C_ON=1'b1;
    defparam blink_counter_2483__i11_LC_6_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i11_LC_6_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i11_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(N__24759),
            .in2(_gnd_net_),
            .in3(N__24753),
            .lcout(n15_adj_2479),
            .ltout(),
            .carryin(n16619),
            .carryout(n16620),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i12_LC_6_22_4.C_ON=1'b1;
    defparam blink_counter_2483__i12_LC_6_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i12_LC_6_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i12_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(N__24750),
            .in2(_gnd_net_),
            .in3(N__24744),
            .lcout(n14_adj_2478),
            .ltout(),
            .carryin(n16620),
            .carryout(n16621),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i13_LC_6_22_5.C_ON=1'b1;
    defparam blink_counter_2483__i13_LC_6_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i13_LC_6_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i13_LC_6_22_5 (
            .in0(_gnd_net_),
            .in1(N__24741),
            .in2(_gnd_net_),
            .in3(N__24735),
            .lcout(n13),
            .ltout(),
            .carryin(n16621),
            .carryout(n16622),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i14_LC_6_22_6.C_ON=1'b1;
    defparam blink_counter_2483__i14_LC_6_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i14_LC_6_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i14_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(N__24891),
            .in2(_gnd_net_),
            .in3(N__24885),
            .lcout(n12),
            .ltout(),
            .carryin(n16622),
            .carryout(n16623),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i15_LC_6_22_7.C_ON=1'b1;
    defparam blink_counter_2483__i15_LC_6_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i15_LC_6_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i15_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(N__24882),
            .in2(_gnd_net_),
            .in3(N__24876),
            .lcout(n11),
            .ltout(),
            .carryin(n16623),
            .carryout(n16624),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i16_LC_6_23_0.C_ON=1'b1;
    defparam blink_counter_2483__i16_LC_6_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i16_LC_6_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i16_LC_6_23_0 (
            .in0(_gnd_net_),
            .in1(N__24873),
            .in2(_gnd_net_),
            .in3(N__24867),
            .lcout(n10_adj_2467),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(n16625),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i17_LC_6_23_1.C_ON=1'b1;
    defparam blink_counter_2483__i17_LC_6_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i17_LC_6_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i17_LC_6_23_1 (
            .in0(_gnd_net_),
            .in1(N__24864),
            .in2(_gnd_net_),
            .in3(N__24858),
            .lcout(n9),
            .ltout(),
            .carryin(n16625),
            .carryout(n16626),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i18_LC_6_23_2.C_ON=1'b1;
    defparam blink_counter_2483__i18_LC_6_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i18_LC_6_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i18_LC_6_23_2 (
            .in0(_gnd_net_),
            .in1(N__24855),
            .in2(_gnd_net_),
            .in3(N__24849),
            .lcout(n8),
            .ltout(),
            .carryin(n16626),
            .carryout(n16627),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i19_LC_6_23_3.C_ON=1'b1;
    defparam blink_counter_2483__i19_LC_6_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i19_LC_6_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i19_LC_6_23_3 (
            .in0(_gnd_net_),
            .in1(N__24846),
            .in2(_gnd_net_),
            .in3(N__24840),
            .lcout(n7_adj_2476),
            .ltout(),
            .carryin(n16627),
            .carryout(n16628),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i20_LC_6_23_4.C_ON=1'b1;
    defparam blink_counter_2483__i20_LC_6_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i20_LC_6_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i20_LC_6_23_4 (
            .in0(_gnd_net_),
            .in1(N__24837),
            .in2(_gnd_net_),
            .in3(N__24831),
            .lcout(n6),
            .ltout(),
            .carryin(n16628),
            .carryout(n16629),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i21_LC_6_23_5.C_ON=1'b1;
    defparam blink_counter_2483__i21_LC_6_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i21_LC_6_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i21_LC_6_23_5 (
            .in0(_gnd_net_),
            .in1(N__24823),
            .in2(_gnd_net_),
            .in3(N__24810),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n16629),
            .carryout(n16630),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i22_LC_6_23_6.C_ON=1'b1;
    defparam blink_counter_2483__i22_LC_6_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i22_LC_6_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i22_LC_6_23_6 (
            .in0(_gnd_net_),
            .in1(N__24982),
            .in2(_gnd_net_),
            .in3(N__24969),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n16630),
            .carryout(n16631),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i23_LC_6_23_7.C_ON=1'b1;
    defparam blink_counter_2483__i23_LC_6_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i23_LC_6_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i23_LC_6_23_7 (
            .in0(_gnd_net_),
            .in1(N__24961),
            .in2(_gnd_net_),
            .in3(N__24948),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n16631),
            .carryout(n16632),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i24_LC_6_24_0.C_ON=1'b1;
    defparam blink_counter_2483__i24_LC_6_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i24_LC_6_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i24_LC_6_24_0 (
            .in0(_gnd_net_),
            .in1(N__24943),
            .in2(_gnd_net_),
            .in3(N__24930),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(n16633),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2483__i25_LC_6_24_1.C_ON=1'b0;
    defparam blink_counter_2483__i25_LC_6_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2483__i25_LC_6_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2483__i25_LC_6_24_1 (
            .in0(_gnd_net_),
            .in1(N__24923),
            .in2(_gnd_net_),
            .in3(N__24927),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15760_3_lut_LC_6_27_7 .C_ON=1'b0;
    defparam \control.i15760_3_lut_LC_6_27_7 .SEQ_MODE=4'b0000;
    defparam \control.i15760_3_lut_LC_6_27_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \control.i15760_3_lut_LC_6_27_7  (
            .in0(N__28461),
            .in1(N__32907),
            .in2(_gnd_net_),
            .in3(N__32862),
            .lcout(\control.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.PHASES_i1_LC_6_29_1 .C_ON=1'b0;
    defparam \control.PHASES_i1_LC_6_29_1 .SEQ_MODE=4'b1000;
    defparam \control.PHASES_i1_LC_6_29_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \control.PHASES_i1_LC_6_29_1  (
            .in0(N__35638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35441),
            .lcout(PIN_1_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49802),
            .ce(N__35723),
            .sr(N__28446));
    defparam \c0.byte_transmit_counter2_i6_LC_7_1_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i6_LC_7_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i6_LC_7_1_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i6_LC_7_1_0  (
            .in0(N__25239),
            .in1(N__25267),
            .in2(N__30659),
            .in3(N__30552),
            .lcout(\c0.byte_transmit_counter2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49851),
            .ce(),
            .sr(N__25131));
    defparam \c0.i1_2_lut_4_lut_adj_771_LC_7_2_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_771_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_771_LC_7_2_0 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_771_LC_7_2_0  (
            .in0(N__25123),
            .in1(N__25069),
            .in2(N__25305),
            .in3(N__33087),
            .lcout(\c0.n4_adj_2203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11047_3_lut_LC_7_2_1 .C_ON=1'b0;
    defparam \c0.i11047_3_lut_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11047_3_lut_LC_7_2_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.i11047_3_lut_LC_7_2_1  (
            .in0(N__48998),
            .in1(N__47960),
            .in2(_gnd_net_),
            .in3(N__48923),
            .lcout(),
            .ltout(\c0.n13808_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_439_LC_7_2_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_439_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_439_LC_7_2_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_439_LC_7_2_2  (
            .in0(N__25218),
            .in1(N__25299),
            .in2(N__25149),
            .in3(N__25260),
            .lcout(\c0.n14064 ),
            .ltout(\c0.n14064_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_2_lut_3_lut_LC_7_2_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_2_lut_3_lut_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_2_lut_3_lut_LC_7_2_3 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \c0.i1_2_lut_2_lut_3_lut_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__29928),
            .in2(N__25146),
            .in3(N__30191),
            .lcout(n612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i5_LC_7_2_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i5_LC_7_2_4 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i5_LC_7_2_4 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i5_LC_7_2_4  (
            .in0(N__25281),
            .in1(N__25300),
            .in2(N__30650),
            .in3(N__30551),
            .lcout(\c0.byte_transmit_counter2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49843),
            .ce(),
            .sr(N__25143));
    defparam \c0.i1_2_lut_4_lut_adj_773_LC_7_2_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_773_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_773_LC_7_2_5 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_773_LC_7_2_5  (
            .in0(N__33088),
            .in1(N__25269),
            .in2(N__25074),
            .in3(N__25124),
            .lcout(\c0.n4_adj_2201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_774_LC_7_2_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_774_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_774_LC_7_2_6 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_774_LC_7_2_6  (
            .in0(N__25125),
            .in1(N__25073),
            .in2(N__25226),
            .in3(N__33089),
            .lcout(\c0.n4_adj_2199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11300_1_lut_LC_7_2_7 .C_ON=1'b0;
    defparam \c0.i11300_1_lut_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11300_1_lut_LC_7_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.i11300_1_lut_LC_7_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30149),
            .lcout(\c0.tx2_transmit_N_1996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_2_lut_LC_7_3_0 .C_ON=1'b1;
    defparam \c0.add_2510_2_lut_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_2_lut_LC_7_3_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_2_lut_LC_7_3_0  (
            .in0(N__25196),
            .in1(N__46160),
            .in2(_gnd_net_),
            .in3(N__25014),
            .lcout(\c0.n18254 ),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(\c0.n16479 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_3_lut_LC_7_3_1 .C_ON=1'b1;
    defparam \c0.add_2510_3_lut_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_3_lut_LC_7_3_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_3_lut_LC_7_3_1  (
            .in0(N__25182),
            .in1(N__48622),
            .in2(_gnd_net_),
            .in3(N__24996),
            .lcout(\c0.n18253 ),
            .ltout(),
            .carryin(\c0.n16479 ),
            .carryout(\c0.n16480 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_4_lut_LC_7_3_2 .C_ON=1'b1;
    defparam \c0.add_2510_4_lut_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_4_lut_LC_7_3_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_4_lut_LC_7_3_2  (
            .in0(N__25200),
            .in1(N__47977),
            .in2(_gnd_net_),
            .in3(N__24987),
            .lcout(\c0.n18314 ),
            .ltout(),
            .carryin(\c0.n16480 ),
            .carryout(\c0.n16481 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_5_lut_LC_7_3_3 .C_ON=1'b1;
    defparam \c0.add_2510_5_lut_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_5_lut_LC_7_3_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_5_lut_LC_7_3_3  (
            .in0(N__25184),
            .in1(N__48986),
            .in2(_gnd_net_),
            .in3(N__25311),
            .lcout(\c0.n18315 ),
            .ltout(),
            .carryin(\c0.n16481 ),
            .carryout(\c0.n16482 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_6_lut_LC_7_3_4 .C_ON=1'b1;
    defparam \c0.add_2510_6_lut_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_6_lut_LC_7_3_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_6_lut_LC_7_3_4  (
            .in0(N__25197),
            .in1(N__48925),
            .in2(_gnd_net_),
            .in3(N__25308),
            .lcout(\c0.n18362 ),
            .ltout(),
            .carryin(\c0.n16482 ),
            .carryout(\c0.n16483 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_7_lut_LC_7_3_5 .C_ON=1'b1;
    defparam \c0.add_2510_7_lut_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_7_lut_LC_7_3_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_7_lut_LC_7_3_5  (
            .in0(N__25183),
            .in1(N__25301),
            .in2(_gnd_net_),
            .in3(N__25272),
            .lcout(\c0.n18316 ),
            .ltout(),
            .carryin(\c0.n16483 ),
            .carryout(\c0.n16484 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_8_lut_LC_7_3_6 .C_ON=1'b1;
    defparam \c0.add_2510_8_lut_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_8_lut_LC_7_3_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_8_lut_LC_7_3_6  (
            .in0(N__25199),
            .in1(N__25268),
            .in2(_gnd_net_),
            .in3(N__25230),
            .lcout(\c0.n18317 ),
            .ltout(),
            .carryin(\c0.n16484 ),
            .carryout(\c0.n16485 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_9_lut_LC_7_3_7 .C_ON=1'b0;
    defparam \c0.add_2510_9_lut_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_9_lut_LC_7_3_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.add_2510_9_lut_LC_7_3_7  (
            .in0(N__25227),
            .in1(N__25198),
            .in2(_gnd_net_),
            .in3(N__25167),
            .lcout(\c0.n18318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15239_4_lut_LC_7_4_0 .C_ON=1'b0;
    defparam \c0.i15239_4_lut_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15239_4_lut_LC_7_4_0 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i15239_4_lut_LC_7_4_0  (
            .in0(N__28892),
            .in1(N__28815),
            .in2(N__40462),
            .in3(N__28868),
            .lcout(),
            .ltout(\c0.n18100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i2_LC_7_4_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i2_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i2_LC_7_4_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i2_LC_7_4_1  (
            .in0(N__28818),
            .in1(N__28989),
            .in2(N__25155),
            .in3(N__28920),
            .lcout(\c0.data_out_frame2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15242_4_lut_LC_7_4_2 .C_ON=1'b0;
    defparam \c0.i15242_4_lut_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15242_4_lut_LC_7_4_2 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i15242_4_lut_LC_7_4_2  (
            .in0(N__28893),
            .in1(N__28816),
            .in2(N__41613),
            .in3(N__28869),
            .lcout(),
            .ltout(\c0.n18103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i1_LC_7_4_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i1_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i1_LC_7_4_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i1_LC_7_4_3  (
            .in0(N__28817),
            .in1(N__28988),
            .in2(N__25152),
            .in3(N__28919),
            .lcout(\c0.data_out_frame2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_665_LC_7_4_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_665_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_665_LC_7_4_4 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \c0.i11_4_lut_adj_665_LC_7_4_4  (
            .in0(N__25442),
            .in1(N__26205),
            .in2(N__25415),
            .in3(N__25398),
            .lcout(\c0.n27_adj_2405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_7_4_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_7_4_5 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_in_frame_0__i27_LC_7_4_5  (
            .in0(N__25391),
            .in1(N__25700),
            .in2(N__26726),
            .in3(N__25557),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11390_2_lut_LC_7_4_6 .C_ON=1'b0;
    defparam \c0.i11390_2_lut_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11390_2_lut_LC_7_4_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i11390_2_lut_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(N__30070),
            .in2(_gnd_net_),
            .in3(N__30132),
            .lcout(\c0.n14161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_7_4_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_7_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i55_LC_7_4_7  (
            .in0(N__27622),
            .in1(N__25370),
            .in2(_gnd_net_),
            .in3(N__25862),
            .lcout(data_in_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_403_LC_7_5_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_403_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_403_LC_7_5_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_4_lut_adj_403_LC_7_5_0  (
            .in0(N__27435),
            .in1(N__27549),
            .in2(N__28155),
            .in3(N__27944),
            .lcout(n158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_633_LC_7_5_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_633_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_633_LC_7_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_633_LC_7_5_1  (
            .in0(N__25356),
            .in1(N__26012),
            .in2(_gnd_net_),
            .in3(N__26069),
            .lcout(\c0.n16982 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_7_5_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_7_5_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_in_frame_0__i29_LC_7_5_2  (
            .in0(N__26111),
            .in1(N__25552),
            .in2(N__26494),
            .in3(N__25677),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_416_LC_7_5_3 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_416_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_416_LC_7_5_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_416_LC_7_5_3  (
            .in0(N__27943),
            .in1(N__28150),
            .in2(_gnd_net_),
            .in3(N__27434),
            .lcout(n135_adj_2463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_7_5_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_7_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i51_LC_7_5_4  (
            .in0(N__26718),
            .in1(N__25331),
            .in2(_gnd_net_),
            .in3(N__25865),
            .lcout(data_in_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_7_5_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_7_5_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_in_frame_0__i31_LC_7_5_5  (
            .in0(N__25553),
            .in1(N__27623),
            .in2(N__25704),
            .in3(N__26093),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_7_5_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_7_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i53_LC_7_5_6  (
            .in0(N__26475),
            .in1(N__26240),
            .in2(_gnd_net_),
            .in3(N__25866),
            .lcout(data_in_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_635_LC_7_5_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_635_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_635_LC_7_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_635_LC_7_5_7  (
            .in0(N__25830),
            .in1(N__25476),
            .in2(_gnd_net_),
            .in3(N__26298),
            .lcout(\c0.n17725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_7_6_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_7_6_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_7_6_0  (
            .in0(N__30372),
            .in1(N__30783),
            .in2(N__30416),
            .in3(N__29850),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_6_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_6_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_7_6_1  (
            .in0(N__25812),
            .in1(N__28020),
            .in2(N__25781),
            .in3(N__25806),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_7_6_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_7_6_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i9_LC_7_6_2  (
            .in0(N__25702),
            .in1(N__25556),
            .in2(N__26646),
            .in3(N__26070),
            .lcout(\c0.data_in_frame_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_7_6_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_7_6_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i13_LC_7_6_3  (
            .in0(N__25555),
            .in1(N__25703),
            .in2(N__26505),
            .in3(N__25945),
            .lcout(\c0.data_in_frame_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_7_6_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_7_6_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_7_6_4  (
            .in0(N__25701),
            .in1(N__25554),
            .in2(N__27135),
            .in3(N__26038),
            .lcout(\c0.data_in_frame_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_631_LC_7_6_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_631_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_631_LC_7_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_631_LC_7_6_6  (
            .in0(N__25494),
            .in1(N__25475),
            .in2(_gnd_net_),
            .in3(N__26037),
            .lcout(),
            .ltout(\c0.n16981_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_652_LC_7_6_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_652_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_652_LC_7_6_7 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i4_4_lut_adj_652_LC_7_6_7  (
            .in0(N__26322),
            .in1(N__26302),
            .in2(N__26271),
            .in3(N__25944),
            .lcout(\c0.n20_adj_2397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_516_LC_7_7_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_516_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_516_LC_7_7_0 .LUT_INIT=16'b1001111111111001;
    LogicCell40 \c0.i4_4_lut_adj_516_LC_7_7_0  (
            .in0(N__26067),
            .in1(N__26247),
            .in2(N__26393),
            .in3(N__26142),
            .lcout(\c0.n20_adj_2350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1016_2_lut_LC_7_7_1 .C_ON=1'b0;
    defparam \c0.i1016_2_lut_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1016_2_lut_LC_7_7_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1016_2_lut_LC_7_7_1  (
            .in0(N__25901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26004),
            .lcout(\c0.n2128 ),
            .ltout(\c0.n2128_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_643_LC_7_7_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_643_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_643_LC_7_7_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i6_4_lut_adj_643_LC_7_7_2  (
            .in0(N__26241),
            .in1(N__26226),
            .in2(N__26208),
            .in3(N__26141),
            .lcout(\c0.n22_adj_2392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1008_2_lut_LC_7_7_3 .C_ON=1'b0;
    defparam \c0.i1008_2_lut_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1008_2_lut_LC_7_7_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1008_2_lut_LC_7_7_3  (
            .in0(N__26192),
            .in1(_gnd_net_),
            .in2(N__26174),
            .in3(_gnd_net_),
            .lcout(\c0.n2120 ),
            .ltout(\c0.n2120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_690_LC_7_7_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_690_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_690_LC_7_7_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i5_4_lut_adj_690_LC_7_7_4  (
            .in0(N__26131),
            .in1(N__26112),
            .in2(N__26097),
            .in3(N__26094),
            .lcout(\c0.n19_adj_2415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_624_LC_7_7_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_624_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_624_LC_7_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_624_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__26066),
            .in2(_gnd_net_),
            .in3(N__26036),
            .lcout(),
            .ltout(\c0.n17721_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_626_LC_7_7_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_626_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_626_LC_7_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_626_LC_7_7_6  (
            .in0(N__26003),
            .in1(N__25940),
            .in2(N__25917),
            .in3(N__25900),
            .lcout(\c0.n10_adj_2390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_7_7_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_7_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i21_LC_7_7_7  (
            .in0(N__26500),
            .in1(N__26389),
            .in2(_gnd_net_),
            .in3(N__26424),
            .lcout(data_in_frame_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_8_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_8_0 .LUT_INIT=16'b0111101000101010;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_8_0  (
            .in0(N__27926),
            .in1(N__26956),
            .in2(N__28136),
            .in3(N__26354),
            .lcout(),
            .ltout(\c0.rx.n18729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.n18729_bdd_4_lut_4_lut_LC_7_8_1 .C_ON=1'b0;
    defparam \c0.rx.n18729_bdd_4_lut_4_lut_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n18729_bdd_4_lut_4_lut_LC_7_8_1 .LUT_INIT=16'b1110000011100101;
    LogicCell40 \c0.rx.n18729_bdd_4_lut_4_lut_LC_7_8_1  (
            .in0(N__28149),
            .in1(N__28287),
            .in2(N__26373),
            .in3(N__28005),
            .lcout(),
            .ltout(\c0.rx.n18732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_7_8_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_7_8_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26370),
            .in3(N__27428),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_7_8_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.rx.i3_4_lut_LC_7_8_3  (
            .in0(N__27542),
            .in1(N__28107),
            .in2(N__27807),
            .in3(N__26660),
            .lcout(\c0.rx.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_7_8_4 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_7_8_4 .LUT_INIT=16'b1001100011001000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_7_8_4  (
            .in0(N__27797),
            .in1(N__26864),
            .in2(N__28137),
            .in3(N__26957),
            .lcout(\c0.rx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_409_LC_7_8_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_409_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_409_LC_7_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_409_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__27541),
            .in2(_gnd_net_),
            .in3(N__26659),
            .lcout(n12582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_418_LC_7_8_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_418_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_418_LC_7_8_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_418_LC_7_8_6  (
            .in0(N__26339),
            .in1(N__27543),
            .in2(_gnd_net_),
            .in3(N__27856),
            .lcout(),
            .ltout(n4_adj_2471_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_8_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_8_7 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_7_8_7  (
            .in0(N__26689),
            .in1(N__28006),
            .in2(N__26325),
            .in3(N__27753),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__0__2285_LC_7_9_0 .C_ON=1'b0;
    defparam \c0.data_in_1__0__2285_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0__2285_LC_7_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_1__0__2285_LC_7_9_0  (
            .in0(N__27039),
            .in1(N__26750),
            .in2(_gnd_net_),
            .in3(N__34195),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_9_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_LC_7_9_1  (
            .in0(N__27846),
            .in1(N__27809),
            .in2(N__27548),
            .in3(N__27748),
            .lcout(\c0.rx.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2__2267_LC_7_9_2 .C_ON=1'b0;
    defparam \c0.data_in_3__2__2267_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2__2267_LC_7_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__2__2267_LC_7_9_2  (
            .in0(N__26705),
            .in1(N__34194),
            .in2(_gnd_net_),
            .in3(N__26572),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_420_LC_7_9_3 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_420_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_420_LC_7_9_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.rx.i1_4_lut_adj_420_LC_7_9_3  (
            .in0(N__28200),
            .in1(N__29143),
            .in2(N__28260),
            .in3(N__28223),
            .lcout(\c0.rx.r_SM_Main_2_N_2088_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2088_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_411_LC_7_9_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_411_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_411_LC_7_9_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_411_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__27845),
            .in2(N__26664),
            .in3(N__26851),
            .lcout(\c0.rx.n161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0__2269_LC_7_9_5 .C_ON=1'b0;
    defparam \c0.data_in_3__0__2269_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0__2269_LC_7_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__0__2269_LC_7_9_5  (
            .in0(N__34193),
            .in1(N__26637),
            .in2(_gnd_net_),
            .in3(N__27062),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2__2275_LC_7_9_6 .C_ON=1'b0;
    defparam \c0.data_in_2__2__2275_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2__2275_LC_7_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__2__2275_LC_7_9_6  (
            .in0(N__26807),
            .in1(N__26573),
            .in2(_gnd_net_),
            .in3(N__34196),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__6__2287_LC_7_9_7 .C_ON=1'b0;
    defparam \c0.data_in_0__6__2287_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6__2287_LC_7_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__6__2287_LC_7_9_7  (
            .in0(N__34192),
            .in1(N__26549),
            .in2(_gnd_net_),
            .in3(N__27258),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6__2271_LC_7_10_0 .C_ON=1'b0;
    defparam \c0.data_in_2__6__2271_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6__2271_LC_7_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__6__2271_LC_7_10_0  (
            .in0(N__27276),
            .in1(N__26527),
            .in2(_gnd_net_),
            .in3(N__34219),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49749),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_613_LC_7_10_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_613_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_613_LC_7_10_1 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.i3_4_lut_adj_613_LC_7_10_1  (
            .in0(N__29279),
            .in1(N__26903),
            .in2(N__26529),
            .in3(N__26768),
            .lcout(\c0.n8_adj_2385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_573_LC_7_10_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_573_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_573_LC_7_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i4_2_lut_adj_573_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__27274),
            .lcout(\c0.n15_adj_2372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2__2283_LC_7_10_3 .C_ON=1'b0;
    defparam \c0.data_in_1__2__2283_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2__2283_LC_7_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__2__2283_LC_7_10_3  (
            .in0(N__34218),
            .in1(N__26904),
            .in2(_gnd_net_),
            .in3(N__26802),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49749),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_422_LC_7_10_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_422_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_422_LC_7_10_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_422_LC_7_10_4  (
            .in0(N__26865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26954),
            .lcout(n12527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7__2286_LC_7_10_5 .C_ON=1'b0;
    defparam \c0.data_in_0__7__2286_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7__2286_LC_7_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__7__2286_LC_7_10_5  (
            .in0(N__34217),
            .in1(N__27009),
            .in2(_gnd_net_),
            .in3(N__26885),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49749),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_417_LC_7_10_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_417_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_417_LC_7_10_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_417_LC_7_10_6  (
            .in0(N__26866),
            .in1(_gnd_net_),
            .in2(N__27857),
            .in3(N__26955),
            .lcout(n151),
            .ltout(n151_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15541_3_lut_LC_7_10_7 .C_ON=1'b0;
    defparam \c0.rx.i15541_3_lut_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15541_3_lut_LC_7_10_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.rx.i15541_3_lut_LC_7_10_7  (
            .in0(N__27529),
            .in1(_gnd_net_),
            .in2(N__26811),
            .in3(N__27808),
            .lcout(\c0.rx.n18194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_563_LC_7_11_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_563_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_563_LC_7_11_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i3_4_lut_adj_563_LC_7_11_1  (
            .in0(N__26803),
            .in1(N__26778),
            .in2(N__27035),
            .in3(N__27696),
            .lcout(),
            .ltout(\c0.n8_adj_2369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_565_LC_7_11_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_565_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_565_LC_7_11_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i1_4_lut_adj_565_LC_7_11_2  (
            .in0(N__27150),
            .in1(N__26982),
            .in2(N__26772),
            .in3(N__27252),
            .lcout(\c0.n10493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6__2279_LC_7_11_3 .C_ON=1'b0;
    defparam \c0.data_in_1__6__2279_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6__2279_LC_7_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_1__6__2279_LC_7_11_3  (
            .in0(N__27253),
            .in1(N__27275),
            .in2(_gnd_net_),
            .in3(N__34211),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_7_11_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_7_11_4 .LUT_INIT=16'b0001000000010101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_7_11_4  (
            .in0(N__27455),
            .in1(N__27234),
            .in2(N__28118),
            .in3(N__28269),
            .lcout(\c0.rx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5__2264_LC_7_11_5 .C_ON=1'b0;
    defparam \c0.data_in_3__5__2264_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5__2264_LC_7_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__5__2264_LC_7_11_5  (
            .in0(N__27219),
            .in1(N__34210),
            .in2(_gnd_net_),
            .in3(N__27151),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1__2268_LC_7_11_6 .C_ON=1'b0;
    defparam \c0.data_in_3__1__2268_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1__2268_LC_7_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__1__2268_LC_7_11_6  (
            .in0(N__34208),
            .in1(N__27134),
            .in2(_gnd_net_),
            .in3(N__34301),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0__2277_LC_7_11_7 .C_ON=1'b0;
    defparam \c0.data_in_2__0__2277_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0__2277_LC_7_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_2__0__2277_LC_7_11_7  (
            .in0(N__27030),
            .in1(N__34209),
            .in2(_gnd_net_),
            .in3(N__27066),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_3_lut_4_lut_LC_7_12_0 .C_ON=1'b0;
    defparam \c0.rx.i3_3_lut_4_lut_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_3_lut_4_lut_LC_7_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i3_3_lut_4_lut_LC_7_12_0  (
            .in0(N__27352),
            .in1(N__27334),
            .in2(N__27318),
            .in3(N__27292),
            .lcout(\c0.rx.n15902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10932_2_lut_LC_7_12_1 .C_ON=1'b0;
    defparam \c0.i10932_2_lut_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10932_2_lut_LC_7_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10932_2_lut_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__27000),
            .in2(_gnd_net_),
            .in3(N__27673),
            .lcout(\c0.n13693 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_3_lut_4_lut_4_lut_LC_7_12_2 .C_ON=1'b0;
    defparam \c0.rx.i13_3_lut_4_lut_4_lut_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_3_lut_4_lut_4_lut_LC_7_12_2 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \c0.rx.i13_3_lut_4_lut_4_lut_LC_7_12_2  (
            .in0(N__27948),
            .in1(N__27450),
            .in2(N__28138),
            .in3(N__26974),
            .lcout(),
            .ltout(\c0.rx.n11041_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_7_12_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_7_12_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_7_12_3  (
            .in0(N__27451),
            .in1(N__34188),
            .in2(N__26922),
            .in3(N__28117),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15577_3_lut_4_lut_LC_7_12_4 .C_ON=1'b0;
    defparam \c0.rx.i15577_3_lut_4_lut_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15577_3_lut_4_lut_LC_7_12_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.rx.i15577_3_lut_4_lut_LC_7_12_4  (
            .in0(N__27858),
            .in1(N__27810),
            .in2(N__27547),
            .in3(N__27752),
            .lcout(\c0.rx.n18196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_559_LC_7_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_559_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_559_LC_7_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_559_LC_7_12_5  (
            .in0(N__27727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27711),
            .lcout(\c0.n6_adj_2368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3__2290_LC_7_12_6 .C_ON=1'b0;
    defparam \c0.data_in_0__3__2290_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3__2290_LC_7_12_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0__3__2290_LC_7_12_6  (
            .in0(N__27674),
            .in1(N__34180),
            .in2(_gnd_net_),
            .in3(N__27690),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1__2292_LC_7_12_7 .C_ON=1'b0;
    defparam \c0.data_in_0__1__2292_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1__2292_LC_7_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__1__2292_LC_7_12_7  (
            .in0(N__34179),
            .in1(N__29283),
            .in2(_gnd_net_),
            .in3(N__27660),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i9777_4_lut_LC_7_13_0 .C_ON=1'b0;
    defparam \c0.rx.i9777_4_lut_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i9777_4_lut_LC_7_13_0 .LUT_INIT=16'b1110110011100000;
    LogicCell40 \c0.rx.i9777_4_lut_LC_7_13_0  (
            .in0(N__27645),
            .in1(N__28023),
            .in2(N__27586),
            .in3(N__27639),
            .lcout(),
            .ltout(\c0.rx.n12552_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_13_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_13_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__27572),
            .in2(N__27630),
            .in3(N__28123),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49714),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_404_LC_7_13_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_404_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_4_lut_adj_404_LC_7_13_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_4_lut_adj_404_LC_7_13_2  (
            .in0(N__27510),
            .in1(N__27456),
            .in2(N__28139),
            .in3(N__27947),
            .lcout(n164_adj_2464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15131_2_lut_LC_7_13_3 .C_ON=1'b0;
    defparam \c0.rx.i15131_2_lut_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15131_2_lut_LC_7_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i15131_2_lut_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__27353),
            .in2(_gnd_net_),
            .in3(N__27335),
            .lcout(),
            .ltout(\c0.rx.n17990_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15163_4_lut_LC_7_13_4 .C_ON=1'b0;
    defparam \c0.rx.i15163_4_lut_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15163_4_lut_LC_7_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i15163_4_lut_LC_7_13_4  (
            .in0(N__28197),
            .in1(N__27316),
            .in2(N__27297),
            .in3(N__27293),
            .lcout(),
            .ltout(\c0.rx.n18024_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_7_13_5 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_7_13_5 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \c0.rx.i2_3_lut_LC_7_13_5  (
            .in0(N__28252),
            .in1(_gnd_net_),
            .in2(N__28290),
            .in3(N__29150),
            .lcout(\c0.rx.n12828 ),
            .ltout(\c0.rx.n12828_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15639_3_lut_LC_7_13_6 .C_ON=1'b0;
    defparam \c0.rx.i15639_3_lut_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15639_3_lut_LC_7_13_6 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \c0.rx.i15639_3_lut_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__28022),
            .in2(N__28272),
            .in3(N__27946),
            .lcout(\c0.rx.n18303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15551_2_lut_3_lut_LC_7_13_7 .C_ON=1'b0;
    defparam \c0.rx.i15551_2_lut_3_lut_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15551_2_lut_3_lut_LC_7_13_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i15551_2_lut_3_lut_LC_7_13_7  (
            .in0(N__28251),
            .in1(N__28222),
            .in2(_gnd_net_),
            .in3(N__28198),
            .lcout(\c0.rx.n18211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_adj_419_LC_7_14_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_adj_419_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_adj_419_LC_7_14_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_adj_419_LC_7_14_0  (
            .in0(N__28086),
            .in1(N__28021),
            .in2(_gnd_net_),
            .in3(N__27945),
            .lcout(\c0.rx.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_LC_7_14_3 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_LC_7_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i4_4_lut_LC_7_14_3  (
            .in0(N__28334),
            .in1(N__28349),
            .in2(N__28386),
            .in3(N__28400),
            .lcout(\c0.tx.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_LC_7_14_4 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_LC_7_14_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.tx.i2_3_lut_LC_7_14_4  (
            .in0(N__28494),
            .in1(N__28304),
            .in2(_gnd_net_),
            .in3(N__28319),
            .lcout(\c0.tx.n54 ),
            .ltout(\c0.tx.n54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i11043_2_lut_4_lut_LC_7_14_5 .C_ON=1'b0;
    defparam \c0.tx.i11043_2_lut_4_lut_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i11043_2_lut_4_lut_LC_7_14_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.tx.i11043_2_lut_4_lut_LC_7_14_5  (
            .in0(N__28366),
            .in1(N__28417),
            .in2(N__27870),
            .in3(N__27866),
            .lcout(\c0.tx.r_SM_Main_2_N_2031_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5_3_lut_LC_7_14_6 .C_ON=1'b0;
    defparam \c0.tx.i5_3_lut_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5_3_lut_LC_7_14_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.tx.i5_3_lut_LC_7_14_6  (
            .in0(N__27867),
            .in1(_gnd_net_),
            .in2(N__28422),
            .in3(N__28367),
            .lcout(),
            .ltout(\c0.tx.n47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_7_14_7 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_7_14_7 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \c0.tx.i1_4_lut_LC_7_14_7  (
            .in0(N__29400),
            .in1(N__28431),
            .in2(N__28425),
            .in3(N__29472),
            .lcout(\c0.tx.n11297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_7_15_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i0_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_7_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__28421),
            .in2(_gnd_net_),
            .in3(N__28404),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\c0.tx.n16524 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i1_LC_7_15_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i1_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_7_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__28401),
            .in2(_gnd_net_),
            .in3(N__28389),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx.n16524 ),
            .carryout(\c0.tx.n16525 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i2_LC_7_15_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i2_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_7_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__28385),
            .in2(_gnd_net_),
            .in3(N__28371),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx.n16525 ),
            .carryout(\c0.tx.n16526 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i3_LC_7_15_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i3_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_7_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__28368),
            .in2(_gnd_net_),
            .in3(N__28353),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx.n16526 ),
            .carryout(\c0.tx.n16527 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i4_LC_7_15_4 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i4_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_7_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__28350),
            .in2(_gnd_net_),
            .in3(N__28338),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx.n16527 ),
            .carryout(\c0.tx.n16528 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i5_LC_7_15_5 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i5_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_7_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__28335),
            .in2(_gnd_net_),
            .in3(N__28323),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx.n16528 ),
            .carryout(\c0.tx.n16529 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i6_LC_7_15_6 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i6_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_7_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__28320),
            .in2(_gnd_net_),
            .in3(N__28308),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx.n16529 ),
            .carryout(\c0.tx.n16530 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i7_LC_7_15_7 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i7_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_7_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__28305),
            .in2(_gnd_net_),
            .in3(N__28293),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx.n16530 ),
            .carryout(\c0.tx.n16531 ),
            .clk(N__49696),
            .ce(N__29484),
            .sr(N__28475));
    defparam \c0.tx.r_Clock_Count__i8_LC_7_16_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_7_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__28493),
            .in2(_gnd_net_),
            .in3(N__28497),
            .lcout(\c0.tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(N__29483),
            .sr(N__28479));
    defparam \control.i15748_2_lut_3_lut_LC_7_27_4 .C_ON=1'b0;
    defparam \control.i15748_2_lut_3_lut_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \control.i15748_2_lut_3_lut_LC_7_27_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \control.i15748_2_lut_3_lut_LC_7_27_4  (
            .in0(N__28460),
            .in1(N__32906),
            .in2(_gnd_net_),
            .in3(N__32858),
            .lcout(\control.n6_adj_2460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i19_3_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \control.i19_3_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \control.i19_3_lut_LC_7_28_4 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \control.i19_3_lut_LC_7_28_4  (
            .in0(N__35663),
            .in1(N__35444),
            .in2(_gnd_net_),
            .in3(N__35512),
            .lcout(\control.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i5146_2_lut_LC_7_29_3 .C_ON=1'b0;
    defparam \control.i5146_2_lut_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \control.i5146_2_lut_LC_7_29_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \control.i5146_2_lut_LC_7_29_3  (
            .in0(N__35443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35664),
            .lcout(\control.PHASES_5_N_2152_1 ),
            .ltout(\control.PHASES_5_N_2152_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i1_2_lut_4_lut_LC_7_29_4 .C_ON=1'b0;
    defparam \control.i1_2_lut_4_lut_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \control.i1_2_lut_4_lut_LC_7_29_4 .LUT_INIT=16'b1111111101110010;
    LogicCell40 \control.i1_2_lut_4_lut_LC_7_29_4  (
            .in0(N__35559),
            .in1(N__35442),
            .in2(N__28449),
            .in3(N__35337),
            .lcout(\control.n10356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_9_1_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_9_1_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_9_1_0  (
            .in0(N__48032),
            .in1(N__48171),
            .in2(N__45336),
            .in3(N__28437),
            .lcout(\c0.n22_adj_2239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15978_LC_9_1_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15978_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15978_LC_9_1_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15978_LC_9_1_1  (
            .in0(N__28575),
            .in1(N__49045),
            .in2(N__40602),
            .in3(N__48031),
            .lcout(\c0.n18843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15914_LC_9_1_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15914_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15914_LC_9_1_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15914_LC_9_1_2  (
            .in0(N__31761),
            .in1(N__48604),
            .in2(N__46212),
            .in3(N__37872),
            .lcout(),
            .ltout(\c0.n18801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18801_bdd_4_lut_LC_9_1_3 .C_ON=1'b0;
    defparam \c0.n18801_bdd_4_lut_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18801_bdd_4_lut_LC_9_1_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18801_bdd_4_lut_LC_9_1_3  (
            .in0(N__48605),
            .in1(N__31809),
            .in2(N__28440),
            .in3(N__40991),
            .lcout(\c0.n18804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18843_bdd_4_lut_LC_9_1_4 .C_ON=1'b0;
    defparam \c0.n18843_bdd_4_lut_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18843_bdd_4_lut_LC_9_1_4 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n18843_bdd_4_lut_LC_9_1_4  (
            .in0(N__49046),
            .in1(N__31644),
            .in2(N__29799),
            .in3(N__28563),
            .lcout(),
            .ltout(\c0.n18846_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_9_1_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_9_1_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_9_1_5  (
            .in0(N__48926),
            .in1(N__49047),
            .in2(N__28557),
            .in3(N__28554),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49866),
            .ce(N__48796),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15814_LC_9_2_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15814_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15814_LC_9_2_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15814_LC_9_2_0  (
            .in0(N__33999),
            .in1(N__48482),
            .in2(N__36087),
            .in3(N__46017),
            .lcout(),
            .ltout(\c0.n18675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18675_bdd_4_lut_LC_9_2_1 .C_ON=1'b0;
    defparam \c0.n18675_bdd_4_lut_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18675_bdd_4_lut_LC_9_2_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18675_bdd_4_lut_LC_9_2_1  (
            .in0(N__48483),
            .in1(N__32991),
            .in2(N__28530),
            .in3(N__45454),
            .lcout(),
            .ltout(\c0.n18678_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_9_2_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_9_2_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_9_2_2  (
            .in0(N__48029),
            .in1(N__35877),
            .in2(N__28527),
            .in3(N__48168),
            .lcout(\c0.n22_adj_2242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15879_LC_9_2_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15879_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15879_LC_9_2_3 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15879_LC_9_2_3  (
            .in0(N__28581),
            .in1(N__49048),
            .in2(N__29784),
            .in3(N__48030),
            .lcout(),
            .ltout(\c0.n18741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18741_bdd_4_lut_LC_9_2_4 .C_ON=1'b0;
    defparam \c0.n18741_bdd_4_lut_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18741_bdd_4_lut_LC_9_2_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18741_bdd_4_lut_LC_9_2_4  (
            .in0(N__49049),
            .in1(N__29742),
            .in2(N__28524),
            .in3(N__31743),
            .lcout(),
            .ltout(\c0.n18744_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_9_2_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_9_2_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_9_2_5  (
            .in0(N__28521),
            .in1(N__49050),
            .in2(N__28515),
            .in3(N__48924),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49859),
            .ce(N__48786),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i4_LC_9_3_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i4_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i4_LC_9_3_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.data_out_frame2_0___i4_LC_9_3_0  (
            .in0(N__28987),
            .in1(N__28656),
            .in2(N__45092),
            .in3(N__28719),
            .lcout(\c0.data_out_frame2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15710_4_lut_4_lut_LC_9_3_1 .C_ON=1'b0;
    defparam \c0.tx2.i15710_4_lut_4_lut_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15710_4_lut_4_lut_LC_9_3_1 .LUT_INIT=16'b1000001110000000;
    LogicCell40 \c0.tx2.i15710_4_lut_4_lut_LC_9_3_1  (
            .in0(N__29841),
            .in1(N__30340),
            .in2(N__30441),
            .in3(N__29926),
            .lcout(),
            .ltout(n17689_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_9_3_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_9_3_2 .LUT_INIT=16'b1000101010111010;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_9_3_2  (
            .in0(N__30184),
            .in1(N__30762),
            .in2(N__28584),
            .in3(N__30435),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18681_bdd_4_lut_LC_9_3_3 .C_ON=1'b0;
    defparam \c0.n18681_bdd_4_lut_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18681_bdd_4_lut_LC_9_3_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18681_bdd_4_lut_LC_9_3_3  (
            .in0(N__48481),
            .in1(N__44806),
            .in2(N__44171),
            .in3(N__37929),
            .lcout(\c0.n18684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_9_3_4 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_9_3_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_9_3_4  (
            .in0(N__29925),
            .in1(N__30434),
            .in2(N__30355),
            .in3(N__30761),
            .lcout(\c0.tx2.n9639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18855_bdd_4_lut_LC_9_3_5 .C_ON=1'b0;
    defparam \c0.n18855_bdd_4_lut_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18855_bdd_4_lut_LC_9_3_5 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18855_bdd_4_lut_LC_9_3_5  (
            .in0(N__48480),
            .in1(N__29733),
            .in2(N__41678),
            .in3(N__41154),
            .lcout(\c0.n18072 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i34_2_lut_LC_9_3_6 .C_ON=1'b0;
    defparam \c0.tx2.i34_2_lut_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i34_2_lut_LC_9_3_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.tx2.i34_2_lut_LC_9_3_6  (
            .in0(N__30339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30430),
            .lcout(),
            .ltout(\c0.tx2.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_4_lut_LC_9_3_7 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_4_lut_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_4_lut_LC_9_3_7 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \c0.tx2.i1_4_lut_4_lut_LC_9_3_7  (
            .in0(N__29876),
            .in1(N__30781),
            .in2(N__28566),
            .in3(N__30810),
            .lcout(\c0.tx2.n11312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_630_LC_9_4_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_630_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_630_LC_9_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_630_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__30067),
            .in2(_gnd_net_),
            .in3(N__28696),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15633_3_lut_4_lut_LC_9_4_1 .C_ON=1'b0;
    defparam \c0.i15633_3_lut_4_lut_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15633_3_lut_4_lut_LC_9_4_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \c0.i15633_3_lut_4_lut_LC_9_4_1  (
            .in0(N__28698),
            .in1(N__30071),
            .in2(N__37741),
            .in3(N__28861),
            .lcout(),
            .ltout(\c0.n18284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i5_LC_9_4_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i5_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i5_LC_9_4_2 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.data_out_frame2_0___i5_LC_9_4_2  (
            .in0(N__37721),
            .in1(N__28984),
            .in2(N__28746),
            .in3(N__28655),
            .lcout(\c0.data_out_frame2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_680_LC_9_4_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_680_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_680_LC_9_4_3 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \c0.i1_4_lut_adj_680_LC_9_4_3  (
            .in0(N__30068),
            .in1(N__28743),
            .in2(N__28593),
            .in3(N__28734),
            .lcout(\c0.n12704 ),
            .ltout(\c0.n12704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15621_3_lut_4_lut_LC_9_4_4 .C_ON=1'b0;
    defparam \c0.i15621_3_lut_4_lut_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15621_3_lut_4_lut_LC_9_4_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.i15621_3_lut_4_lut_LC_9_4_4  (
            .in0(N__45077),
            .in1(N__30069),
            .in2(N__28722),
            .in3(N__28697),
            .lcout(\c0.n18287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15636_3_lut_4_lut_LC_9_4_5 .C_ON=1'b0;
    defparam \c0.i15636_3_lut_4_lut_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15636_3_lut_4_lut_LC_9_4_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \c0.i15636_3_lut_4_lut_LC_9_4_5  (
            .in0(N__28699),
            .in1(N__30072),
            .in2(N__50664),
            .in3(N__28862),
            .lcout(),
            .ltout(\c0.n18289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i3_LC_9_4_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i3_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i3_LC_9_4_6 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.data_out_frame2_0___i3_LC_9_4_6  (
            .in0(N__50655),
            .in1(N__28983),
            .in2(N__28659),
            .in3(N__28654),
            .lcout(\c0.data_out_frame2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6035_bdd_4_lut_4_lut_LC_9_4_7 .C_ON=1'b0;
    defparam \c0.n6035_bdd_4_lut_4_lut_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6035_bdd_4_lut_4_lut_LC_9_4_7 .LUT_INIT=16'b0101100011111000;
    LogicCell40 \c0.n6035_bdd_4_lut_4_lut_LC_9_4_7  (
            .in0(N__28982),
            .in1(N__28924),
            .in2(N__28804),
            .in3(N__33083),
            .lcout(\c0.n18831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15218_4_lut_LC_9_5_0 .C_ON=1'b0;
    defparam \c0.i15218_4_lut_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15218_4_lut_LC_9_5_0 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \c0.i15218_4_lut_LC_9_5_0  (
            .in0(N__28859),
            .in1(N__37843),
            .in2(N__28803),
            .in3(N__28824),
            .lcout(),
            .ltout(\c0.n18079_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i8_LC_9_5_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i8_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i8_LC_9_5_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.data_out_frame2_0___i8_LC_9_5_1  (
            .in0(N__28934),
            .in1(N__28793),
            .in2(N__28641),
            .in3(N__28986),
            .lcout(\c0.data_out_frame2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49835),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_661_LC_9_5_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_661_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_661_LC_9_5_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i12_4_lut_adj_661_LC_9_5_2  (
            .in0(N__28638),
            .in1(N__28629),
            .in2(N__28617),
            .in3(N__28605),
            .lcout(\c0.n28_adj_2403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15224_4_lut_LC_9_5_3 .C_ON=1'b0;
    defparam \c0.i15224_4_lut_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15224_4_lut_LC_9_5_3 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i15224_4_lut_LC_9_5_3  (
            .in0(N__28883),
            .in1(N__28791),
            .in2(N__44367),
            .in3(N__28860),
            .lcout(),
            .ltout(\c0.n18085_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i6_LC_9_5_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i6_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i6_LC_9_5_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i6_LC_9_5_4  (
            .in0(N__28792),
            .in1(N__28985),
            .in2(N__28938),
            .in3(N__28933),
            .lcout(\c0.data_out_frame2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49835),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15221_4_lut_LC_9_5_5 .C_ON=1'b0;
    defparam \c0.i15221_4_lut_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15221_4_lut_LC_9_5_5 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i15221_4_lut_LC_9_5_5  (
            .in0(N__28882),
            .in1(N__28787),
            .in2(N__41811),
            .in3(N__28858),
            .lcout(\c0.n18082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15527_3_lut_4_lut_LC_9_5_6 .C_ON=1'b0;
    defparam \c0.i15527_3_lut_4_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15527_3_lut_4_lut_LC_9_5_6 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \c0.i15527_3_lut_4_lut_LC_9_5_6  (
            .in0(N__30161),
            .in1(N__37842),
            .in2(N__30599),
            .in3(N__30049),
            .lcout(\c0.n18270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_707_LC_9_5_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_707_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_707_LC_9_5_7 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \c0.i1_4_lut_adj_707_LC_9_5_7  (
            .in0(N__33176),
            .in1(N__33283),
            .in2(N__30066),
            .in3(N__30124),
            .lcout(\c0.n6035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_9_6_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i0_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_9_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__30213),
            .in2(_gnd_net_),
            .in3(N__28758),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\c0.tx2.n16539 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i1_LC_9_6_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i1_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_9_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__30227),
            .in2(_gnd_net_),
            .in3(N__28755),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx2.n16539 ),
            .carryout(\c0.tx2.n16540 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i2_LC_9_6_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i2_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_9_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__30240),
            .in2(_gnd_net_),
            .in3(N__28752),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx2.n16540 ),
            .carryout(\c0.tx2.n16541 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i3_LC_9_6_3 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i3_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_9_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__30830),
            .in2(_gnd_net_),
            .in3(N__28749),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx2.n16541 ),
            .carryout(\c0.tx2.n16542 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i4_LC_9_6_4 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i4_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_9_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__30252),
            .in2(_gnd_net_),
            .in3(N__29100),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx2.n16542 ),
            .carryout(\c0.tx2.n16543 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i5_LC_9_6_5 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i5_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_9_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__30854),
            .in2(_gnd_net_),
            .in3(N__29097),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx2.n16543 ),
            .carryout(\c0.tx2.n16544 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i6_LC_9_6_6 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i6_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_9_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__29087),
            .in2(_gnd_net_),
            .in3(N__29073),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx2.n16544 ),
            .carryout(\c0.tx2.n16545 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i7_LC_9_6_7 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i7_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_9_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__29063),
            .in2(_gnd_net_),
            .in3(N__29049),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx2.n16545 ),
            .carryout(\c0.tx2.n16546 ),
            .clk(N__49827),
            .ce(N__30726),
            .sr(N__29021));
    defparam \c0.tx2.r_Clock_Count__i8_LC_9_7_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_9_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__29036),
            .in2(_gnd_net_),
            .in3(N__29046),
            .lcout(\c0.tx2.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49815),
            .ce(N__30725),
            .sr(N__29022));
    defparam \c0.add_2506_2_lut_LC_9_8_0 .C_ON=1'b1;
    defparam \c0.add_2506_2_lut_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_2_lut_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_2_lut_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__29127),
            .in2(N__42799),
            .in3(_gnd_net_),
            .lcout(\c0.tx_transmit_N_1947_0 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\c0.n16517 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_3_lut_LC_9_8_1 .C_ON=1'b1;
    defparam \c0.add_2506_3_lut_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_3_lut_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_3_lut_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__34774),
            .in2(_gnd_net_),
            .in3(N__28998),
            .lcout(\c0.tx_transmit_N_1947_1 ),
            .ltout(),
            .carryin(\c0.n16517 ),
            .carryout(\c0.n16518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_4_lut_LC_9_8_2 .C_ON=1'b1;
    defparam \c0.add_2506_4_lut_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_4_lut_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_4_lut_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__35144),
            .in2(_gnd_net_),
            .in3(N__28995),
            .lcout(\c0.tx_transmit_N_1947_2 ),
            .ltout(),
            .carryin(\c0.n16518 ),
            .carryout(\c0.n16519 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_5_lut_LC_9_8_3 .C_ON=1'b1;
    defparam \c0.add_2506_5_lut_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_5_lut_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_5_lut_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__35049),
            .in2(_gnd_net_),
            .in3(N__28992),
            .lcout(tx_transmit_N_1947_3),
            .ltout(),
            .carryin(\c0.n16519 ),
            .carryout(\c0.n16520 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_6_lut_LC_9_8_4 .C_ON=1'b1;
    defparam \c0.add_2506_6_lut_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_6_lut_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_6_lut_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__32484),
            .in2(_gnd_net_),
            .in3(N__29250),
            .lcout(tx_transmit_N_1947_4),
            .ltout(),
            .carryin(\c0.n16520 ),
            .carryout(\c0.n16521 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_7_lut_LC_9_8_5 .C_ON=1'b1;
    defparam \c0.add_2506_7_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_7_lut_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_7_lut_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__30927),
            .in2(_gnd_net_),
            .in3(N__29247),
            .lcout(\c0.tx_transmit_N_1947_5 ),
            .ltout(),
            .carryin(\c0.n16521 ),
            .carryout(\c0.n16522 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_8_lut_LC_9_8_6 .C_ON=1'b1;
    defparam \c0.add_2506_8_lut_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_8_lut_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_8_lut_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__30887),
            .in2(_gnd_net_),
            .in3(N__29244),
            .lcout(tx_transmit_N_1947_6),
            .ltout(),
            .carryin(\c0.n16522 ),
            .carryout(\c0.n16523 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_9_lut_LC_9_8_7 .C_ON=1'b0;
    defparam \c0.add_2506_9_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_9_lut_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_9_lut_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__31035),
            .in2(_gnd_net_),
            .in3(N__29241),
            .lcout(tx_transmit_N_1947_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i0_LC_9_9_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i0_LC_9_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i0_LC_9_9_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.byte_transmit_counter2_i0_LC_9_9_0  (
            .in0(N__30554),
            .in1(N__29238),
            .in2(N__30642),
            .in3(N__45952),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49791),
            .ce(),
            .sr(N__29223));
    defparam \c0.i1_2_lut_adj_759_LC_9_9_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_759_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_759_LC_9_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_759_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__36051),
            .in2(_gnd_net_),
            .in3(N__31911),
            .lcout(\c0.n10782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_9_9_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_9_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__29208),
            .in2(_gnd_net_),
            .in3(N__29181),
            .lcout(\c0.rx.n73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_9_9_5 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_9_9_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__29289),
            .in2(_gnd_net_),
            .in3(N__32120),
            .lcout(\c0.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_9_9_7 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_9_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29354),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_9_10_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_9_10_0  (
            .in0(N__32180),
            .in1(N__31347),
            .in2(N__31294),
            .in3(N__31398),
            .lcout(n9667),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__3__2253_LC_9_10_1 .C_ON=1'b0;
    defparam \c0.data_out_0__3__2253_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__3__2253_LC_9_10_1 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.data_out_0__3__2253_LC_9_10_1  (
            .in0(N__43411),
            .in1(N__36584),
            .in2(_gnd_net_),
            .in3(N__46960),
            .lcout(data_out_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_2167_LC_9_10_2 .C_ON=1'b0;
    defparam \c0.tx_active_prev_2167_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_2167_LC_9_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx_active_prev_2167_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32130),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1__2284_LC_9_10_3 .C_ON=1'b0;
    defparam \c0.data_in_1__1__2284_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1__2284_LC_9_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__1__2284_LC_9_10_3  (
            .in0(N__34227),
            .in1(N__29274),
            .in2(_gnd_net_),
            .in3(N__34281),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__7__2241_LC_9_10_4 .C_ON=1'b0;
    defparam \c0.data_out_1__7__2241_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__7__2241_LC_9_10_4 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \c0.data_out_1__7__2241_LC_9_10_4  (
            .in0(N__46959),
            .in1(N__43412),
            .in2(_gnd_net_),
            .in3(N__29322),
            .lcout(data_out_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_585_LC_9_10_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_585_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_585_LC_9_10_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_585_LC_9_10_5  (
            .in0(N__47228),
            .in1(N__47685),
            .in2(_gnd_net_),
            .in3(N__46958),
            .lcout(n10973),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_9_10_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_9_10_6 .LUT_INIT=16'b0101111100001100;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_9_10_6  (
            .in0(N__29328),
            .in1(N__30906),
            .in2(N__31295),
            .in3(N__32129),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_10_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_9_10_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_9_10_7  (
            .in0(N__33706),
            .in1(N__33748),
            .in2(_gnd_net_),
            .in3(N__33914),
            .lcout(r_Bit_Index_0_adj_2519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15180_3_lut_LC_9_11_0 .C_ON=1'b0;
    defparam \c0.tx.i15180_3_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15180_3_lut_LC_9_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx.i15180_3_lut_LC_9_11_0  (
            .in0(N__32322),
            .in1(N__31632),
            .in2(_gnd_net_),
            .in3(N__31149),
            .lcout(\c0.tx.n18041 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18747_bdd_4_lut_LC_9_11_1 .C_ON=1'b0;
    defparam \c0.n18747_bdd_4_lut_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18747_bdd_4_lut_LC_9_11_1 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18747_bdd_4_lut_LC_9_11_1  (
            .in0(N__35220),
            .in1(N__29493),
            .in2(N__31578),
            .in3(N__34359),
            .lcout(n18750),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_11_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_11_2 .LUT_INIT=16'b1101110110011001;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_11_2  (
            .in0(N__31348),
            .in1(N__31285),
            .in2(_gnd_net_),
            .in3(N__29301),
            .lcout(),
            .ltout(n3_adj_2525_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_9_11_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_9_11_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__29353),
            .in2(N__29370),
            .in3(N__29479),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_3_lut_LC_9_11_4 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_3_lut_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_3_lut_LC_9_11_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.tx.i2_3_lut_3_lut_LC_9_11_4  (
            .in0(N__31349),
            .in1(N__31399),
            .in2(_gnd_net_),
            .in3(N__31215),
            .lcout(\c0.tx.n17697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15687_2_lut_LC_9_11_5 .C_ON=1'b0;
    defparam \c0.i15687_2_lut_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15687_2_lut_LC_9_11_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i15687_2_lut_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__42707),
            .in2(_gnd_net_),
            .in3(N__29321),
            .lcout(\c0.n18354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_4_lut_LC_9_11_6 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_4_lut_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_4_lut_LC_9_11_6 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx.i1_3_lut_4_lut_LC_9_11_6  (
            .in0(N__31350),
            .in1(N__31400),
            .in2(N__31296),
            .in3(N__31216),
            .lcout(),
            .ltout(\c0.tx.n11030_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_9_11_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_9_11_7 .LUT_INIT=16'b0000101001001010;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_9_11_7  (
            .in0(N__31150),
            .in1(N__31289),
            .in2(N__29310),
            .in3(N__31074),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n18711_bdd_4_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \c0.tx.n18711_bdd_4_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n18711_bdd_4_lut_LC_9_12_3 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \c0.tx.n18711_bdd_4_lut_LC_9_12_3  (
            .in0(N__31413),
            .in1(N__29307),
            .in2(N__31461),
            .in3(N__31434),
            .lcout(\c0.tx.o_Tx_Serial_N_2062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15306_3_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \c0.tx.i15306_3_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15306_3_lut_LC_9_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i15306_3_lut_LC_9_12_4  (
            .in0(N__31154),
            .in1(N__29381),
            .in2(_gnd_net_),
            .in3(N__29408),
            .lcout(\c0.tx.n18167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_817_LC_9_12_5.C_ON=1'b0;
    defparam i24_4_lut_adj_817_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_817_LC_9_12_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 i24_4_lut_adj_817_LC_9_12_5 (
            .in0(N__35230),
            .in1(N__29295),
            .in2(N__30897),
            .in3(N__35081),
            .lcout(),
            .ltout(n10_adj_2532_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_9_12_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_12_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_9_12_6  (
            .in0(N__32523),
            .in1(N__32570),
            .in2(N__29412),
            .in3(N__29409),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49750),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_528_LC_9_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_528_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_528_LC_9_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_528_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__32352),
            .in2(_gnd_net_),
            .in3(N__37335),
            .lcout(\c0.n10749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_9_13_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_9_13_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_9_13_1  (
            .in0(N__31214),
            .in1(N__31327),
            .in2(N__31293),
            .in3(N__31395),
            .lcout(\c0.tx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_9_13_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_9_13_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_9_13_2  (
            .in0(N__31396),
            .in1(N__31275),
            .in2(N__31345),
            .in3(N__31213),
            .lcout(\c0.tx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15125_2_lut_LC_9_13_3 .C_ON=1'b0;
    defparam \c0.tx.i15125_2_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15125_2_lut_LC_9_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i15125_2_lut_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__31252),
            .in2(_gnd_net_),
            .in3(N__31326),
            .lcout(\c0.tx.n17984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__4__2188_LC_9_13_4 .C_ON=1'b0;
    defparam \c0.data_out_8__4__2188_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__4__2188_LC_9_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__4__2188_LC_9_13_4  (
            .in0(N__46847),
            .in1(N__38058),
            .in2(_gnd_net_),
            .in3(N__36708),
            .lcout(data_out_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_9_13_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_9_13_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_9_13_5  (
            .in0(N__42812),
            .in1(N__31407),
            .in2(N__36663),
            .in3(N__34870),
            .lcout(),
            .ltout(n10_adj_2537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_815_LC_9_13_6.C_ON=1'b0;
    defparam i24_4_lut_adj_815_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_815_LC_9_13_6.LUT_INIT=16'b0100010011100100;
    LogicCell40 i24_4_lut_adj_815_LC_9_13_6 (
            .in0(N__35092),
            .in1(N__29433),
            .in2(N__29388),
            .in3(N__35246),
            .lcout(),
            .ltout(n10_adj_2535_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_9_13_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_9_13_7  (
            .in0(N__32585),
            .in1(N__29382),
            .in2(N__29385),
            .in3(N__32529),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15574_2_lut_LC_9_14_0 .C_ON=1'b0;
    defparam \c0.i15574_2_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15574_2_lut_LC_9_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15574_2_lut_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__29427),
            .in2(_gnd_net_),
            .in3(N__42808),
            .lcout(\c0.n18188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__7__2185_LC_9_14_1 .C_ON=1'b0;
    defparam \c0.data_out_8__7__2185_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__7__2185_LC_9_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__7__2185_LC_9_14_1  (
            .in0(N__46855),
            .in1(N__38748),
            .in2(_gnd_net_),
            .in3(N__32357),
            .lcout(data_out_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_603_LC_9_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_603_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_603_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_603_LC_9_14_2  (
            .in0(N__32681),
            .in1(N__42606),
            .in2(_gnd_net_),
            .in3(N__34565),
            .lcout(\c0.n17883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_1_lut_LC_9_14_5 .C_ON=1'b0;
    defparam \c0.tx.i2_1_lut_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_1_lut_LC_9_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.i2_1_lut_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31380),
            .lcout(n5155),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18753_bdd_4_lut_LC_9_14_7 .C_ON=1'b0;
    defparam \c0.n18753_bdd_4_lut_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18753_bdd_4_lut_LC_9_14_7 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18753_bdd_4_lut_LC_9_14_7  (
            .in0(N__29538),
            .in1(N__31554),
            .in2(N__29445),
            .in3(N__35245),
            .lcout(n18756),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__6__2226_LC_9_15_0 .C_ON=1'b0;
    defparam \c0.data_out_3__6__2226_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6__2226_LC_9_15_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.data_out_3__6__2226_LC_9_15_0  (
            .in0(N__47668),
            .in1(N__29426),
            .in2(N__43409),
            .in3(N__47121),
            .lcout(\c0.data_out_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_9_15_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_9_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_9_15_1  (
            .in0(N__42800),
            .in1(N__39908),
            .in2(_gnd_net_),
            .in3(N__36776),
            .lcout(\c0.n5_adj_2241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_9_15_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_9_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_9_15_3  (
            .in0(N__42801),
            .in1(N__31610),
            .in2(_gnd_net_),
            .in3(N__31698),
            .lcout(\c0.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__7__2233_LC_9_16_2 .C_ON=1'b0;
    defparam \c0.data_out_2__7__2233_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__7__2233_LC_9_16_2 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \c0.data_out_2__7__2233_LC_9_16_2  (
            .in0(N__47115),
            .in1(_gnd_net_),
            .in2(N__29550),
            .in3(N__43372),
            .lcout(data_out_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49704),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__6__2242_LC_9_16_5 .C_ON=1'b0;
    defparam \c0.data_out_1__6__2242_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6__2242_LC_9_16_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.data_out_1__6__2242_LC_9_16_5  (
            .in0(N__31599),
            .in1(N__47400),
            .in2(N__43410),
            .in3(N__47117),
            .lcout(data_out_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49704),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__7__2225_LC_9_16_6 .C_ON=1'b0;
    defparam \c0.data_out_3__7__2225_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7__2225_LC_9_16_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_3__7__2225_LC_9_16_6  (
            .in0(N__47116),
            .in1(N__43376),
            .in2(N__29562),
            .in3(N__47401),
            .lcout(data_out_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49704),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_9_16_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_9_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_9_16_7  (
            .in0(N__42811),
            .in1(N__29558),
            .in2(_gnd_net_),
            .in3(N__29546),
            .lcout(\c0.n2_adj_2229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_1266_i1_3_lut_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.mux_1266_i1_3_lut_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_1266_i1_3_lut_LC_9_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_1266_i1_3_lut_LC_9_17_0  (
            .in0(N__47677),
            .in1(N__47394),
            .in2(_gnd_net_),
            .in3(N__47111),
            .lcout(n2837),
            .ltout(n2837_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__5__2251_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.data_out_0__5__2251_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5__2251_LC_9_17_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_out_0__5__2251_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__43319),
            .in2(N__29529),
            .in3(N__29526),
            .lcout(data_out_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15651_2_lut_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.i15651_2_lut_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15651_2_lut_LC_9_18_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15651_2_lut_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__29525),
            .in2(_gnd_net_),
            .in3(N__42860),
            .lcout(\c0.n18189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i2658_4_lut_LC_9_22_5 .C_ON=1'b0;
    defparam \control.i2658_4_lut_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \control.i2658_4_lut_LC_9_22_5 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \control.i2658_4_lut_LC_9_22_5  (
            .in0(N__29642),
            .in1(N__29627),
            .in2(N__29661),
            .in3(N__29675),
            .lcout(),
            .ltout(\control.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i2661_4_lut_LC_9_22_6 .C_ON=1'b0;
    defparam \control.i2661_4_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \control.i2661_4_lut_LC_9_22_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \control.i2661_4_lut_LC_9_22_6  (
            .in0(N__29597),
            .in1(N__29583),
            .in2(N__29514),
            .in3(N__29612),
            .lcout(\control.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i0_LC_9_23_0 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i0_LC_9_23_0 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i0_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i0_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__29511),
            .in2(_gnd_net_),
            .in3(N__29505),
            .lcout(\control.n10 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\control.n16647 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i1_LC_9_23_1 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i1_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i1_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i1_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__29502),
            .in2(_gnd_net_),
            .in3(N__29496),
            .lcout(\control.n9_adj_2459 ),
            .ltout(),
            .carryin(\control.n16647 ),
            .carryout(\control.n16648 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i2_LC_9_23_2 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i2_LC_9_23_2 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i2_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i2_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__29676),
            .in2(_gnd_net_),
            .in3(N__29664),
            .lcout(\control.pwm_delay_2 ),
            .ltout(),
            .carryin(\control.n16648 ),
            .carryout(\control.n16649 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i3_LC_9_23_3 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i3_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i3_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i3_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__29660),
            .in2(_gnd_net_),
            .in3(N__29646),
            .lcout(\control.pwm_delay_3 ),
            .ltout(),
            .carryin(\control.n16649 ),
            .carryout(\control.n16650 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i4_LC_9_23_4 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i4_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i4_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i4_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__29643),
            .in2(_gnd_net_),
            .in3(N__29631),
            .lcout(\control.pwm_delay_4 ),
            .ltout(),
            .carryin(\control.n16650 ),
            .carryout(\control.n16651 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i5_LC_9_23_5 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i5_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i5_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i5_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__29628),
            .in2(_gnd_net_),
            .in3(N__29616),
            .lcout(\control.pwm_delay_5 ),
            .ltout(),
            .carryin(\control.n16651 ),
            .carryout(\control.n16652 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i6_LC_9_23_6 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i6_LC_9_23_6 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i6_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i6_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__29613),
            .in2(_gnd_net_),
            .in3(N__29601),
            .lcout(\control.pwm_delay_6 ),
            .ltout(),
            .carryin(\control.n16652 ),
            .carryout(\control.n16653 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i7_LC_9_23_7 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i7_LC_9_23_7 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i7_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i7_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__29598),
            .in2(_gnd_net_),
            .in3(N__29586),
            .lcout(\control.pwm_delay_7 ),
            .ltout(),
            .carryin(\control.n16653 ),
            .carryout(\control.n16654 ),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i8_LC_9_24_0 .C_ON=1'b1;
    defparam \control.pwm_delay_2485__i8_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i8_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i8_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__29582),
            .in2(_gnd_net_),
            .in3(N__29568),
            .lcout(\control.pwm_delay_8 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\control.n16655 ),
            .clk(N__49778),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.pwm_delay_2485__i9_LC_9_24_1 .C_ON=1'b0;
    defparam \control.pwm_delay_2485__i9_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \control.pwm_delay_2485__i9_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \control.pwm_delay_2485__i9_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__32900),
            .in2(_gnd_net_),
            .in3(N__29565),
            .lcout(\control.pwm_delay_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18885_bdd_4_lut_LC_10_1_0 .C_ON=1'b0;
    defparam \c0.n18885_bdd_4_lut_LC_10_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18885_bdd_4_lut_LC_10_1_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18885_bdd_4_lut_LC_10_1_0  (
            .in0(N__49075),
            .in1(N__29754),
            .in2(N__31731),
            .in3(N__29694),
            .lcout(),
            .ltout(\c0.n18888_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_10_1_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_10_1_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_10_1_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_10_1_1  (
            .in0(N__29700),
            .in1(N__49076),
            .in2(N__29709),
            .in3(N__48927),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49867),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15904_LC_10_1_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15904_LC_10_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15904_LC_10_1_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15904_LC_10_1_2  (
            .in0(N__31827),
            .in1(N__48602),
            .in2(N__31659),
            .in3(N__46162),
            .lcout(),
            .ltout(\c0.n18789_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18789_bdd_4_lut_LC_10_1_3 .C_ON=1'b0;
    defparam \c0.n18789_bdd_4_lut_LC_10_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18789_bdd_4_lut_LC_10_1_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18789_bdd_4_lut_LC_10_1_3  (
            .in0(N__48603),
            .in1(N__29724),
            .in2(N__29706),
            .in3(N__35904),
            .lcout(),
            .ltout(\c0.n18792_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_10_1_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_10_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_10_1_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_10_1_4  (
            .in0(N__48035),
            .in1(N__37899),
            .in2(N__29703),
            .in3(N__48170),
            .lcout(\c0.n22_adj_2270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_10_1_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_10_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_10_1_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_10_1_5  (
            .in0(N__33531),
            .in1(N__49074),
            .in2(N__29685),
            .in3(N__48034),
            .lcout(\c0.n18885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_494_LC_10_2_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_494_LC_10_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_494_LC_10_2_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_494_LC_10_2_0  (
            .in0(N__43661),
            .in1(N__40751),
            .in2(N__45801),
            .in3(N__40976),
            .lcout(\c0.n10816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_758_LC_10_2_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_758_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_758_LC_10_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_758_LC_10_2_1  (
            .in0(_gnd_net_),
            .in1(N__41082),
            .in2(_gnd_net_),
            .in3(N__46415),
            .lcout(),
            .ltout(\c0.n10861_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_775_LC_10_2_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_775_LC_10_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_775_LC_10_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_775_LC_10_2_2  (
            .in0(N__45357),
            .in1(N__40437),
            .in2(N__29688),
            .in3(N__40803),
            .lcout(\c0.n20_adj_2442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18795_bdd_4_lut_LC_10_2_3 .C_ON=1'b0;
    defparam \c0.n18795_bdd_4_lut_LC_10_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18795_bdd_4_lut_LC_10_2_3 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18795_bdd_4_lut_LC_10_2_3  (
            .in0(N__48623),
            .in1(N__31767),
            .in2(N__41722),
            .in3(N__33333),
            .lcout(\c0.n18798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_780_LC_10_2_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_780_LC_10_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_780_LC_10_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_780_LC_10_2_4  (
            .in0(_gnd_net_),
            .in1(N__31857),
            .in2(_gnd_net_),
            .in3(N__45202),
            .lcout(\c0.n10893 ),
            .ltout(\c0.n10893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_781_LC_10_2_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_781_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_781_LC_10_2_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_781_LC_10_2_5  (
            .in0(N__41674),
            .in1(N__36335),
            .in2(N__29727),
            .in3(N__44167),
            .lcout(\c0.n17886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_705_LC_10_2_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_705_LC_10_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_705_LC_10_2_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_705_LC_10_2_6  (
            .in0(_gnd_net_),
            .in1(N__33383),
            .in2(_gnd_net_),
            .in3(N__31856),
            .lcout(\c0.n18_adj_2423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_483_LC_10_2_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_483_LC_10_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_483_LC_10_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_483_LC_10_2_7  (
            .in0(N__45815),
            .in1(N__41036),
            .in2(_gnd_net_),
            .in3(N__43662),
            .lcout(\c0.n17911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_10_3_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_10_3_0 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_10_3_0  (
            .in0(N__46090),
            .in1(N__40844),
            .in2(N__50743),
            .in3(_gnd_net_),
            .lcout(\c0.n5_adj_2433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_3_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_3_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_3_1  (
            .in0(N__48161),
            .in1(N__31773),
            .in2(N__48033),
            .in3(N__31716),
            .lcout(\c0.n22_adj_2373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_788_LC_10_3_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_788_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_788_LC_10_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_788_LC_10_3_2  (
            .in0(N__41078),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37139),
            .lcout(\c0.n17748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_508_LC_10_3_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_508_LC_10_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_508_LC_10_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_508_LC_10_3_3  (
            .in0(N__37138),
            .in1(N__41077),
            .in2(_gnd_net_),
            .in3(N__45206),
            .lcout(\c0.n10688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_10_3_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_10_3_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_10_3_4 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_10_3_4  (
            .in0(N__30773),
            .in1(N__29889),
            .in2(N__30366),
            .in3(N__29842),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i138_LC_10_3_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i138_LC_10_3_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i138_LC_10_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i138_LC_10_3_5  (
            .in0(N__38660),
            .in1(N__29723),
            .in2(_gnd_net_),
            .in3(N__50451),
            .lcout(data_out_frame2_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_10_3_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_10_3_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_10_3_6  (
            .in0(N__46091),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__41190),
            .lcout(),
            .ltout(\c0.n5_adj_2435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_3_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_3_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_3_7  (
            .in0(N__48624),
            .in1(N__44660),
            .in2(N__29802),
            .in3(N__46092),
            .lcout(\c0.n6_adj_2223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_10_4_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_10_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_10_4_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_10_4_0  (
            .in0(N__30439),
            .in1(N__30774),
            .in2(N__29849),
            .in3(N__30368),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15828_LC_10_4_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15828_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15828_LC_10_4_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15828_LC_10_4_1  (
            .in0(N__46187),
            .in1(N__36049),
            .in2(N__48649),
            .in3(N__45248),
            .lcout(),
            .ltout(\c0.n18687_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18687_bdd_4_lut_LC_10_4_2 .C_ON=1'b0;
    defparam \c0.n18687_bdd_4_lut_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18687_bdd_4_lut_LC_10_4_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18687_bdd_4_lut_LC_10_4_2  (
            .in0(N__48556),
            .in1(N__44624),
            .in2(N__29787),
            .in3(N__36314),
            .lcout(\c0.n18690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_518_LC_10_4_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_518_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_518_LC_10_4_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_518_LC_10_4_3  (
            .in0(N__44742),
            .in1(N__44899),
            .in2(N__44805),
            .in3(N__41405),
            .lcout(\c0.n17795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_4_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_4_4 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_4_4  (
            .in0(N__48557),
            .in1(N__31854),
            .in2(N__29772),
            .in3(N__46188),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_10_4_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_10_4_5 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_10_4_5  (
            .in0(N__46189),
            .in1(N__44820),
            .in2(N__37792),
            .in3(N__48558),
            .lcout(\c0.n6_adj_2354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15973_LC_10_4_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15973_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15973_LC_10_4_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15973_LC_10_4_6  (
            .in0(N__43656),
            .in1(N__44741),
            .in2(N__48648),
            .in3(N__46186),
            .lcout(\c0.n18855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i46_LC_10_4_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i46_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i46_LC_10_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i46_LC_10_4_7  (
            .in0(N__37785),
            .in1(N__39354),
            .in2(_gnd_net_),
            .in3(N__50445),
            .lcout(data_out_frame2_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10936_2_lut_LC_10_5_0 .C_ON=1'b0;
    defparam \c0.i10936_2_lut_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10936_2_lut_LC_10_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i10936_2_lut_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__29918),
            .in2(_gnd_net_),
            .in3(N__30192),
            .lcout(\c0.n12359 ),
            .ltout(\c0.n12359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_782_LC_10_5_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_782_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_782_LC_10_5_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.i2_4_lut_adj_782_LC_10_5_1  (
            .in0(N__30162),
            .in1(N__33175),
            .in2(N__30138),
            .in3(N__33290),
            .lcout(),
            .ltout(\c0.n6_adj_2443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_2261_LC_10_5_2 .C_ON=1'b0;
    defparam \c0.tx2_transmit_2261_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_2261_LC_10_5_2 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \c0.tx2_transmit_2261_LC_10_5_2  (
            .in0(N__33291),
            .in1(N__33177),
            .in2(N__30135),
            .in3(N__30050),
            .lcout(\c0.r_SM_Main_2_N_2034_0_adj_2213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49836),
            .ce(),
            .sr(N__30131));
    defparam \c0.i1_2_lut_adj_448_LC_10_5_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_448_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_448_LC_10_5_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i1_2_lut_adj_448_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__30045),
            .in2(_gnd_net_),
            .in3(N__33174),
            .lcout(\c0.n10958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4167_4_lut_LC_10_5_4 .C_ON=1'b0;
    defparam \c0.tx2.i4167_4_lut_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4167_4_lut_LC_10_5_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.tx2.i4167_4_lut_LC_10_5_4  (
            .in0(N__30450),
            .in1(N__29828),
            .in2(N__29927),
            .in3(N__30438),
            .lcout(n6707),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11346_2_lut_4_lut_LC_10_5_5 .C_ON=1'b0;
    defparam \c0.tx2.i11346_2_lut_4_lut_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11346_2_lut_4_lut_LC_10_5_5 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \c0.tx2.i11346_2_lut_4_lut_LC_10_5_5  (
            .in0(N__29877),
            .in1(N__30855),
            .in2(N__30831),
            .in3(N__30201),
            .lcout(r_SM_Main_2_N_2031_1),
            .ltout(r_SM_Main_2_N_2031_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15154_3_lut_4_lut_LC_10_5_6 .C_ON=1'b0;
    defparam \c0.tx2.i15154_3_lut_4_lut_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15154_3_lut_4_lut_LC_10_5_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \c0.tx2.i15154_3_lut_4_lut_LC_10_5_6  (
            .in0(N__30356),
            .in1(N__30436),
            .in2(N__29808),
            .in3(N__30769),
            .lcout(n18014),
            .ltout(n18014_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15159_3_lut_LC_10_5_7 .C_ON=1'b0;
    defparam \c0.tx2.i15159_3_lut_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15159_3_lut_LC_10_5_7 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \c0.tx2.i15159_3_lut_LC_10_5_7  (
            .in0(N__30437),
            .in1(_gnd_net_),
            .in2(N__29805),
            .in3(N__30449),
            .lcout(n11545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i4_LC_10_6_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i4_LC_10_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i4_LC_10_6_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i4_LC_10_6_0  (
            .in0(N__30675),
            .in1(N__48891),
            .in2(N__30600),
            .in3(N__30553),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49828),
            .ce(),
            .sr(N__30459));
    defparam \c0.tx2.i1_2_lut_LC_10_6_5 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_LC_10_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i1_2_lut_LC_10_6_5  (
            .in0(N__33885),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33938),
            .lcout(n4_adj_2472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_LC_10_6_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_10_6_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_LC_10_6_6  (
            .in0(N__33937),
            .in1(N__33680),
            .in2(_gnd_net_),
            .in3(N__33884),
            .lcout(\c0.tx2.n13800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15201_3_lut_LC_10_6_7 .C_ON=1'b0;
    defparam \c0.tx2.i15201_3_lut_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15201_3_lut_LC_10_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx2.i15201_3_lut_LC_10_6_7  (
            .in0(N__42387),
            .in1(N__43074),
            .in2(_gnd_net_),
            .in3(N__33936),
            .lcout(\c0.tx2.n18062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_7_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_7_0 .LUT_INIT=16'b1011101110011001;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_7_0  (
            .in0(N__30440),
            .in1(N__30367),
            .in2(_gnd_net_),
            .in3(N__30258),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_1__bdd_4_lut_LC_10_7_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_1__bdd_4_lut_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_1__bdd_4_lut_LC_10_7_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.tx2.r_Bit_Index_1__bdd_4_lut_LC_10_7_1  (
            .in0(N__33883),
            .in1(N__30294),
            .in2(N__33681),
            .in3(N__30282),
            .lcout(),
            .ltout(\c0.tx2.n18717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18717_bdd_4_lut_LC_10_7_2 .C_ON=1'b0;
    defparam \c0.tx2.n18717_bdd_4_lut_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18717_bdd_4_lut_LC_10_7_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.tx2.n18717_bdd_4_lut_LC_10_7_2  (
            .in0(N__30267),
            .in1(N__30789),
            .in2(N__30261),
            .in3(N__33679),
            .lcout(\c0.tx2.o_Tx_Serial_N_2062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4_4_lut_LC_10_7_3 .C_ON=1'b0;
    defparam \c0.tx2.i4_4_lut_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4_4_lut_LC_10_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx2.i4_4_lut_LC_10_7_3  (
            .in0(N__30251),
            .in1(N__30239),
            .in2(N__30228),
            .in3(N__30212),
            .lcout(\c0.tx2.n10 ),
            .ltout(\c0.tx2.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5_3_lut_LC_10_7_4 .C_ON=1'b0;
    defparam \c0.tx2.i5_3_lut_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5_3_lut_LC_10_7_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.tx2.i5_3_lut_LC_10_7_4  (
            .in0(N__30853),
            .in1(_gnd_net_),
            .in2(N__30834),
            .in3(N__30829),
            .lcout(\c0.tx2.n12775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15200_3_lut_LC_10_7_5 .C_ON=1'b0;
    defparam \c0.tx2.i15200_3_lut_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15200_3_lut_LC_10_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx2.i15200_3_lut_LC_10_7_5  (
            .in0(N__30798),
            .in1(N__49179),
            .in2(_gnd_net_),
            .in3(N__33939),
            .lcout(\c0.tx2.n18061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i13_1_lut_LC_10_7_7 .C_ON=1'b0;
    defparam \c0.tx2.i13_1_lut_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i13_1_lut_LC_10_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.i13_1_lut_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30782),
            .lcout(n11096),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15706_3_lut_4_lut_LC_10_8_0 .C_ON=1'b0;
    defparam \c0.i15706_3_lut_4_lut_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15706_3_lut_4_lut_LC_10_8_0 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \c0.i15706_3_lut_4_lut_LC_10_8_0  (
            .in0(N__33834),
            .in1(N__33450),
            .in2(N__47672),
            .in3(N__33794),
            .lcout(),
            .ltout(\c0.n18260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_2168_LC_10_8_1 .C_ON=1'b0;
    defparam \c0.tx_transmit_2168_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_2168_LC_10_8_1 .LUT_INIT=16'b0000001000010011;
    LogicCell40 \c0.tx_transmit_2168_LC_10_8_1  (
            .in0(N__30690),
            .in1(N__30696),
            .in2(N__30699),
            .in3(N__33765),
            .lcout(\c0.r_SM_Main_2_N_2034_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49805),
            .ce(),
            .sr(N__30684));
    defparam \c0.i1_2_lut_3_lut_adj_637_LC_10_8_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_637_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_637_LC_10_8_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_637_LC_10_8_2  (
            .in0(N__32132),
            .in1(_gnd_net_),
            .in2(N__32178),
            .in3(N__47291),
            .lcout(\c0.n130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10860_2_lut_LC_10_8_3 .C_ON=1'b0;
    defparam \c0.i10860_2_lut_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10860_2_lut_LC_10_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i10860_2_lut_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__32164),
            .in2(_gnd_net_),
            .in3(N__32131),
            .lcout(n12227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_LC_10_8_5 .C_ON=1'b0;
    defparam \c0.i6_3_lut_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_LC_10_8_5 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \c0.i6_3_lut_LC_10_8_5  (
            .in0(N__47292),
            .in1(_gnd_net_),
            .in2(N__47691),
            .in3(N__47059),
            .lcout(\c0.n3465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_10_8_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_10_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_10_8_6  (
            .in0(N__47058),
            .in1(N__47681),
            .in2(_gnd_net_),
            .in3(N__47293),
            .lcout(\c0.n4806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_10_8_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_10_8_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_10_8_7  (
            .in0(N__33515),
            .in1(N__33490),
            .in2(_gnd_net_),
            .in3(N__33469),
            .lcout(\c0.n85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_10_9_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_10_9_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_10_9_1  (
            .in0(N__30876),
            .in1(N__30888),
            .in2(N__31005),
            .in3(N__30950),
            .lcout(byte_transmit_counter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_533_LC_10_9_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_533_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_533_LC_10_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_533_LC_10_9_2  (
            .in0(N__31016),
            .in1(N__30875),
            .in2(N__30867),
            .in3(N__31046),
            .lcout(\c0.n14068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_10_9_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_10_9_3 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_10_9_3  (
            .in0(N__32506),
            .in1(N__30866),
            .in2(N__31004),
            .in3(N__30949),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_10_9_4.C_ON=1'b0;
    defparam i2_4_lut_LC_10_9_4.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_10_9_4.LUT_INIT=16'b0000000100000000;
    LogicCell40 i2_4_lut_LC_10_9_4 (
            .in0(N__32019),
            .in1(N__33402),
            .in2(N__31920),
            .in3(N__32187),
            .lcout(UART_TRANSMITTER_state_7_N_1223_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_10_9_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_10_9_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_10_9_5  (
            .in0(N__30993),
            .in1(N__35071),
            .in2(N__33858),
            .in3(N__30948),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_10_9_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i1_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_10_9_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_10_9_6  (
            .in0(N__30951),
            .in1(N__30989),
            .in2(N__34856),
            .in3(N__33491),
            .lcout(byte_transmit_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_10_9_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_10_9_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_10_9_7  (
            .in0(N__35190),
            .in1(N__33470),
            .in2(N__31003),
            .in3(N__30952),
            .lcout(byte_transmit_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_10_10_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i0_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_10_10_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_10_10_0  (
            .in0(N__33516),
            .in1(N__42798),
            .in2(N__31001),
            .in3(N__30953),
            .lcout(byte_transmit_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_437_LC_10_10_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_437_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_437_LC_10_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_437_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__47260),
            .in2(_gnd_net_),
            .in3(N__32293),
            .lcout(),
            .ltout(\c0.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_10_10_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_10_10_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \c0.i2_4_lut_LC_10_10_2  (
            .in0(N__30982),
            .in1(N__34376),
            .in2(N__31056),
            .in3(N__30912),
            .lcout(n5341),
            .ltout(n5341_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_10_10_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_10_10_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_10_10_3  (
            .in0(N__31000),
            .in1(N__31034),
            .in2(N__31053),
            .in3(N__31050),
            .lcout(byte_transmit_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_10_10_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_10_10_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_10_10_4  (
            .in0(N__30926),
            .in1(N__31020),
            .in2(N__31002),
            .in3(N__30954),
            .lcout(\c0.byte_transmit_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15139_4_lut_LC_10_10_5 .C_ON=1'b0;
    defparam \c0.i15139_4_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15139_4_lut_LC_10_10_5 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \c0.i15139_4_lut_LC_10_10_5  (
            .in0(N__32024),
            .in1(N__47259),
            .in2(N__47615),
            .in3(N__32193),
            .lcout(\c0.n17998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15079_2_lut_3_lut_3_lut_LC_10_10_7 .C_ON=1'b0;
    defparam \c0.tx.i15079_2_lut_3_lut_3_lut_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15079_2_lut_3_lut_3_lut_LC_10_10_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.tx.i15079_2_lut_3_lut_3_lut_LC_10_10_7  (
            .in0(N__32179),
            .in1(N__31346),
            .in2(_gnd_net_),
            .in3(N__31397),
            .lcout(\c0.tx.n17938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i2_LC_10_11_0 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i2_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i2_LC_10_11_0 .LUT_INIT=16'b1010011011000110;
    LogicCell40 \c0.UART_TRANSMITTER_state__i2_LC_10_11_0  (
            .in0(N__46962),
            .in1(N__47257),
            .in2(N__47614),
            .in3(N__32262),
            .lcout(UART_TRANSMITTER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i1_LC_10_11_1 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_10_11_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.UART_TRANSMITTER_state__i1_LC_10_11_1  (
            .in0(N__47256),
            .in1(N__32241),
            .in2(N__47669),
            .in3(N__32280),
            .lcout(UART_TRANSMITTER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_10_11_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_10_11_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_10_11_2  (
            .in0(N__37101),
            .in1(N__34844),
            .in2(N__31083),
            .in3(N__42708),
            .lcout(n10_adj_2536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2723_2_lut_LC_10_11_3 .C_ON=1'b0;
    defparam \c0.tx.i2723_2_lut_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2723_2_lut_LC_10_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx.i2723_2_lut_LC_10_11_3  (
            .in0(N__31152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31487),
            .lcout(),
            .ltout(n5440_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_10_11_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_11_4 .LUT_INIT=16'b1001110000000000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_10_11_4  (
            .in0(N__31170),
            .in1(N__31459),
            .in2(N__31095),
            .in3(N__31092),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15156_2_lut_3_lut_LC_10_11_5 .C_ON=1'b0;
    defparam \c0.tx.i15156_2_lut_3_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15156_2_lut_3_lut_LC_10_11_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.tx.i15156_2_lut_3_lut_LC_10_11_5  (
            .in0(N__31291),
            .in1(N__31073),
            .in2(_gnd_net_),
            .in3(N__31168),
            .lcout(n18016),
            .ltout(n18016_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_10_11_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_10_11_6 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_10_11_6  (
            .in0(N__31169),
            .in1(N__31488),
            .in2(N__31086),
            .in3(N__31153),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_636_LC_10_11_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_636_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_636_LC_10_11_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_636_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__47536),
            .in2(_gnd_net_),
            .in3(N__46961),
            .lcout(n9_adj_2477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_10_12_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_10_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_10_12_1  (
            .in0(N__42781),
            .in1(N__34492),
            .in2(_gnd_net_),
            .in3(N__37443),
            .lcout(\c0.n8_adj_2207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_10_12_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_10_12_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_10_12_2  (
            .in0(N__31427),
            .in1(N__32226),
            .in2(N__32600),
            .in3(N__32524),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_LC_10_12_3 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_LC_10_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_LC_10_12_3  (
            .in0(N__31151),
            .in1(N__31486),
            .in2(_gnd_net_),
            .in3(N__31455),
            .lcout(\c0.tx.n13802 ),
            .ltout(\c0.tx.n13802_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4255_4_lut_LC_10_12_4 .C_ON=1'b0;
    defparam \c0.tx.i4255_4_lut_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4255_4_lut_LC_10_12_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.tx.i4255_4_lut_LC_10_12_4  (
            .in0(N__31292),
            .in1(N__31217),
            .in2(N__31062),
            .in3(N__32181),
            .lcout(),
            .ltout(\c0.tx.n6796_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_10_12_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_10_12_5 .LUT_INIT=16'b0001000100110000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_10_12_5  (
            .in0(N__31218),
            .in1(N__31401),
            .in2(N__31059),
            .in3(N__31344),
            .lcout(\c0.tx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49751),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_6  (
            .in0(N__31485),
            .in1(N__31467),
            .in2(N__31460),
            .in3(N__31101),
            .lcout(\c0.tx.n18711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15179_3_lut_LC_10_12_7 .C_ON=1'b0;
    defparam \c0.tx.i15179_3_lut_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15179_3_lut_LC_10_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx.i15179_3_lut_LC_10_12_7  (
            .in0(N__31428),
            .in1(N__32457),
            .in2(_gnd_net_),
            .in3(N__31148),
            .lcout(\c0.tx.n18040 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_10_13_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_10_13_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_10_13_0  (
            .in0(N__31110),
            .in1(N__31521),
            .in2(N__32613),
            .in3(N__32530),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_10_13_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_10_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_10_13_1  (
            .in0(N__42804),
            .in1(N__34728),
            .in2(_gnd_net_),
            .in3(N__32353),
            .lcout(\c0.n8_adj_2205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__5__2187_LC_10_13_2 .C_ON=1'b0;
    defparam \c0.data_out_8__5__2187_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__5__2187_LC_10_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__5__2187_LC_10_13_2  (
            .in0(N__46846),
            .in1(N__38034),
            .in2(_gnd_net_),
            .in3(N__37390),
            .lcout(data_out_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_10_13_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_10_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_10_13_3  (
            .in0(N__42803),
            .in1(N__34336),
            .in2(_gnd_net_),
            .in3(N__36557),
            .lcout(\c0.n8_adj_2232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_10_13_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_10_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_10_13_4  (
            .in0(N__32674),
            .in1(N__37389),
            .in2(_gnd_net_),
            .in3(N__42802),
            .lcout(\c0.n8_adj_2209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15152_3_lut_4_lut_LC_10_13_6 .C_ON=1'b0;
    defparam \c0.tx.i15152_3_lut_4_lut_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15152_3_lut_4_lut_LC_10_13_6 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \c0.tx.i15152_3_lut_4_lut_LC_10_13_6  (
            .in0(N__31379),
            .in1(N__31325),
            .in2(N__31290),
            .in3(N__31207),
            .lcout(n18012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15305_3_lut_LC_10_13_7 .C_ON=1'b0;
    defparam \c0.tx.i15305_3_lut_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15305_3_lut_LC_10_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i15305_3_lut_LC_10_13_7  (
            .in0(N__31155),
            .in1(N__31109),
            .in2(_gnd_net_),
            .in3(N__32646),
            .lcout(\c0.tx.n18166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15948_LC_10_14_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15948_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15948_LC_10_14_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15948_LC_10_14_0  (
            .in0(N__32625),
            .in1(N__35192),
            .in2(N__31563),
            .in3(N__34833),
            .lcout(\c0.n18753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18873_bdd_4_lut_LC_10_14_1 .C_ON=1'b0;
    defparam \c0.n18873_bdd_4_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18873_bdd_4_lut_LC_10_14_1 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18873_bdd_4_lut_LC_10_14_1  (
            .in0(N__35193),
            .in1(N__31548),
            .in2(N__31539),
            .in3(N__31512),
            .lcout(),
            .ltout(n18876_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_819_LC_10_14_2.C_ON=1'b0;
    defparam i24_4_lut_adj_819_LC_10_14_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_819_LC_10_14_2.LUT_INIT=16'b0011000010111000;
    LogicCell40 i24_4_lut_adj_819_LC_10_14_2 (
            .in0(N__31494),
            .in1(N__35080),
            .in2(N__31524),
            .in3(N__35194),
            .lcout(n10_adj_2531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_10_14_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_10_14_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_10_14_3  (
            .in0(N__39941),
            .in1(N__42821),
            .in2(_gnd_net_),
            .in3(N__36745),
            .lcout(),
            .ltout(\c0.n5_adj_2196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_14_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_14_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_14_4  (
            .in0(N__31683),
            .in1(N__35191),
            .in2(N__31515),
            .in3(N__34834),
            .lcout(\c0.n18873 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_10_14_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_10_14_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_10_14_5  (
            .in0(N__36854),
            .in1(N__42820),
            .in2(_gnd_net_),
            .in3(N__34563),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i43_4_lut_LC_10_14_6.C_ON=1'b0;
    defparam i43_4_lut_LC_10_14_6.SEQ_MODE=4'b0000;
    defparam i43_4_lut_LC_10_14_6.LUT_INIT=16'b1111000010001000;
    LogicCell40 i43_4_lut_LC_10_14_6 (
            .in0(N__42822),
            .in1(N__37336),
            .in2(N__31506),
            .in3(N__34832),
            .lcout(n24_adj_2523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_10_14_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_10_14_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_10_14_7  (
            .in0(N__34835),
            .in1(N__42823),
            .in2(N__31503),
            .in3(N__34683),
            .lcout(n10_adj_2533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15533_3_lut_LC_10_15_0 .C_ON=1'b0;
    defparam \c0.i15533_3_lut_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15533_3_lut_LC_10_15_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15533_3_lut_LC_10_15_0  (
            .in0(N__37340),
            .in1(N__47646),
            .in2(_gnd_net_),
            .in3(N__39837),
            .lcout(\c0.n18230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_825_LC_10_15_1.C_ON=1'b0;
    defparam i24_4_lut_adj_825_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_825_LC_10_15_1.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_825_LC_10_15_1 (
            .in0(N__34923),
            .in1(N__35093),
            .in2(N__32370),
            .in3(N__35247),
            .lcout(),
            .ltout(n10_adj_2528_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_10_15_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_15_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_10_15_2  (
            .in0(N__32614),
            .in1(N__31628),
            .in2(N__31635),
            .in3(N__32531),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15731_2_lut_3_lut_LC_10_15_3 .C_ON=1'b0;
    defparam \c0.i15731_2_lut_3_lut_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15731_2_lut_3_lut_LC_10_15_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i15731_2_lut_3_lut_LC_10_15_3  (
            .in0(N__43368),
            .in1(N__47634),
            .in2(_gnd_net_),
            .in3(N__47072),
            .lcout(\c0.n11016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_549_LC_10_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_549_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_549_LC_10_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_549_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__34347),
            .in2(_gnd_net_),
            .in3(N__37284),
            .lcout(\c0.n10558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__5__2227_LC_10_15_5 .C_ON=1'b0;
    defparam \c0.data_out_3__5__2227_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5__2227_LC_10_15_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_3__5__2227_LC_10_15_5  (
            .in0(N__47345),
            .in1(N__43346),
            .in2(N__31614),
            .in3(N__47073),
            .lcout(data_out_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49717),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6__2250_LC_10_16_0 .C_ON=1'b0;
    defparam \c0.data_out_0__6__2250_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__6__2250_LC_10_16_0 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \c0.data_out_0__6__2250_LC_10_16_0  (
            .in0(N__47680),
            .in1(N__47118),
            .in2(N__43393),
            .in3(N__31587),
            .lcout(\c0.data_out_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_16_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_16_2  (
            .in0(N__31598),
            .in1(N__31586),
            .in2(_gnd_net_),
            .in3(N__42810),
            .lcout(\c0.n1_adj_2272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15707_3_lut_LC_10_16_4 .C_ON=1'b0;
    defparam \c0.i15707_3_lut_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15707_3_lut_LC_10_16_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15707_3_lut_LC_10_16_4  (
            .in0(N__47679),
            .in1(N__36891),
            .in2(_gnd_net_),
            .in3(N__37485),
            .lcout(\c0.n18184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15958_LC_10_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15958_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15958_LC_10_16_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15958_LC_10_16_5  (
            .in0(N__32718),
            .in1(N__35195),
            .in2(N__32655),
            .in3(N__34867),
            .lcout(\c0.n18849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15604_2_lut_LC_10_16_6 .C_ON=1'b0;
    defparam \c0.i15604_2_lut_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15604_2_lut_LC_10_16_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i15604_2_lut_LC_10_16_6  (
            .in0(N__31673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42809),
            .lcout(\c0.n18377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__5__2235_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.data_out_2__5__2235_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__5__2235_LC_10_17_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \c0.data_out_2__5__2235_LC_10_17_1  (
            .in0(N__43269),
            .in1(N__47119),
            .in2(_gnd_net_),
            .in3(N__31697),
            .lcout(data_out_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15657_2_lut_LC_10_17_3 .C_ON=1'b0;
    defparam \c0.i15657_2_lut_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15657_2_lut_LC_10_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15657_2_lut_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__37484),
            .in2(_gnd_net_),
            .in3(N__42712),
            .lcout(\c0.n18335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3__2237_LC_10_17_7 .C_ON=1'b0;
    defparam \c0.data_out_2__3__2237_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__3__2237_LC_10_17_7 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \c0.data_out_2__3__2237_LC_10_17_7  (
            .in0(N__47678),
            .in1(N__31674),
            .in2(N__43318),
            .in3(N__47120),
            .lcout(\c0.data_out_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15068_2_lut_LC_10_27_4 .C_ON=1'b0;
    defparam \control.i15068_2_lut_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \control.i15068_2_lut_LC_10_27_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \control.i15068_2_lut_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__35574),
            .in2(_gnd_net_),
            .in3(N__35665),
            .lcout(\control.n17926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15091_2_lut_LC_10_29_7 .C_ON=1'b0;
    defparam \control.i15091_2_lut_LC_10_29_7 .SEQ_MODE=4'b0000;
    defparam \control.i15091_2_lut_LC_10_29_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \control.i15091_2_lut_LC_10_29_7  (
            .in0(_gnd_net_),
            .in1(N__35575),
            .in2(_gnd_net_),
            .in3(N__32921),
            .lcout(\control.n17950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_11_1_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_11_1_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_11_1_0  (
            .in0(N__37859),
            .in1(N__37653),
            .in2(N__40406),
            .in3(N__33332),
            .lcout(),
            .ltout(\c0.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i154_LC_11_1_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i154_LC_11_1_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i154_LC_11_1_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_frame2_0___i154_LC_11_1_1  (
            .in0(N__32964),
            .in1(_gnd_net_),
            .in2(N__31662),
            .in3(N__31650),
            .lcout(\c0.data_out_frame2_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__50444),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_11_1_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_11_1_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_11_1_2  (
            .in0(N__41724),
            .in1(N__40791),
            .in2(N__36012),
            .in3(N__45455),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15649_3_lut_LC_11_1_3 .C_ON=1'b0;
    defparam \c0.i15649_3_lut_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15649_3_lut_LC_11_1_3 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \c0.i15649_3_lut_LC_11_1_3  (
            .in0(_gnd_net_),
            .in1(N__46205),
            .in2(N__48682),
            .in3(N__37858),
            .lcout(\c0.n18266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15206_3_lut_LC_11_1_4 .C_ON=1'b0;
    defparam \c0.i15206_3_lut_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15206_3_lut_LC_11_1_4 .LUT_INIT=16'b1100001011000010;
    LogicCell40 \c0.i15206_3_lut_LC_11_1_4  (
            .in0(N__37740),
            .in1(N__48591),
            .in2(N__46210),
            .in3(_gnd_net_),
            .lcout(\c0.n18067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15557_2_lut_3_lut_LC_11_1_5 .C_ON=1'b0;
    defparam \c0.i15557_2_lut_3_lut_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15557_2_lut_3_lut_LC_11_1_5 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \c0.i15557_2_lut_3_lut_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__46201),
            .in2(N__48681),
            .in3(N__50671),
            .lcout(\c0.n18221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15606_3_lut_LC_11_1_6 .C_ON=1'b0;
    defparam \c0.i15606_3_lut_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15606_3_lut_LC_11_1_6 .LUT_INIT=16'b0011001000110010;
    LogicCell40 \c0.i15606_3_lut_LC_11_1_6  (
            .in0(N__44374),
            .in1(N__48595),
            .in2(N__46211),
            .in3(_gnd_net_),
            .lcout(\c0.n18360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15608_3_lut_LC_11_1_7 .C_ON=1'b0;
    defparam \c0.i15608_3_lut_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15608_3_lut_LC_11_1_7 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \c0.i15608_3_lut_LC_11_1_7  (
            .in0(_gnd_net_),
            .in1(N__46206),
            .in2(N__48683),
            .in3(N__40468),
            .lcout(\c0.n18256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_11_2_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_11_2_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_11_2_0  (
            .in0(N__40940),
            .in1(N__40983),
            .in2(N__44172),
            .in3(N__37559),
            .lcout(),
            .ltout(\c0.n14_adj_2359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i161_LC_11_2_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i161_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i161_LC_11_2_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i161_LC_11_2_1  (
            .in0(N__31704),
            .in1(N__31710),
            .in2(N__31719),
            .in3(N__37761),
            .lcout(\c0.data_out_frame2_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49868),
            .ce(N__50426),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_721_LC_11_2_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_721_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_721_LC_11_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_721_LC_11_2_2  (
            .in0(N__44973),
            .in1(N__46262),
            .in2(N__44589),
            .in3(N__45669),
            .lcout(\c0.n15_adj_2429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_527_LC_11_2_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_527_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_527_LC_11_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_527_LC_11_2_3  (
            .in0(N__44286),
            .in1(N__43819),
            .in2(_gnd_net_),
            .in3(N__43865),
            .lcout(\c0.n17847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_798_LC_11_2_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_798_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_798_LC_11_2_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_798_LC_11_2_4  (
            .in0(N__43818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33324),
            .lcout(\c0.n10867 ),
            .ltout(\c0.n10867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_806_LC_11_2_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_806_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_806_LC_11_2_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_806_LC_11_2_5  (
            .in0(N__33644),
            .in1(N__36153),
            .in2(N__31791),
            .in3(N__45696),
            .lcout(\c0.n17_adj_2449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i59_LC_11_3_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i59_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i59_LC_11_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i59_LC_11_3_0  (
            .in0(N__50263),
            .in1(N__38568),
            .in2(_gnd_net_),
            .in3(N__50742),
            .lcout(data_out_frame2_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_789_LC_11_3_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_789_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_789_LC_11_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_789_LC_11_3_1  (
            .in0(N__46638),
            .in1(N__43745),
            .in2(_gnd_net_),
            .in3(N__50703),
            .lcout(),
            .ltout(\c0.n17739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_709_LC_11_3_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_709_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_709_LC_11_3_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_709_LC_11_3_2  (
            .in0(N__31866),
            .in1(N__44659),
            .in2(N__31788),
            .in3(N__43892),
            .lcout(\c0.n28_adj_2425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i137_LC_11_3_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i137_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i137_LC_11_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i137_LC_11_3_3  (
            .in0(N__38720),
            .in1(N__31784),
            .in2(_gnd_net_),
            .in3(N__50261),
            .lcout(data_out_frame2_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18837_bdd_4_lut_LC_11_3_4 .C_ON=1'b0;
    defparam \c0.n18837_bdd_4_lut_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18837_bdd_4_lut_LC_11_3_4 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18837_bdd_4_lut_LC_11_3_4  (
            .in0(N__48487),
            .in1(N__31833),
            .in2(N__31785),
            .in3(N__37188),
            .lcout(\c0.n18840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i136_LC_11_3_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i136_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i136_LC_11_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i136_LC_11_3_5  (
            .in0(N__42098),
            .in1(N__40984),
            .in2(_gnd_net_),
            .in3(N__50260),
            .lcout(data_out_frame2_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15909_LC_11_3_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15909_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15909_LC_11_3_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15909_LC_11_3_6  (
            .in0(N__35985),
            .in1(N__40389),
            .in2(N__48606),
            .in3(N__46190),
            .lcout(\c0.n18795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i152_LC_11_3_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i152_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i152_LC_11_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i152_LC_11_3_7  (
            .in0(N__42099),
            .in1(N__31757),
            .in2(_gnd_net_),
            .in3(N__50262),
            .lcout(data_out_frame2_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i88_LC_11_4_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i88_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i88_LC_11_4_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i88_LC_11_4_0  (
            .in0(N__50137),
            .in1(_gnd_net_),
            .in2(N__39633),
            .in3(N__44749),
            .lcout(data_out_frame2_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i42_LC_11_4_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i42_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i42_LC_11_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i42_LC_11_4_1  (
            .in0(N__39503),
            .in1(N__31855),
            .in2(_gnd_net_),
            .in3(N__50134),
            .lcout(data_out_frame2_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i54_LC_11_4_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i54_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i54_LC_11_4_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i54_LC_11_4_2  (
            .in0(N__50135),
            .in1(N__38846),
            .in2(_gnd_net_),
            .in3(N__44888),
            .lcout(data_out_frame2_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i114_LC_11_4_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i114_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i114_LC_11_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i114_LC_11_4_3  (
            .in0(N__39087),
            .in1(N__40396),
            .in2(_gnd_net_),
            .in3(N__50131),
            .lcout(data_out_frame2_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15953_LC_11_4_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15953_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15953_LC_11_4_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15953_LC_11_4_4  (
            .in0(N__46185),
            .in1(N__48524),
            .in2(N__37602),
            .in3(N__33344),
            .lcout(\c0.n18837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i83_LC_11_4_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i83_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i83_LC_11_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i83_LC_11_4_5  (
            .in0(N__40891),
            .in1(N__36183),
            .in2(_gnd_net_),
            .in3(N__50136),
            .lcout(data_out_frame2_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i146_LC_11_4_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i146_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i146_LC_11_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i146_LC_11_4_6  (
            .in0(N__50133),
            .in1(N__38336),
            .in2(_gnd_net_),
            .in3(N__31823),
            .lcout(data_out_frame2_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i144_LC_11_4_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i144_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i144_LC_11_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i144_LC_11_4_7  (
            .in0(N__39232),
            .in1(N__31805),
            .in2(_gnd_net_),
            .in3(N__50132),
            .lcout(data_out_frame2_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i50_LC_11_5_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i50_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i50_LC_11_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i50_LC_11_5_0  (
            .in0(N__50254),
            .in1(N__39085),
            .in2(_gnd_net_),
            .in3(N__44040),
            .lcout(data_out_frame2_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i84_LC_11_5_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i84_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i84_LC_11_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i84_LC_11_5_2  (
            .in0(N__50256),
            .in1(N__38982),
            .in2(_gnd_net_),
            .in3(N__41406),
            .lcout(data_out_frame2_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i99_LC_11_5_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i99_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i99_LC_11_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i99_LC_11_5_3  (
            .in0(N__38271),
            .in1(N__41076),
            .in2(_gnd_net_),
            .in3(N__50259),
            .lcout(data_out_frame2_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i96_LC_11_5_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i96_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i96_LC_11_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i96_LC_11_5_4  (
            .in0(N__50258),
            .in1(N__39234),
            .in2(_gnd_net_),
            .in3(N__43660),
            .lcout(data_out_frame2_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i128_LC_11_5_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i128_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i128_LC_11_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i128_LC_11_5_5  (
            .in0(N__39233),
            .in1(N__40928),
            .in2(_gnd_net_),
            .in3(N__50253),
            .lcout(data_out_frame2_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i53_LC_11_5_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i53_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i53_LC_11_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i53_LC_11_5_6  (
            .in0(N__50255),
            .in1(N__38907),
            .in2(_gnd_net_),
            .in3(N__36220),
            .lcout(data_out_frame2_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i87_LC_11_5_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i87_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i87_LC_11_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i87_LC_11_5_7  (
            .in0(N__39705),
            .in1(N__50789),
            .in2(_gnd_net_),
            .in3(N__50257),
            .lcout(data_out_frame2_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_682_LC_11_6_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_682_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_682_LC_11_6_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_682_LC_11_6_0  (
            .in0(N__41624),
            .in1(N__44967),
            .in2(N__36363),
            .in3(N__37128),
            .lcout(\c0.n16_adj_2412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_479_LC_11_6_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_479_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_479_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_479_LC_11_6_1  (
            .in0(N__45789),
            .in1(N__43655),
            .in2(_gnd_net_),
            .in3(N__40739),
            .lcout(\c0.n17727 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i110_LC_11_6_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i110_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i110_LC_11_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i110_LC_11_6_2  (
            .in0(N__50313),
            .in1(N__39343),
            .in2(_gnd_net_),
            .in3(N__44792),
            .lcout(data_out_frame2_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i151_LC_11_6_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i151_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i151_LC_11_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i151_LC_11_6_4  (
            .in0(N__50314),
            .in1(N__41284),
            .in2(_gnd_net_),
            .in3(N__42368),
            .lcout(data_out_frame2_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_11_6_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_11_6_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_11_6_5  (
            .in0(N__36216),
            .in1(_gnd_net_),
            .in2(N__44972),
            .in3(N__46139),
            .lcout(\c0.n5_adj_2436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i82_LC_11_6_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i82_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i82_LC_11_6_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i82_LC_11_6_6  (
            .in0(N__50316),
            .in1(_gnd_net_),
            .in2(N__40750),
            .in3(N__39086),
            .lcout(data_out_frame2_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i58_LC_11_6_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i58_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i58_LC_11_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i58_LC_11_6_7  (
            .in0(N__38650),
            .in1(N__31903),
            .in2(_gnd_net_),
            .in3(N__50315),
            .lcout(data_out_frame2_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i0_LC_11_7_0 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i0_LC_11_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__32097),
            .in2(N__33573),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\c0.n16634 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i1_LC_11_7_1 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i1_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i1_LC_11_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__33420),
            .in2(_gnd_net_),
            .in3(N__31884),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n16634 ),
            .carryout(\c0.n16635 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i2_LC_11_7_2 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i2_LC_11_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__31952),
            .in2(_gnd_net_),
            .in3(N__31881),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n16635 ),
            .carryout(\c0.n16636 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i3_LC_11_7_3 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i3_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i3_LC_11_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__33617),
            .in2(_gnd_net_),
            .in3(N__31878),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n16636 ),
            .carryout(\c0.n16637 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i4_LC_11_7_4 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i4_LC_11_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__32060),
            .in2(_gnd_net_),
            .in3(N__31875),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n16637 ),
            .carryout(\c0.n16638 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i5_LC_11_7_5 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i5_LC_11_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__31934),
            .in2(_gnd_net_),
            .in3(N__31872),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n16638 ),
            .carryout(\c0.n16639 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i6_LC_11_7_6 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i6_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i6_LC_11_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__33543),
            .in2(_gnd_net_),
            .in3(N__31869),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n16639 ),
            .carryout(\c0.n16640 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i7_LC_11_7_7 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i7_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i7_LC_11_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__32045),
            .in2(_gnd_net_),
            .in3(N__31974),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(\c0.n16640 ),
            .carryout(\c0.n16641 ),
            .clk(N__49829),
            .ce(N__36516),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i8_LC_11_8_0 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i8_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i8_LC_11_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i8_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__33603),
            .in2(_gnd_net_),
            .in3(N__31971),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\c0.n16642 ),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i9_LC_11_8_1 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i9_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i9_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i9_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__33432),
            .in2(_gnd_net_),
            .in3(N__31968),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(\c0.n16642 ),
            .carryout(\c0.n16643 ),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i10_LC_11_8_2 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i10_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i10_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i10_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__33585),
            .in2(_gnd_net_),
            .in3(N__31965),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(\c0.n16643 ),
            .carryout(\c0.n16644 ),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i11_LC_11_8_3 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i11_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i11_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i11_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__32088),
            .in2(_gnd_net_),
            .in3(N__31962),
            .lcout(\c0.delay_counter_11 ),
            .ltout(),
            .carryin(\c0.n16644 ),
            .carryout(\c0.n16645 ),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i12_LC_11_8_4 .C_ON=1'b1;
    defparam \c0.delay_counter_2484__i12_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i12_LC_11_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i12_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__32076),
            .in2(_gnd_net_),
            .in3(N__31959),
            .lcout(\c0.delay_counter_12 ),
            .ltout(),
            .carryin(\c0.n16645 ),
            .carryout(\c0.n16646 ),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2484__i13_LC_11_8_5 .C_ON=1'b0;
    defparam \c0.delay_counter_2484__i13_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2484__i13_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2484__i13_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__33557),
            .in2(_gnd_net_),
            .in3(N__31956),
            .lcout(\c0.delay_counter_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49816),
            .ce(N__36512),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_11_9_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_11_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_LC_11_9_0  (
            .in0(N__31953),
            .in1(N__33591),
            .in2(N__31938),
            .in3(N__32031),
            .lcout(n26_adj_2466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_438_LC_11_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_438_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_438_LC_11_9_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_438_LC_11_9_1  (
            .in0(N__33789),
            .in1(N__32023),
            .in2(_gnd_net_),
            .in3(N__33851),
            .lcout(\c0.n98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15158_4_lut_LC_11_9_2 .C_ON=1'b0;
    defparam \c0.i15158_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15158_4_lut_LC_11_9_2 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \c0.i15158_4_lut_LC_11_9_2  (
            .in0(N__33852),
            .in1(N__33446),
            .in2(N__47128),
            .in3(N__33790),
            .lcout(\c0.n18019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_441_LC_11_9_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_441_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_441_LC_11_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_441_LC_11_9_3  (
            .in0(N__33788),
            .in1(N__33850),
            .in2(_gnd_net_),
            .in3(N__33806),
            .lcout(n129),
            .ltout(n129_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_567_LC_11_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_567_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_567_LC_11_9_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_567_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__32168),
            .in2(N__32139),
            .in3(N__32136),
            .lcout(\c0.n1707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_11_9_5 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_11_9_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_LC_11_9_5  (
            .in0(N__32087),
            .in1(N__32075),
            .in2(N__32064),
            .in3(N__32046),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_11_9_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_11_9_6 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_11_9_6  (
            .in0(N__33853),
            .in1(N__33445),
            .in2(N__32025),
            .in3(N__33787),
            .lcout(n574),
            .ltout(n574_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_618_LC_11_9_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_618_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_618_LC_11_9_7 .LUT_INIT=16'b0001000011011100;
    LogicCell40 \c0.i1_4_lut_adj_618_LC_11_9_7  (
            .in0(N__47258),
            .in1(N__47085),
            .in2(N__31998),
            .in3(N__31995),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3__2205_LC_11_10_0 .C_ON=1'b0;
    defparam \c0.data_out_6__3__2205_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3__2205_LC_11_10_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__3__2205_LC_11_10_0  (
            .in0(N__38931),
            .in1(N__47237),
            .in2(N__31989),
            .in3(N__46974),
            .lcout(\c0.data_out_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49793),
            .ce(N__43425),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2__2206_LC_11_10_1 .C_ON=1'b0;
    defparam \c0.data_out_6__2__2206_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2__2206_LC_11_10_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_6__2__2206_LC_11_10_1  (
            .in0(N__46973),
            .in1(N__39006),
            .in2(N__32235),
            .in3(N__47255),
            .lcout(\c0.data_out_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49793),
            .ce(N__43425),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_587_LC_11_10_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_587_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_587_LC_11_10_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_587_LC_11_10_2  (
            .in0(N__47254),
            .in1(N__46970),
            .in2(_gnd_net_),
            .in3(N__32295),
            .lcout(n6_adj_2470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15119_2_lut_3_lut_LC_11_10_3.C_ON=1'b0;
    defparam i15119_2_lut_3_lut_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam i15119_2_lut_3_lut_LC_11_10_3.LUT_INIT=16'b1111111111101110;
    LogicCell40 i15119_2_lut_3_lut_LC_11_10_3 (
            .in0(N__46968),
            .in1(N__32270),
            .in2(_gnd_net_),
            .in3(N__32256),
            .lcout(),
            .ltout(n17978_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15531_4_lut_LC_11_10_4.C_ON=1'b0;
    defparam i15531_4_lut_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam i15531_4_lut_LC_11_10_4.LUT_INIT=16'b0101111100011111;
    LogicCell40 i15531_4_lut_LC_11_10_4 (
            .in0(N__47550),
            .in1(N__46971),
            .in2(N__32298),
            .in3(N__32294),
            .lcout(n18202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15708_4_lut_LC_11_10_6.C_ON=1'b0;
    defparam i15708_4_lut_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam i15708_4_lut_LC_11_10_6.LUT_INIT=16'b0001000100010000;
    LogicCell40 i15708_4_lut_LC_11_10_6 (
            .in0(N__32258),
            .in1(N__47236),
            .in2(N__32274),
            .in3(N__46972),
            .lcout(n18368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_11_10_7.C_ON=1'b0;
    defparam i1_2_lut_LC_11_10_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_11_10_7.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_LC_11_10_7 (
            .in0(N__46969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32257),
            .lcout(n22_adj_2522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15560_3_lut_LC_11_11_0 .C_ON=1'b0;
    defparam \c0.i15560_3_lut_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15560_3_lut_LC_11_11_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15560_3_lut_LC_11_11_0  (
            .in0(N__47549),
            .in1(N__42493),
            .in2(_gnd_net_),
            .in3(N__37341),
            .lcout(\c0.n18226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i42_4_lut_LC_11_11_2.C_ON=1'b0;
    defparam i42_4_lut_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam i42_4_lut_LC_11_11_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 i42_4_lut_LC_11_11_2 (
            .in0(N__33957),
            .in1(N__35072),
            .in2(N__32769),
            .in3(N__35218),
            .lcout(n21_adj_2524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i3_LC_11_11_3 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i3_LC_11_11_3 .LUT_INIT=16'b0001000010111010;
    LogicCell40 \c0.UART_TRANSMITTER_state__i3_LC_11_11_3  (
            .in0(N__47554),
            .in1(N__32220),
            .in2(N__47798),
            .in3(N__32214),
            .lcout(UART_TRANSMITTER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15963_LC_11_11_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15963_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15963_LC_11_11_4 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15963_LC_11_11_4  (
            .in0(N__34008),
            .in1(N__34852),
            .in2(N__42561),
            .in3(N__35216),
            .lcout(),
            .ltout(\c0.n18861_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18861_bdd_4_lut_LC_11_11_5 .C_ON=1'b0;
    defparam \c0.n18861_bdd_4_lut_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18861_bdd_4_lut_LC_11_11_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18861_bdd_4_lut_LC_11_11_5  (
            .in0(N__35217),
            .in1(N__36570),
            .in2(N__32208),
            .in3(N__32205),
            .lcout(),
            .ltout(n18864_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_823_LC_11_11_6.C_ON=1'b0;
    defparam i24_4_lut_adj_823_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_823_LC_11_11_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 i24_4_lut_adj_823_LC_11_11_6 (
            .in0(N__32307),
            .in1(N__35073),
            .in2(N__32328),
            .in3(N__35219),
            .lcout(),
            .ltout(n10_adj_2529_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_11_11_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_11_11_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_11_11_7  (
            .in0(N__32601),
            .in1(N__32321),
            .in2(N__32325),
            .in3(N__32513),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_496_LC_11_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_496_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_496_LC_11_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_496_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__34701),
            .in2(_gnd_net_),
            .in3(N__32424),
            .lcout(\c0.n17850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_11_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_11_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_727_LC_11_12_1  (
            .in0(N__34679),
            .in1(N__34593),
            .in2(N__37368),
            .in3(N__42494),
            .lcout(\c0.n6_adj_2276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_11_12_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_11_12_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_11_12_3  (
            .in0(N__34699),
            .in1(N__34851),
            .in2(N__36603),
            .in3(N__42780),
            .lcout(n10_adj_2499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_543_LC_11_12_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_543_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_543_LC_11_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_543_LC_11_12_4  (
            .in0(N__39834),
            .in1(N__36858),
            .in2(N__34525),
            .in3(N__36777),
            .lcout(\c0.n10550 ),
            .ltout(\c0.n10550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_712_LC_11_12_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_712_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_712_LC_11_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_712_LC_11_12_5  (
            .in0(N__34700),
            .in1(N__32682),
            .in2(N__32301),
            .in3(N__32438),
            .lcout(\c0.n14_adj_2320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_540_LC_11_12_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_540_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_540_LC_11_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_540_LC_11_12_6  (
            .in0(N__34592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34678),
            .lcout(\c0.n10524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_11_12_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_11_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_11_12_7  (
            .in0(N__32712),
            .in1(N__43437),
            .in2(_gnd_net_),
            .in3(N__42779),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_545_LC_11_13_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_545_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_545_LC_11_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_545_LC_11_13_0  (
            .in0(N__34494),
            .in1(N__32439),
            .in2(N__36659),
            .in3(N__32423),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_537_LC_11_13_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_537_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_537_LC_11_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_537_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__34408),
            .in2(_gnd_net_),
            .in3(N__43148),
            .lcout(\c0.n6_adj_2361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_531_LC_11_13_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_531_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_531_LC_11_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_531_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__36462),
            .in2(_gnd_net_),
            .in3(N__36709),
            .lcout(\c0.n10746 ),
            .ltout(\c0.n10746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_538_LC_11_13_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_538_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_538_LC_11_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_538_LC_11_13_4  (
            .in0(N__32397),
            .in1(N__32385),
            .in2(N__32391),
            .in3(N__34439),
            .lcout(n17758),
            .ltout(n17758_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__2__2182_LC_11_13_5 .C_ON=1'b0;
    defparam \c0.data_out_9__2__2182_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__2__2182_LC_11_13_5 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \c0.data_out_9__2__2182_LC_11_13_5  (
            .in0(N__46853),
            .in1(N__34343),
            .in2(N__32388),
            .in3(N__37097),
            .lcout(data_out_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49752),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_666_LC_11_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_666_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_666_LC_11_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_666_LC_11_13_6  (
            .in0(N__37442),
            .in1(N__37388),
            .in2(_gnd_net_),
            .in3(N__42469),
            .lcout(\c0.n10734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_11_13_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_11_13_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_11_13_7  (
            .in0(N__34409),
            .in1(N__34871),
            .in2(N__32379),
            .in3(N__42830),
            .lcout(n10_adj_2461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_487_LC_11_14_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_487_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_487_LC_11_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_487_LC_11_14_1  (
            .in0(N__34533),
            .in1(N__39751),
            .in2(N__37047),
            .in3(N__32358),
            .lcout(\c0.n17742 ),
            .ltout(\c0.n17742_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__4__2180_LC_11_14_2 .C_ON=1'b0;
    defparam \c0.data_out_9__4__2180_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__4__2180_LC_11_14_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__4__2180_LC_11_14_2  (
            .in0(N__34962),
            .in1(N__36485),
            .in2(N__32331),
            .in3(N__43152),
            .lcout(\c0.data_out_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49739),
            .ce(N__46854),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__5__2179_LC_11_14_4 .C_ON=1'b0;
    defparam \c0.data_out_9__5__2179_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__5__2179_LC_11_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__5__2179_LC_11_14_4  (
            .in0(N__32697),
            .in1(N__34656),
            .in2(N__32691),
            .in3(N__42540),
            .lcout(\c0.data_out_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49739),
            .ce(N__46854),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_11_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_621_LC_11_14_5  (
            .in0(N__34337),
            .in1(N__39750),
            .in2(_gnd_net_),
            .in3(N__37282),
            .lcout(),
            .ltout(\c0.n6_adj_2365_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_551_LC_11_14_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_551_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_551_LC_11_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_551_LC_11_14_6  (
            .in0(N__34968),
            .in1(N__42937),
            .in2(N__32658),
            .in3(N__36746),
            .lcout(\c0.n17768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_11_15_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_11_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_11_15_0  (
            .in0(N__37537),
            .in1(N__43147),
            .in2(_gnd_net_),
            .in3(N__42817),
            .lcout(\c0.n5_adj_2220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_15_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_15_1  (
            .in0(N__42818),
            .in1(N__50924),
            .in2(_gnd_net_),
            .in3(N__34532),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_11_15_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_15_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_11_15_2  (
            .in0(N__32525),
            .in1(N__32618),
            .in2(N__32645),
            .in3(N__35019),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_579_LC_11_15_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_579_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_579_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_579_LC_11_15_3  (
            .in0(N__39984),
            .in1(N__50925),
            .in2(_gnd_net_),
            .in3(N__39893),
            .lcout(\c0.n10537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15584_2_lut_LC_11_15_4 .C_ON=1'b0;
    defparam \c0.i15584_2_lut_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15584_2_lut_LC_11_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15584_2_lut_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__43527),
            .in2(_gnd_net_),
            .in3(N__42816),
            .lcout(\c0.n18265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_11_15_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_11_15_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_11_15_5  (
            .in0(N__32453),
            .in1(N__32748),
            .in2(N__32619),
            .in3(N__32535),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10351_3_lut_LC_11_15_6 .C_ON=1'b0;
    defparam \c0.i10351_3_lut_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10351_3_lut_LC_11_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i10351_3_lut_LC_11_15_6  (
            .in0(N__34590),
            .in1(N__39985),
            .in2(_gnd_net_),
            .in3(N__34857),
            .lcout(),
            .ltout(\c0.n1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_LC_11_15_7 .C_ON=1'b0;
    defparam \c0.i29_4_lut_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_LC_11_15_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.i29_4_lut_LC_11_15_7  (
            .in0(N__42819),
            .in1(N__34858),
            .in2(N__32772),
            .in3(N__37043),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18849_bdd_4_lut_LC_11_16_0 .C_ON=1'b0;
    defparam \c0.n18849_bdd_4_lut_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18849_bdd_4_lut_LC_11_16_0 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18849_bdd_4_lut_LC_11_16_0  (
            .in0(N__40236),
            .in1(N__32757),
            .in2(N__32742),
            .in3(N__35234),
            .lcout(),
            .ltout(n18852_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_11_16_1.C_ON=1'b0;
    defparam i24_4_lut_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_11_16_1.LUT_INIT=16'b0100010011110000;
    LogicCell40 i24_4_lut_LC_11_16_1 (
            .in0(N__35235),
            .in1(N__32724),
            .in2(N__32751),
            .in3(N__35088),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15580_2_lut_LC_11_16_2 .C_ON=1'b0;
    defparam \c0.i15580_2_lut_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15580_2_lut_LC_11_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15580_2_lut_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__32945),
            .in2(_gnd_net_),
            .in3(N__42814),
            .lcout(\c0.n18264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_11_16_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_11_16_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_11_16_3  (
            .in0(N__42815),
            .in1(N__34632),
            .in2(N__32733),
            .in3(N__34878),
            .lcout(n10_adj_2527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__4__2244_LC_11_16_5 .C_ON=1'b0;
    defparam \c0.data_out_1__4__2244_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__4__2244_LC_11_16_5 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \c0.data_out_1__4__2244_LC_11_16_5  (
            .in0(N__47632),
            .in1(N__47081),
            .in2(N__43317),
            .in3(N__35003),
            .lcout(\c0.data_out_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49718),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15643_2_lut_LC_11_16_6 .C_ON=1'b0;
    defparam \c0.i15643_2_lut_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15643_2_lut_LC_11_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15643_2_lut_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__42485),
            .in2(_gnd_net_),
            .in3(N__42813),
            .lcout(\c0.n18322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__1__2255_LC_11_16_7 .C_ON=1'b0;
    defparam \c0.data_out_0__1__2255_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__1__2255_LC_11_16_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \c0.data_out_0__1__2255_LC_11_16_7  (
            .in0(N__43260),
            .in1(N__47080),
            .in2(_gnd_net_),
            .in3(N__32711),
            .lcout(data_out_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49718),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15737_4_lut_4_lut_4_lut_3_lut_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.i15737_4_lut_4_lut_4_lut_3_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15737_4_lut_4_lut_4_lut_3_lut_LC_11_17_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \c0.i15737_4_lut_4_lut_4_lut_3_lut_LC_11_17_6  (
            .in0(N__47625),
            .in1(N__47320),
            .in2(_gnd_net_),
            .in3(N__47070),
            .lcout(n11017),
            .ltout(n11017_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__0__2256_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.data_out_0__0__2256_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0__2256_LC_11_17_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.data_out_0__0__2256_LC_11_17_7  (
            .in0(N__47071),
            .in1(N__32946),
            .in2(N__32949),
            .in3(N__47346),
            .lcout(data_out_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49705),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__4__2228_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.data_out_3__4__2228_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4__2228_LC_11_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_3__4__2228_LC_11_18_2  (
            .in0(N__32934),
            .in1(N__40277),
            .in2(_gnd_net_),
            .in3(N__43270),
            .lcout(data_out_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49719),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15603_2_lut_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.i15603_2_lut_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15603_2_lut_LC_11_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15603_2_lut_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__32933),
            .in2(_gnd_net_),
            .in3(N__42861),
            .lcout(\c0.n18191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i1_2_lut_4_lut_adj_814_LC_11_27_4 .C_ON=1'b0;
    defparam \control.i1_2_lut_4_lut_adj_814_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \control.i1_2_lut_4_lut_adj_814_LC_11_27_4 .LUT_INIT=16'b0011101111111111;
    LogicCell40 \control.i1_2_lut_4_lut_adj_814_LC_11_27_4  (
            .in0(N__35679),
            .in1(N__32905),
            .in2(N__35471),
            .in3(N__32857),
            .lcout(\control.n17251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i1_3_lut_LC_11_28_1 .C_ON=1'b0;
    defparam \control.i1_3_lut_LC_11_28_1 .SEQ_MODE=4'b0000;
    defparam \control.i1_3_lut_LC_11_28_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \control.i1_3_lut_LC_11_28_1  (
            .in0(N__35567),
            .in1(N__32925),
            .in2(_gnd_net_),
            .in3(N__35315),
            .lcout(\control.n10490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15757_2_lut_LC_11_28_5 .C_ON=1'b0;
    defparam \control.i15757_2_lut_LC_11_28_5 .SEQ_MODE=4'b0000;
    defparam \control.i15757_2_lut_LC_11_28_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \control.i15757_2_lut_LC_11_28_5  (
            .in0(_gnd_net_),
            .in1(N__32904),
            .in2(_gnd_net_),
            .in3(N__32856),
            .lcout(\control.PHASES_5__N_2160 ),
            .ltout(\control.PHASES_5__N_2160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15769_4_lut_LC_11_28_6 .C_ON=1'b0;
    defparam \control.i15769_4_lut_LC_11_28_6 .SEQ_MODE=4'b0000;
    defparam \control.i15769_4_lut_LC_11_28_6 .LUT_INIT=16'b1111010011111110;
    LogicCell40 \control.i15769_4_lut_LC_11_28_6  (
            .in0(N__35463),
            .in1(N__32823),
            .in2(N__32817),
            .in3(N__32813),
            .lcout(\control.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i1_2_lut_LC_11_28_7 .C_ON=1'b0;
    defparam \control.i1_2_lut_LC_11_28_7 .SEQ_MODE=4'b0000;
    defparam \control.i1_2_lut_LC_11_28_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \control.i1_2_lut_LC_11_28_7  (
            .in0(N__35690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35566),
            .lcout(\control.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.i15762_4_lut_LC_11_29_0 .C_ON=1'b0;
    defparam \control.i15762_4_lut_LC_11_29_0 .SEQ_MODE=4'b0000;
    defparam \control.i15762_4_lut_LC_11_29_0 .LUT_INIT=16'b1111111101110010;
    LogicCell40 \control.i15762_4_lut_LC_11_29_0  (
            .in0(N__35462),
            .in1(N__32814),
            .in2(N__32802),
            .in3(N__35324),
            .lcout(\control.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i57_LC_12_1_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i57_LC_12_1_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i57_LC_12_1_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i57_LC_12_1_0  (
            .in0(N__50425),
            .in1(_gnd_net_),
            .in2(N__38724),
            .in3(N__40536),
            .lcout(data_out_frame2_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i122_LC_12_1_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i122_LC_12_1_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i122_LC_12_1_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i122_LC_12_1_1  (
            .in0(N__38661),
            .in1(N__35980),
            .in2(_gnd_net_),
            .in3(N__50423),
            .lcout(data_out_frame2_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i130_LC_12_1_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i130_LC_12_1_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i130_LC_12_1_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i130_LC_12_1_2  (
            .in0(N__50424),
            .in1(N__38340),
            .in2(_gnd_net_),
            .in3(N__35898),
            .lcout(data_out_frame2_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15784_LC_12_1_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15784_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15784_LC_12_1_3 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15784_LC_12_1_3  (
            .in0(N__48488),
            .in1(N__50711),
            .in2(N__50621),
            .in3(N__46197),
            .lcout(),
            .ltout(\c0.n18639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18639_bdd_4_lut_LC_12_1_4 .C_ON=1'b0;
    defparam \c0.n18639_bdd_4_lut_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18639_bdd_4_lut_LC_12_1_4 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18639_bdd_4_lut_LC_12_1_4  (
            .in0(N__37221),
            .in1(N__41089),
            .in2(N__32970),
            .in3(N__48489),
            .lcout(\c0.n18642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_689_LC_12_1_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_689_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_689_LC_12_1_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_689_LC_12_1_5  (
            .in0(_gnd_net_),
            .in1(N__35979),
            .in2(_gnd_net_),
            .in3(N__44853),
            .lcout(\c0.n10700 ),
            .ltout(\c0.n10700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_535_LC_12_1_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_535_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_535_LC_12_1_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_535_LC_12_1_6  (
            .in0(N__42054),
            .in1(N__43950),
            .in2(N__32967),
            .in3(N__35897),
            .lcout(\c0.n17841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_12_1_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_12_1_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_12_1_7  (
            .in0(N__33030),
            .in1(N__33645),
            .in2(N__32958),
            .in3(N__33024),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_12_2_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_12_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__46261),
            .in2(_gnd_net_),
            .in3(N__37183),
            .lcout(\c0.n17804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_710_LC_12_2_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_710_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_710_LC_12_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_710_LC_12_2_2  (
            .in0(N__36104),
            .in1(N__40355),
            .in2(N__37622),
            .in3(N__45146),
            .lcout(\c0.n29_adj_2427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_432_LC_12_2_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_432_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_432_LC_12_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_432_LC_12_2_3  (
            .in0(N__36184),
            .in1(N__33320),
            .in2(_gnd_net_),
            .in3(N__48220),
            .lcout(\c0.n10849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_426_LC_12_2_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_426_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_426_LC_12_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_426_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(N__44898),
            .in2(_gnd_net_),
            .in3(N__41415),
            .lcout(\c0.n17874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_757_LC_12_2_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_757_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_757_LC_12_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_757_LC_12_2_5  (
            .in0(N__45627),
            .in1(N__44457),
            .in2(_gnd_net_),
            .in3(N__45695),
            .lcout(\c0.n17908 ),
            .ltout(\c0.n17908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_706_LC_12_2_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_706_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_706_LC_12_2_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_706_LC_12_2_6  (
            .in0(N__33018),
            .in1(N__45486),
            .in2(N__33009),
            .in3(N__44490),
            .lcout(),
            .ltout(\c0.n30_adj_2424_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_717_LC_12_2_7 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_717_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_717_LC_12_2_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_717_LC_12_2_7  (
            .in0(N__36387),
            .in1(N__33006),
            .in2(N__33000),
            .in3(N__32997),
            .lcout(\c0.n10577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i62_LC_12_3_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i62_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i62_LC_12_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i62_LC_12_3_0  (
            .in0(N__50141),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__44852),
            .lcout(data_out_frame2_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i142_LC_12_3_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i142_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i142_LC_12_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i142_LC_12_3_1  (
            .in0(N__38459),
            .in1(N__32984),
            .in2(_gnd_net_),
            .in3(N__50139),
            .lcout(data_out_frame2_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i74_LC_12_3_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i74_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i74_LC_12_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i74_LC_12_3_2  (
            .in0(N__50142),
            .in1(N__39510),
            .in2(_gnd_net_),
            .in3(N__43949),
            .lcout(data_out_frame2_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i147_LC_12_3_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i147_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i147_LC_12_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i147_LC_12_3_3  (
            .in0(N__38277),
            .in1(N__43052),
            .in2(_gnd_net_),
            .in3(N__50140),
            .lcout(data_out_frame2_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i98_LC_12_3_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i98_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i98_LC_12_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i98_LC_12_3_4  (
            .in0(N__50143),
            .in1(N__38335),
            .in2(_gnd_net_),
            .in3(N__33328),
            .lcout(data_out_frame2_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_800_LC_12_3_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_800_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_800_LC_12_3_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_800_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__36306),
            .in2(_gnd_net_),
            .in3(N__40664),
            .lcout(\c0.n10829 ),
            .ltout(\c0.n10829_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_747_LC_12_3_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_747_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_747_LC_12_3_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_747_LC_12_3_6  (
            .in0(N__36255),
            .in1(N__37637),
            .in2(N__33294),
            .in3(N__46562),
            .lcout(\c0.n17755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i115_LC_12_3_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i115_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i115_LC_12_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i115_LC_12_3_7  (
            .in0(N__40899),
            .in1(N__50613),
            .in2(_gnd_net_),
            .in3(N__50138),
            .lcout(data_out_frame2_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i97_LC_12_4_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i97_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i97_LC_12_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i97_LC_12_4_0  (
            .in0(N__50123),
            .in1(N__38400),
            .in2(_gnd_net_),
            .in3(N__45766),
            .lcout(data_out_frame2_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i131_LC_12_4_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i131_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i131_LC_12_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i131_LC_12_4_1  (
            .in0(N__38275),
            .in1(N__46637),
            .in2(_gnd_net_),
            .in3(N__50120),
            .lcout(data_out_frame2_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i61_LC_12_4_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i61_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i61_LC_12_4_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i61_LC_12_4_2  (
            .in0(N__50121),
            .in1(N__50529),
            .in2(_gnd_net_),
            .in3(N__44949),
            .lcout(data_out_frame2_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_430_LC_12_4_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_430_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_430_LC_12_4_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.i3_4_lut_adj_430_LC_12_4_3  (
            .in0(N__33289),
            .in1(N__33192),
            .in2(N__33183),
            .in3(N__33090),
            .lcout(n11114),
            .ltout(n11114_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i123_LC_12_4_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i123_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i123_LC_12_4_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_out_frame2_0___i123_LC_12_4_4  (
            .in0(N__38563),
            .in1(_gnd_net_),
            .in2(N__33033),
            .in3(N__50710),
            .lcout(data_out_frame2_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i106_LC_12_4_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i106_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i106_LC_12_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i106_LC_12_4_5  (
            .in0(N__39502),
            .in1(N__41703),
            .in2(_gnd_net_),
            .in3(N__50118),
            .lcout(data_out_frame2_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i127_LC_12_4_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i127_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i127_LC_12_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i127_LC_12_4_6  (
            .in0(N__50119),
            .in1(N__39287),
            .in2(_gnd_net_),
            .in3(N__41751),
            .lcout(data_out_frame2_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i70_LC_12_4_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i70_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i70_LC_12_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i70_LC_12_4_7  (
            .in0(N__44231),
            .in1(N__36313),
            .in2(_gnd_net_),
            .in3(N__50122),
            .lcout(data_out_frame2_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i71_LC_12_5_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i71_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i71_LC_12_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i71_LC_12_5_0  (
            .in0(N__50148),
            .in1(N__41289),
            .in2(_gnd_net_),
            .in3(N__37129),
            .lcout(data_out_frame2_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i145_LC_12_5_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i145_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i145_LC_12_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i145_LC_12_5_1  (
            .in0(N__38392),
            .in1(N__33345),
            .in2(_gnd_net_),
            .in3(N__50144),
            .lcout(data_out_frame2_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i86_LC_12_5_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i86_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i86_LC_12_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i86_LC_12_5_2  (
            .in0(N__50150),
            .in1(N__38847),
            .in2(_gnd_net_),
            .in3(N__36039),
            .lcout(data_out_frame2_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i56_LC_12_5_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i56_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i56_LC_12_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i56_LC_12_5_3  (
            .in0(N__39625),
            .in1(N__33372),
            .in2(_gnd_net_),
            .in3(N__50147),
            .lcout(data_out_frame2_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i148_LC_12_5_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i148_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i148_LC_12_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i148_LC_12_5_4  (
            .in0(N__50145),
            .in1(N__38186),
            .in2(_gnd_net_),
            .in3(N__41999),
            .lcout(data_out_frame2_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i89_LC_12_5_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i89_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i89_LC_12_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i89_LC_12_5_5  (
            .in0(N__38719),
            .in1(N__46467),
            .in2(_gnd_net_),
            .in3(N__50151),
            .lcout(data_out_frame2_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i45_LC_12_5_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i45_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i45_LC_12_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i45_LC_12_5_6  (
            .in0(N__50146),
            .in1(_gnd_net_),
            .in2(N__41508),
            .in3(N__46697),
            .lcout(data_out_frame2_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i72_LC_12_5_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i72_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i72_LC_12_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i72_LC_12_5_7  (
            .in0(N__42091),
            .in1(N__41657),
            .in2(_gnd_net_),
            .in3(N__50149),
            .lcout(data_out_frame2_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49855),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_744_LC_12_6_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_744_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_744_LC_12_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_744_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__45394),
            .in2(_gnd_net_),
            .in3(N__42165),
            .lcout(\c0.n10887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i134_LC_12_6_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i134_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i134_LC_12_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i134_LC_12_6_1  (
            .in0(N__50299),
            .in1(N__44232),
            .in2(_gnd_net_),
            .in3(N__45444),
            .lcout(data_out_frame2_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i111_LC_12_6_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i111_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i111_LC_12_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i111_LC_12_6_2  (
            .in0(N__40149),
            .in1(N__42166),
            .in2(_gnd_net_),
            .in3(N__50297),
            .lcout(data_out_frame2_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i69_LC_12_6_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i69_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i69_LC_12_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i69_LC_12_6_3  (
            .in0(N__50301),
            .in1(N__38107),
            .in2(_gnd_net_),
            .in3(N__50869),
            .lcout(data_out_frame2_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i67_LC_12_6_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i67_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i67_LC_12_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i67_LC_12_6_4  (
            .in0(N__38276),
            .in1(N__43759),
            .in2(_gnd_net_),
            .in3(N__50300),
            .lcout(data_out_frame2_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i126_LC_12_6_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i126_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i126_LC_12_6_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i126_LC_12_6_5  (
            .in0(N__50298),
            .in1(_gnd_net_),
            .in2(N__45403),
            .in3(N__38450),
            .lcout(data_out_frame2_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15789_LC_12_6_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15789_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15789_LC_12_6_6 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15789_LC_12_6_6  (
            .in0(N__45650),
            .in1(N__46081),
            .in2(N__48490),
            .in3(N__36185),
            .lcout(\c0.n18645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i73_LC_12_6_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i73_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i73_LC_12_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i73_LC_12_6_7  (
            .in0(N__50302),
            .in1(N__39555),
            .in2(_gnd_net_),
            .in3(N__46382),
            .lcout(data_out_frame2_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i156_LC_12_7_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i156_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i156_LC_12_7_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i156_LC_12_7_0  (
            .in0(N__41413),
            .in1(N__33382),
            .in2(N__36264),
            .in3(N__36285),
            .lcout(\c0.data_out_frame2_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49839),
            .ce(N__50350),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_435_LC_12_7_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_435_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_435_LC_12_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_adj_435_LC_12_7_2  (
            .in0(N__33584),
            .in1(N__33569),
            .in2(N__33558),
            .in3(N__33542),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18807_bdd_4_lut_LC_12_7_4 .C_ON=1'b0;
    defparam \c0.n18807_bdd_4_lut_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18807_bdd_4_lut_LC_12_7_4 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n18807_bdd_4_lut_LC_12_7_4  (
            .in0(N__43954),
            .in1(N__33390),
            .in2(N__48689),
            .in3(N__44329),
            .lcout(\c0.n18810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15695_3_lut_LC_12_7_6 .C_ON=1'b0;
    defparam \c0.i15695_3_lut_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15695_3_lut_LC_12_7_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.i15695_3_lut_LC_12_7_6  (
            .in0(N__48635),
            .in1(N__45088),
            .in2(_gnd_net_),
            .in3(N__46089),
            .lcout(\c0.n18371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15704_3_lut_LC_12_7_7 .C_ON=1'b0;
    defparam \c0.i15704_3_lut_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15704_3_lut_LC_12_7_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \c0.i15704_3_lut_LC_12_7_7  (
            .in0(N__46088),
            .in1(N__41620),
            .in2(_gnd_net_),
            .in3(N__48636),
            .lcout(\c0.n18374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i156_2_lut_3_lut_LC_12_8_0 .C_ON=1'b0;
    defparam \c0.i156_2_lut_3_lut_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i156_2_lut_3_lut_LC_12_8_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \c0.i156_2_lut_3_lut_LC_12_8_0  (
            .in0(N__33514),
            .in1(N__33492),
            .in2(_gnd_net_),
            .in3(N__33471),
            .lcout(\c0.n155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_436_LC_12_8_1 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_436_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_436_LC_12_8_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i11_3_lut_adj_436_LC_12_8_1  (
            .in0(N__33431),
            .in1(N__33419),
            .in2(_gnd_net_),
            .in3(N__33408),
            .lcout(n25_adj_2468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i81_LC_12_8_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i81_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i81_LC_12_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i81_LC_12_8_2  (
            .in0(N__39155),
            .in1(N__46520),
            .in2(_gnd_net_),
            .in3(N__50429),
            .lcout(data_out_frame2_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15919_LC_12_8_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15919_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15919_LC_12_8_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15919_LC_12_8_3  (
            .in0(N__46117),
            .in1(N__45575),
            .in2(N__48491),
            .in3(N__40746),
            .lcout(\c0.n18807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15207_4_lut_LC_12_8_4 .C_ON=1'b0;
    defparam \c0.i15207_4_lut_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15207_4_lut_LC_12_8_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \c0.i15207_4_lut_LC_12_8_4  (
            .in0(N__33951),
            .in1(N__48389),
            .in2(N__46708),
            .in3(N__46118),
            .lcout(\c0.n18068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4698_2_lut_LC_12_8_5 .C_ON=1'b0;
    defparam \c0.i4698_2_lut_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4698_2_lut_LC_12_8_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i4698_2_lut_LC_12_8_5  (
            .in0(N__46116),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48372),
            .lcout(\c0.n7263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i101_LC_12_8_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i101_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i101_LC_12_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i101_LC_12_8_6  (
            .in0(N__38109),
            .in1(N__45185),
            .in2(_gnd_net_),
            .in3(N__50427),
            .lcout(data_out_frame2_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i65_LC_12_8_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i65_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i65_LC_12_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i65_LC_12_8_7  (
            .in0(N__50428),
            .in1(N__38399),
            .in2(_gnd_net_),
            .in3(N__46345),
            .lcout(data_out_frame2_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_12_9_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_12_9_0 .LUT_INIT=16'b1010011000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_12_9_0  (
            .in0(N__33882),
            .in1(N__33940),
            .in2(N__33753),
            .in3(N__33707),
            .lcout(r_Bit_Index_1_adj_2518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15579_3_lut_4_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \c0.i15579_3_lut_4_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15579_3_lut_4_lut_LC_12_9_1 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \c0.i15579_3_lut_4_lut_LC_12_9_1  (
            .in0(N__33857),
            .in1(N__33813),
            .in2(N__47670),
            .in3(N__33795),
            .lcout(\c0.n18259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_12_9_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_12_9_4 .LUT_INIT=16'b1001110000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_12_9_4  (
            .in0(N__33752),
            .in1(N__33667),
            .in2(N__33723),
            .in3(N__33708),
            .lcout(r_Bit_Index_2_adj_2517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_811_LC_12_9_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_811_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_811_LC_12_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_811_LC_12_9_5  (
            .in0(N__50871),
            .in1(N__41090),
            .in2(_gnd_net_),
            .in3(N__46341),
            .lcout(\c0.n17715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_LC_12_9_6 .C_ON=1'b0;
    defparam \c0.i4_2_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_LC_12_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i4_2_lut_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__33618),
            .in2(_gnd_net_),
            .in3(N__33602),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i52_LC_12_9_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i52_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i52_LC_12_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i52_LC_12_9_7  (
            .in0(N__38981),
            .in1(N__44087),
            .in2(_gnd_net_),
            .in3(N__50430),
            .lcout(data_out_frame2_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1__2276_LC_12_10_0 .C_ON=1'b0;
    defparam \c0.data_in_2__1__2276_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1__2276_LC_12_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_2__1__2276_LC_12_10_0  (
            .in0(N__34229),
            .in1(N__34273),
            .in2(_gnd_net_),
            .in3(N__34308),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3__2274_LC_12_10_1 .C_ON=1'b0;
    defparam \c0.data_in_2__3__2274_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3__2274_LC_12_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_2__3__2274_LC_12_10_1  (
            .in0(N__34257),
            .in1(N__34029),
            .in2(_gnd_net_),
            .in3(N__34230),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15693_2_lut_LC_12_10_2 .C_ON=1'b0;
    defparam \c0.i15693_2_lut_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15693_2_lut_LC_12_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15693_2_lut_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__39755),
            .in2(_gnd_net_),
            .in3(N__42797),
            .lcout(\c0.n18365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i100_LC_12_10_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i100_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i100_LC_12_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i100_LC_12_10_3  (
            .in0(N__38187),
            .in1(N__43797),
            .in2(_gnd_net_),
            .in3(N__50431),
            .lcout(data_out_frame2_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i150_LC_12_10_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i150_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i150_LC_12_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i150_LC_12_10_4  (
            .in0(N__50433),
            .in1(N__44229),
            .in2(_gnd_net_),
            .in3(N__33989),
            .lcout(data_out_frame2_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i55_LC_12_10_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i55_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i55_LC_12_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i55_LC_12_10_5  (
            .in0(N__39700),
            .in1(N__40657),
            .in2(_gnd_net_),
            .in3(N__50434),
            .lcout(data_out_frame2_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i113_LC_12_10_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i113_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i113_LC_12_10_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i113_LC_12_10_6  (
            .in0(N__50432),
            .in1(_gnd_net_),
            .in2(N__39159),
            .in3(N__46287),
            .lcout(data_out_frame2_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(_gnd_net_));
    defparam i41_4_lut_LC_12_11_0.C_ON=1'b0;
    defparam i41_4_lut_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam i41_4_lut_LC_12_11_0.LUT_INIT=16'b1111010000000100;
    LogicCell40 i41_4_lut_LC_12_11_0 (
            .in0(N__34869),
            .in1(N__33975),
            .in2(N__35248),
            .in3(N__33969),
            .lcout(n18_adj_2526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__3__2189_LC_12_11_1 .C_ON=1'b0;
    defparam \c0.data_out_8__3__2189_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__3__2189_LC_12_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_8__3__2189_LC_12_11_1  (
            .in0(N__36624),
            .in1(N__46851),
            .in2(_gnd_net_),
            .in3(N__38133),
            .lcout(data_out_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_586_LC_12_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_586_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_586_LC_12_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_586_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__36539),
            .in2(_gnd_net_),
            .in3(N__36623),
            .lcout(\c0.n17761 ),
            .ltout(\c0.n17761_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_536_LC_12_11_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_536_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_536_LC_12_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_536_LC_12_11_3  (
            .in0(N__34630),
            .in1(N__40310),
            .in2(N__34383),
            .in3(N__36802),
            .lcout(\c0.n17844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__2__2190_LC_12_11_4 .C_ON=1'b0;
    defparam \c0.data_out_8__2__2190_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__2__2190_LC_12_11_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.data_out_8__2__2190_LC_12_11_4  (
            .in0(N__34380),
            .in1(N__47313),
            .in2(N__38217),
            .in3(N__36540),
            .lcout(data_out_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_601_LC_12_11_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_601_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_601_LC_12_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_601_LC_12_11_5  (
            .in0(N__34365),
            .in1(N__34485),
            .in2(N__39993),
            .in3(N__36803),
            .lcout(\c0.n17826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i44_LC_12_11_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i44_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i44_LC_12_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i44_LC_12_11_6  (
            .in0(N__42150),
            .in1(N__43845),
            .in2(_gnd_net_),
            .in3(N__50435),
            .lcout(data_out_frame2_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49794),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15869_LC_12_11_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15869_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15869_LC_12_11_7 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15869_LC_12_11_7  (
            .in0(N__42897),
            .in1(N__35236),
            .in2(N__36444),
            .in3(N__34868),
            .lcout(\c0.n18747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_555_LC_12_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_555_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_555_LC_12_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_555_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__35857),
            .in2(_gnd_net_),
            .in3(N__37545),
            .lcout(),
            .ltout(\c0.n17807_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__2__2174_LC_12_12_1 .C_ON=1'b0;
    defparam \c0.data_out_10__2__2174_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__2__2174_LC_12_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__2__2174_LC_12_12_1  (
            .in0(N__34458),
            .in1(N__34342),
            .in2(N__34350),
            .in3(N__42942),
            .lcout(\c0.data_out_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49781),
            .ce(N__46856),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_12_12_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_12_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_715_LC_12_12_2  (
            .in0(N__34341),
            .in1(N__36937),
            .in2(_gnd_net_),
            .in3(N__37283),
            .lcout(),
            .ltout(\c0.n6_adj_2318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__6__2178_LC_12_12_3 .C_ON=1'b0;
    defparam \c0.data_out_9__6__2178_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__6__2178_LC_12_12_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__6__2178_LC_12_12_3  (
            .in0(N__35858),
            .in1(N__37017),
            .in2(N__34536),
            .in3(N__34519),
            .lcout(\c0.data_out_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49781),
            .ce(N__46856),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_615_LC_12_12_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_615_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_615_LC_12_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_615_LC_12_12_4  (
            .in0(N__39942),
            .in1(N__47733),
            .in2(N__34493),
            .in3(N__39907),
            .lcout(\c0.n6_adj_2367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__3__2181_LC_12_12_5 .C_ON=1'b0;
    defparam \c0.data_out_9__3__2181_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__3__2181_LC_12_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__3__2181_LC_12_12_5  (
            .in0(N__34452),
            .in1(N__36646),
            .in2(N__34446),
            .in3(N__37361),
            .lcout(\c0.data_out_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49781),
            .ce(N__46856),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_590_LC_12_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_590_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_590_LC_12_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_590_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__34723),
            .in2(_gnd_net_),
            .in3(N__34698),
            .lcout(\c0.n17835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_499_LC_12_13_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_499_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_499_LC_12_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_499_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__37093),
            .in2(_gnd_net_),
            .in3(N__36968),
            .lcout(),
            .ltout(\c0.data_out_9__2__N_367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_502_LC_12_13_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_502_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_502_LC_12_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_502_LC_12_13_2  (
            .in0(N__40334),
            .in1(N__34710),
            .in2(N__34425),
            .in3(N__34607),
            .lcout(),
            .ltout(\c0.n15_adj_2319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__7__2177_LC_12_13_3 .C_ON=1'b0;
    defparam \c0.data_out_9__7__2177_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__7__2177_LC_12_13_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__7__2177_LC_12_13_3  (
            .in0(N__34394),
            .in1(N__36489),
            .in2(N__34422),
            .in3(N__34419),
            .lcout(\c0.data_out_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49766),
            .ce(N__46821),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__6__2170_LC_12_13_4 .C_ON=1'b0;
    defparam \c0.data_out_10__6__2170_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__6__2170_LC_12_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__6__2170_LC_12_13_4  (
            .in0(N__34912),
            .in1(N__34410),
            .in2(N__50923),
            .in3(N__34395),
            .lcout(data_out_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49766),
            .ce(N__46821),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_610_LC_12_13_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_610_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_610_LC_12_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_610_LC_12_13_5  (
            .in0(N__34631),
            .in1(N__34911),
            .in2(N__34955),
            .in3(N__37544),
            .lcout(\c0.n17718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_564_LC_12_13_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_564_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_564_LC_12_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_564_LC_12_13_6  (
            .in0(N__50914),
            .in1(N__34724),
            .in2(N__43533),
            .in3(N__39864),
            .lcout(\c0.n17774 ),
            .ltout(\c0.n17774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__3__2173_LC_12_13_7 .C_ON=1'b0;
    defparam \c0.data_out_10__3__2173_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__3__2173_LC_12_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_10__3__2173_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__36938),
            .in2(N__34704),
            .in3(N__34569),
            .lcout(\c0.data_out_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49766),
            .ce(N__46821),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__5__2171_LC_12_14_0 .C_ON=1'b0;
    defparam \c0.data_out_10__5__2171_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__5__2171_LC_12_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__5__2171_LC_12_14_0  (
            .in0(N__36831),
            .in1(N__34591),
            .in2(N__36558),
            .in3(N__34647),
            .lcout(\c0.data_out_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49753),
            .ce(N__46843),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_490_LC_12_14_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_490_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_490_LC_12_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_490_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__34677),
            .in2(_gnd_net_),
            .in3(N__36853),
            .lcout(\c0.n6_adj_2314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_568_LC_12_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_568_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_568_LC_12_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_568_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__34913),
            .in2(_gnd_net_),
            .in3(N__37534),
            .lcout(),
            .ltout(\c0.n10801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__0__2176_LC_12_14_3 .C_ON=1'b0;
    defparam \c0.data_out_10__0__2176_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__0__2176_LC_12_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__0__2176_LC_12_14_3  (
            .in0(N__34646),
            .in1(N__36747),
            .in2(N__34635),
            .in3(N__36897),
            .lcout(\c0.data_out_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49753),
            .ce(N__46843),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_552_LC_12_14_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_552_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_552_LC_12_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_552_LC_12_14_5  (
            .in0(N__34914),
            .in1(N__34608),
            .in2(N__34956),
            .in3(N__36830),
            .lcout(),
            .ltout(\c0.n10_adj_2366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__1__2175_LC_12_14_6 .C_ON=1'b0;
    defparam \c0.data_out_10__1__2175_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__1__2175_LC_12_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__1__2175_LC_12_14_6  (
            .in0(N__35859),
            .in1(N__37535),
            .in2(N__34596),
            .in3(N__36909),
            .lcout(\c0.data_out_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49753),
            .ce(N__46843),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_577_LC_12_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_577_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_577_LC_12_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_577_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__42600),
            .in2(_gnd_net_),
            .in3(N__34564),
            .lcout(\c0.n17819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_485_LC_12_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_485_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_485_LC_12_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_485_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__39836),
            .in2(_gnd_net_),
            .in3(N__37433),
            .lcout(\c0.n6_adj_2277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_12_15_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_12_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_12_15_1  (
            .in0(N__42870),
            .in1(N__34948),
            .in2(_gnd_net_),
            .in3(N__36716),
            .lcout(),
            .ltout(\c0.n8_adj_2211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_12_15_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_12_15_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_12_15_2  (
            .in0(N__34876),
            .in1(N__40309),
            .in2(N__34932),
            .in3(N__42871),
            .lcout(n10_adj_2505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__6__2186_LC_12_15_3 .C_ON=1'b0;
    defparam \c0.data_out_8__6__2186_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__6__2186_LC_12_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_8__6__2186_LC_12_15_3  (
            .in0(N__37434),
            .in1(N__46852),
            .in2(_gnd_net_),
            .in3(N__38772),
            .lcout(data_out_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15528_2_lut_LC_12_15_4 .C_ON=1'b0;
    defparam \c0.i15528_2_lut_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15528_2_lut_LC_12_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15528_2_lut_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__39835),
            .in2(_gnd_net_),
            .in3(N__42868),
            .lcout(),
            .ltout(\c0.n18222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15864_LC_12_15_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15864_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15864_LC_12_15_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15864_LC_12_15_5  (
            .in0(N__34884),
            .in1(N__35249),
            .in2(N__34929),
            .in3(N__34877),
            .lcout(),
            .ltout(\c0.n18693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18693_bdd_4_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \c0.n18693_bdd_4_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18693_bdd_4_lut_LC_12_15_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18693_bdd_4_lut_LC_12_15_6  (
            .in0(N__35250),
            .in1(N__35802),
            .in2(N__34926),
            .in3(N__34983),
            .lcout(n18696),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_12_15_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_12_15_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_12_15_7  (
            .in0(N__42869),
            .in1(N__37071),
            .in2(_gnd_net_),
            .in3(N__34910),
            .lcout(\c0.n5_adj_2347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15968_LC_12_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15968_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15968_LC_12_16_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15968_LC_12_16_0  (
            .in0(N__35231),
            .in1(N__34974),
            .in2(N__35013),
            .in3(N__34872),
            .lcout(),
            .ltout(\c0.n18867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18867_bdd_4_lut_LC_12_16_1 .C_ON=1'b0;
    defparam \c0.n18867_bdd_4_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18867_bdd_4_lut_LC_12_16_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18867_bdd_4_lut_LC_12_16_1  (
            .in0(N__35262),
            .in1(N__34989),
            .in2(N__35253),
            .in3(N__35232),
            .lcout(),
            .ltout(n18870_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_821_LC_12_16_2.C_ON=1'b0;
    defparam i24_4_lut_adj_821_LC_12_16_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_821_LC_12_16_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 i24_4_lut_adj_821_LC_12_16_2 (
            .in0(N__35233),
            .in1(N__35106),
            .in2(N__35097),
            .in3(N__35094),
            .lcout(n10_adj_2530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__7__2193_LC_12_16_3 .C_ON=1'b0;
    defparam \c0.data_out_7__7__2193_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7__2193_LC_12_16_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_7__7__2193_LC_12_16_3  (
            .in0(N__39183),
            .in1(N__47871),
            .in2(N__47810),
            .in3(N__39900),
            .lcout(\c0.data_out_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_16_4  (
            .in0(N__35853),
            .in1(N__36807),
            .in2(_gnd_net_),
            .in3(N__42872),
            .lcout(\c0.n5_adj_2214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15601_2_lut_LC_12_16_6 .C_ON=1'b0;
    defparam \c0.i15601_2_lut_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15601_2_lut_LC_12_16_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i15601_2_lut_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__35004),
            .in2(_gnd_net_),
            .in3(N__42873),
            .lcout(\c0.n18190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__2__2246_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.data_out_1__2__2246_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2__2246_LC_12_17_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_1__2__2246_LC_12_17_0  (
            .in0(N__47142),
            .in1(N__43264),
            .in2(N__35814),
            .in3(N__47690),
            .lcout(\c0.data_out_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15721_2_lut_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.i15721_2_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15721_2_lut_LC_12_17_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.i15721_2_lut_LC_12_17_1  (
            .in0(N__47127),
            .in1(N__43259),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n11277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_17_3  (
            .in0(N__42866),
            .in1(N__35822),
            .in2(_gnd_net_),
            .in3(N__35793),
            .lcout(\c0.n2_adj_2348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15666_2_lut_LC_12_17_4 .C_ON=1'b0;
    defparam \c0.i15666_2_lut_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15666_2_lut_LC_12_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15666_2_lut_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__37249),
            .in2(_gnd_net_),
            .in3(N__42865),
            .lcout(\c0.n18334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4__2196_LC_12_17_5 .C_ON=1'b0;
    defparam \c0.data_out_7__4__2196_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4__2196_LC_12_17_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_7__4__2196_LC_12_17_5  (
            .in0(N__38487),
            .in1(N__47883),
            .in2(N__47814),
            .in3(N__35852),
            .lcout(\c0.data_out_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__2__2230_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.data_out_3__2__2230_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2__2230_LC_12_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_3__2__2230_LC_12_17_6  (
            .in0(N__35823),
            .in1(N__40270),
            .in2(_gnd_net_),
            .in3(N__43265),
            .lcout(data_out_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15665_2_lut_LC_12_17_7 .C_ON=1'b0;
    defparam \c0.i15665_2_lut_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15665_2_lut_LC_12_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15665_2_lut_LC_12_17_7  (
            .in0(N__42867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35810),
            .lcout(\c0.n18223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__2__2238_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.data_out_2__2__2238_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__2__2238_LC_12_19_1 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \c0.data_out_2__2__2238_LC_12_19_1  (
            .in0(N__43347),
            .in1(N__35792),
            .in2(_gnd_net_),
            .in3(N__47123),
            .lcout(data_out_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49741),
            .ce(),
            .sr(_gnd_net_));
    defparam \control.PHASES_i4_LC_12_27_2 .C_ON=1'b0;
    defparam \control.PHASES_i4_LC_12_27_2 .SEQ_MODE=4'b1000;
    defparam \control.PHASES_i4_LC_12_27_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \control.PHASES_i4_LC_12_27_2  (
            .in0(N__35689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35576),
            .lcout(PIN_24_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49838),
            .ce(N__35760),
            .sr(N__35748));
    defparam \control.PHASES_i5_LC_12_28_6 .C_ON=1'b0;
    defparam \control.PHASES_i5_LC_12_28_6 .SEQ_MODE=4'b1000;
    defparam \control.PHASES_i5_LC_12_28_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \control.PHASES_i5_LC_12_28_6  (
            .in0(_gnd_net_),
            .in1(N__35470),
            .in2(_gnd_net_),
            .in3(N__35545),
            .lcout(PIN_23_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49847),
            .ce(N__35727),
            .sr(N__35700));
    defparam \control.i1_4_lut_LC_12_29_5 .C_ON=1'b0;
    defparam \control.i1_4_lut_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \control.i1_4_lut_LC_12_29_5 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \control.i1_4_lut_LC_12_29_5  (
            .in0(N__35691),
            .in1(N__35577),
            .in2(N__35472),
            .in3(N__35325),
            .lcout(\control.PHASES_5_N_2130_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_786_LC_13_1_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_786_LC_13_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_786_LC_13_1_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_786_LC_13_1_0  (
            .in0(N__44437),
            .in1(N__50823),
            .in2(N__35277),
            .in3(N__41324),
            .lcout(\c0.n15_adj_2445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_802_LC_13_1_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_802_LC_13_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_802_LC_13_1_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_802_LC_13_1_1  (
            .in0(_gnd_net_),
            .in1(N__35899),
            .in2(_gnd_net_),
            .in3(N__35984),
            .lcout(\c0.n10890 ),
            .ltout(\c0.n10890_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_805_LC_13_1_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_805_LC_13_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_805_LC_13_1_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_805_LC_13_1_2  (
            .in0(N__50620),
            .in1(N__35961),
            .in2(N__35949),
            .in3(N__40560),
            .lcout(),
            .ltout(\c0.n16_adj_2448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i155_LC_13_1_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i155_LC_13_1_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i155_LC_13_1_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i155_LC_13_1_3  (
            .in0(N__35931),
            .in1(N__35946),
            .in2(N__35934),
            .in3(N__41897),
            .lcout(\c0.data_out_frame2_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__50419),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_784_LC_13_1_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_784_LC_13_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_784_LC_13_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_784_LC_13_1_4  (
            .in0(N__35930),
            .in1(N__40535),
            .in2(_gnd_net_),
            .in3(N__36243),
            .lcout(),
            .ltout(\c0.n14_adj_2444_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i157_LC_13_1_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i157_LC_13_1_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i157_LC_13_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i157_LC_13_1_5  (
            .in0(N__36138),
            .in1(N__35913),
            .in2(N__35907),
            .in3(N__40703),
            .lcout(\c0.data_out_frame2_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__50419),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_693_LC_13_1_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_693_LC_13_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_693_LC_13_1_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_693_LC_13_1_6  (
            .in0(N__35900),
            .in1(_gnd_net_),
            .in2(N__43958),
            .in3(_gnd_net_),
            .lcout(\c0.n10825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i166_LC_13_2_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i166_LC_13_2_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i166_LC_13_2_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i166_LC_13_2_0  (
            .in0(N__36072),
            .in1(N__44913),
            .in2(N__35868),
            .in3(N__37743),
            .lcout(\c0.data_out_frame2_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49879),
            .ce(N__50467),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_adj_532_LC_13_2_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_adj_532_LC_13_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_adj_532_LC_13_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_2_lut_3_lut_adj_532_LC_13_2_1  (
            .in0(N__37802),
            .in1(N__44160),
            .in2(_gnd_net_),
            .in3(N__46475),
            .lcout(\c0.n16_adj_2358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_428_LC_13_2_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_428_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_428_LC_13_2_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_428_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(N__36228),
            .in2(_gnd_net_),
            .in3(N__40777),
            .lcout(),
            .ltout(\c0.n10720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_783_LC_13_2_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_783_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_783_LC_13_2_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_783_LC_13_2_3  (
            .in0(N__36149),
            .in1(N__36070),
            .in2(N__36192),
            .in3(N__42978),
            .lcout(\c0.n17838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_797_LC_13_2_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_797_LC_13_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_797_LC_13_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_797_LC_13_2_4  (
            .in0(_gnd_net_),
            .in1(N__46535),
            .in2(_gnd_net_),
            .in3(N__36189),
            .lcout(\c0.n10819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_LC_13_2_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_LC_13_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_LC_13_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_2_lut_3_lut_LC_13_2_5  (
            .in0(N__36134),
            .in1(N__41564),
            .in2(_gnd_net_),
            .in3(N__50885),
            .lcout(),
            .ltout(\c0.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i158_LC_13_2_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i158_LC_13_2_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i158_LC_13_2_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i158_LC_13_2_6  (
            .in0(N__36071),
            .in1(N__36117),
            .in2(N__36108),
            .in3(N__36105),
            .lcout(\c0.data_out_frame2_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49879),
            .ce(N__50467),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_778_LC_13_2_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_778_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_778_LC_13_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_778_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(N__41950),
            .in2(_gnd_net_),
            .in3(N__36429),
            .lcout(\c0.n10839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i68_LC_13_3_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i68_LC_13_3_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i68_LC_13_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i68_LC_13_3_0  (
            .in0(N__38182),
            .in1(N__40776),
            .in2(_gnd_net_),
            .in3(N__50244),
            .lcout(data_out_frame2_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i120_LC_13_3_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i120_LC_13_3_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i120_LC_13_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i120_LC_13_3_1  (
            .in0(N__50241),
            .in1(N__39632),
            .in2(_gnd_net_),
            .in3(N__40197),
            .lcout(data_out_frame2_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_792_LC_13_3_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_792_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_792_LC_13_3_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_792_LC_13_3_2  (
            .in0(N__36060),
            .in1(N__36050),
            .in2(N__37583),
            .in3(N__36239),
            .lcout(),
            .ltout(\c0.n12_adj_2446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_793_LC_13_3_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_793_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_793_LC_13_3_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_793_LC_13_3_3  (
            .in0(N__36011),
            .in1(N__45506),
            .in2(N__35988),
            .in3(N__42052),
            .lcout(\c0.n17792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i112_LC_13_3_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i112_LC_13_3_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i112_LC_13_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i112_LC_13_3_4  (
            .in0(N__40096),
            .in1(N__42223),
            .in2(_gnd_net_),
            .in3(N__50240),
            .lcout(data_out_frame2_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i139_LC_13_3_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i139_LC_13_3_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i139_LC_13_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i139_LC_13_3_5  (
            .in0(N__50243),
            .in1(N__38564),
            .in2(_gnd_net_),
            .in3(N__43019),
            .lcout(data_out_frame2_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_803_LC_13_3_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_803_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_803_LC_13_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_803_LC_13_3_6  (
            .in0(N__36227),
            .in1(N__40775),
            .in2(_gnd_net_),
            .in3(N__46534),
            .lcout(\c0.n17859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i135_LC_13_3_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i135_LC_13_3_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i135_LC_13_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i135_LC_13_3_7  (
            .in0(N__50242),
            .in1(N__41288),
            .in2(_gnd_net_),
            .in3(N__42261),
            .lcout(data_out_frame2_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i48_LC_13_4_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i48_LC_13_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i48_LC_13_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i48_LC_13_4_0  (
            .in0(N__50128),
            .in1(N__40098),
            .in2(_gnd_net_),
            .in3(N__44649),
            .lcout(data_out_frame2_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i107_LC_13_4_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i107_LC_13_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i107_LC_13_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i107_LC_13_4_1  (
            .in0(N__39425),
            .in1(N__37212),
            .in2(_gnd_net_),
            .in3(N__50124),
            .lcout(data_out_frame2_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i43_LC_13_4_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i43_LC_13_4_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i43_LC_13_4_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i43_LC_13_4_2  (
            .in0(N__50127),
            .in1(N__39426),
            .in2(_gnd_net_),
            .in3(N__41555),
            .lcout(data_out_frame2_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i78_LC_13_4_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i78_LC_13_4_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i78_LC_13_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i78_LC_13_4_3  (
            .in0(N__39350),
            .in1(N__44613),
            .in2(_gnd_net_),
            .in3(N__50130),
            .lcout(data_out_frame2_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i132_LC_13_4_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i132_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i132_LC_13_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i132_LC_13_4_4  (
            .in0(N__50126),
            .in1(N__38174),
            .in2(_gnd_net_),
            .in3(N__41946),
            .lcout(data_out_frame2_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i64_LC_13_4_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i64_LC_13_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i64_LC_13_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i64_LC_13_4_5  (
            .in0(N__39231),
            .in1(N__41184),
            .in2(_gnd_net_),
            .in3(N__50129),
            .lcout(data_out_frame2_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i129_LC_13_4_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i129_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i129_LC_13_4_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i129_LC_13_4_6  (
            .in0(N__50125),
            .in1(_gnd_net_),
            .in2(N__38388),
            .in3(N__37178),
            .lcout(data_out_frame2_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_506_LC_13_4_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_506_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_506_LC_13_4_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_506_LC_13_4_7  (
            .in0(N__43752),
            .in1(N__50702),
            .in2(N__46645),
            .in3(N__41366),
            .lcout(\c0.n10864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i124_LC_13_5_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i124_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i124_LC_13_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i124_LC_13_5_0  (
            .in0(N__41451),
            .in1(N__36426),
            .in2(_gnd_net_),
            .in3(N__50246),
            .lcout(data_out_frame2_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i66_LC_13_5_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i66_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i66_LC_13_5_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i66_LC_13_5_1  (
            .in0(N__50249),
            .in1(_gnd_net_),
            .in2(N__38320),
            .in3(N__44309),
            .lcout(data_out_frame2_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i116_LC_13_5_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i116_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i116_LC_13_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i116_LC_13_5_2  (
            .in0(N__38980),
            .in1(N__45040),
            .in2(_gnd_net_),
            .in3(N__50245),
            .lcout(data_out_frame2_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i92_LC_13_5_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i92_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i92_LC_13_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i92_LC_13_5_3  (
            .in0(N__50251),
            .in1(N__41452),
            .in2(_gnd_net_),
            .in3(N__45614),
            .lcout(data_out_frame2_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i47_LC_13_5_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i47_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i47_LC_13_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i47_LC_13_5_4  (
            .in0(N__40148),
            .in1(N__41853),
            .in2(_gnd_net_),
            .in3(N__50248),
            .lcout(data_out_frame2_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i90_LC_13_5_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i90_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i90_LC_13_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i90_LC_13_5_5  (
            .in0(N__50250),
            .in1(N__38639),
            .in2(_gnd_net_),
            .in3(N__45574),
            .lcout(data_out_frame2_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i94_LC_13_5_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i94_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i94_LC_13_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i94_LC_13_5_6  (
            .in0(N__38445),
            .in1(N__45234),
            .in2(_gnd_net_),
            .in3(N__50252),
            .lcout(data_out_frame2_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i133_LC_13_5_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i133_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i133_LC_13_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i133_LC_13_5_7  (
            .in0(N__50247),
            .in1(N__38083),
            .in2(_gnd_net_),
            .in3(N__48219),
            .lcout(data_out_frame2_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i85_LC_13_6_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i85_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i85_LC_13_6_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i85_LC_13_6_0  (
            .in0(N__50402),
            .in1(_gnd_net_),
            .in2(N__38905),
            .in3(N__41025),
            .lcout(data_out_frame2_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i143_LC_13_6_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i143_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i143_LC_13_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i143_LC_13_6_1  (
            .in0(N__39282),
            .in1(N__42290),
            .in2(_gnd_net_),
            .in3(N__50401),
            .lcout(data_out_frame2_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_678_LC_13_6_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_678_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_678_LC_13_6_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_678_LC_13_6_2  (
            .in0(N__45613),
            .in1(N__45654),
            .in2(N__46474),
            .in3(N__45570),
            .lcout(\c0.n10_adj_2411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i105_LC_13_6_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i105_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i105_LC_13_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i105_LC_13_6_3  (
            .in0(N__39554),
            .in1(N__45849),
            .in2(_gnd_net_),
            .in3(N__50398),
            .lcout(data_out_frame2_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i117_LC_13_6_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i117_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i117_LC_13_6_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i117_LC_13_6_4  (
            .in0(N__50399),
            .in1(_gnd_net_),
            .in2(N__38904),
            .in3(N__44418),
            .lcout(data_out_frame2_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i91_LC_13_6_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i91_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i91_LC_13_6_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i91_LC_13_6_5  (
            .in0(N__45655),
            .in1(_gnd_net_),
            .in2(N__38556),
            .in3(N__50403),
            .lcout(data_out_frame2_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i125_LC_13_6_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i125_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i125_LC_13_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i125_LC_13_6_6  (
            .in0(N__50400),
            .in1(N__50505),
            .in2(_gnd_net_),
            .in3(N__45003),
            .lcout(data_out_frame2_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_762_LC_13_6_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_762_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_762_LC_13_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_762_LC_13_6_7  (
            .in0(N__45039),
            .in1(N__45233),
            .in2(_gnd_net_),
            .in3(N__41325),
            .lcout(\c0.n10_adj_2440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_530_LC_13_7_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_530_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_530_LC_13_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_530_LC_13_7_0  (
            .in0(N__44994),
            .in1(N__41357),
            .in2(_gnd_net_),
            .in3(N__45435),
            .lcout(\c0.n6_adj_2357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15983_LC_13_7_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15983_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15983_LC_13_7_1 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15983_LC_13_7_1  (
            .in0(N__41015),
            .in1(N__46120),
            .in2(N__48688),
            .in3(N__50586),
            .lcout(),
            .ltout(\c0.n18879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18879_bdd_4_lut_LC_13_7_2 .C_ON=1'b0;
    defparam \c0.n18879_bdd_4_lut_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18879_bdd_4_lut_LC_13_7_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n18879_bdd_4_lut_LC_13_7_2  (
            .in0(N__41227),
            .in1(N__48631),
            .in2(N__36366),
            .in3(N__50868),
            .lcout(\c0.n18160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15799_LC_13_7_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15799_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15799_LC_13_7_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15799_LC_13_7_3  (
            .in0(N__36428),
            .in1(N__45041),
            .in2(N__48687),
            .in3(N__46119),
            .lcout(\c0.n18657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_694_LC_13_7_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_694_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_694_LC_13_7_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_694_LC_13_7_4  (
            .in0(N__41228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41865),
            .lcout(\c0.n10852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_794_LC_13_7_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_794_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_794_LC_13_7_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_794_LC_13_7_5  (
            .in0(N__40689),
            .in1(N__44330),
            .in2(N__36348),
            .in3(N__36315),
            .lcout(\c0.n14_adj_2447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i108_LC_13_7_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i108_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i108_LC_13_7_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i108_LC_13_7_6  (
            .in0(N__42039),
            .in1(_gnd_net_),
            .in2(N__42148),
            .in3(N__50404),
            .lcout(data_out_frame2_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i63_LC_13_7_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i63_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i63_LC_13_7_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i63_LC_13_7_7  (
            .in0(N__50405),
            .in1(_gnd_net_),
            .in2(N__39288),
            .in3(N__44683),
            .lcout(data_out_frame2_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15809_LC_13_8_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15809_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15809_LC_13_8_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15809_LC_13_8_0  (
            .in0(N__36398),
            .in1(N__48637),
            .in2(N__36279),
            .in3(N__46122),
            .lcout(\c0.n18669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_13_8_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_13_8_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_13_8_1  (
            .in0(N__46121),
            .in1(_gnd_net_),
            .in2(N__37679),
            .in3(N__40551),
            .lcout(\c0.n5_adj_2274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15690_3_lut_LC_13_8_2 .C_ON=1'b0;
    defparam \c0.i15690_3_lut_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15690_3_lut_LC_13_8_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15690_3_lut_LC_13_8_2  (
            .in0(N__41815),
            .in1(N__48638),
            .in2(_gnd_net_),
            .in3(N__46123),
            .lcout(\c0.n18308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_702_LC_13_8_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_702_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_702_LC_13_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_702_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__37179),
            .in2(_gnd_net_),
            .in3(N__44677),
            .lcout(),
            .ltout(\c0.n6_adj_2422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_704_LC_13_8_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_704_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_704_LC_13_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_704_LC_13_8_4  (
            .in0(N__46397),
            .in1(N__36427),
            .in2(N__36402),
            .in3(N__42977),
            .lcout(\c0.n17780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i149_LC_13_8_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i149_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i149_LC_13_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i149_LC_13_8_5  (
            .in0(N__38108),
            .in1(N__36399),
            .in2(_gnd_net_),
            .in3(N__50463),
            .lcout(data_out_frame2_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i41_LC_13_8_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i41_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i41_LC_13_8_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i41_LC_13_8_6  (
            .in0(N__50464),
            .in1(_gnd_net_),
            .in2(N__39552),
            .in3(N__41365),
            .lcout(data_out_frame2_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i49_LC_13_8_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i49_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i49_LC_13_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i49_LC_13_8_7  (
            .in0(N__37675),
            .in1(N__39136),
            .in2(_gnd_net_),
            .in3(N__50465),
            .lcout(data_out_frame2_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_808_LC_13_9_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_808_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_808_LC_13_9_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_808_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__46331),
            .in2(_gnd_net_),
            .in3(N__50870),
            .lcout(),
            .ltout(\c0.n10870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_713_LC_13_9_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_713_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_713_LC_13_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_713_LC_13_9_2  (
            .in0(N__37671),
            .in1(N__37213),
            .in2(N__36390),
            .in3(N__44086),
            .lcout(\c0.n27_adj_2428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_741_LC_13_9_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_741_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_741_LC_13_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_741_LC_13_9_4  (
            .in0(N__45856),
            .in1(N__44810),
            .in2(N__46719),
            .in3(N__40656),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_9_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_9_6 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_9_6  (
            .in0(N__48690),
            .in1(N__46064),
            .in2(N__36375),
            .in3(N__41364),
            .lcout(\c0.n6_adj_2275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_594_LC_13_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_594_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_594_LC_13_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_594_LC_13_9_7  (
            .in0(N__39986),
            .in1(N__36553),
            .in2(_gnd_net_),
            .in3(N__36630),
            .lcout(\c0.n10542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15726_2_lut_3_lut_LC_13_10_2 .C_ON=1'b0;
    defparam \c0.i15726_2_lut_3_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15726_2_lut_3_lut_LC_13_10_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i15726_2_lut_3_lut_LC_13_10_2  (
            .in0(N__47686),
            .in1(N__47354),
            .in2(_gnd_net_),
            .in3(N__47137),
            .lcout(\c0.n11056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15522_2_lut_LC_13_10_4 .C_ON=1'b0;
    defparam \c0.i15522_2_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15522_2_lut_LC_13_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15522_2_lut_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__38507),
            .in2(_gnd_net_),
            .in3(N__47353),
            .lcout(),
            .ltout(\c0.n18199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2__2198_LC_13_10_5 .C_ON=1'b0;
    defparam \c0.data_out_7__2__2198_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2__2198_LC_13_10_5 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.data_out_7__2__2198_LC_13_10_5  (
            .in0(N__47138),
            .in1(N__47687),
            .in2(N__36492),
            .in3(N__42941),
            .lcout(\c0.data_out_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49818),
            .ce(N__47898),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_498_LC_13_10_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_498_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_498_LC_13_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_498_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__40311),
            .in2(_gnd_net_),
            .in3(N__37066),
            .lcout(\c0.n17832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7__2201_LC_13_11_0 .C_ON=1'b0;
    defparam \c0.data_out_6__7__2201_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7__2201_LC_13_11_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.data_out_6__7__2201_LC_13_11_0  (
            .in0(N__47065),
            .in1(N__47358),
            .in2(N__39576),
            .in3(N__36435),
            .lcout(\c0.data_out_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49807),
            .ce(N__43424),
            .sr(_gnd_net_));
    defparam \c0.i15536_3_lut_LC_13_11_1 .C_ON=1'b0;
    defparam \c0.i15536_3_lut_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15536_3_lut_LC_13_11_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15536_3_lut_LC_13_11_1  (
            .in0(N__37483),
            .in1(N__47603),
            .in2(_gnd_net_),
            .in3(N__37278),
            .lcout(),
            .ltout(\c0.n18242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6__2202_LC_13_11_2 .C_ON=1'b0;
    defparam \c0.data_out_6__6__2202_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6__2202_LC_13_11_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_6__6__2202_LC_13_11_2  (
            .in0(N__47064),
            .in1(N__39654),
            .in2(N__36465),
            .in3(N__47357),
            .lcout(\c0.data_out_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49807),
            .ce(N__43424),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_13_11_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_13_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_13_11_3  (
            .in0(N__47734),
            .in1(N__36458),
            .in2(_gnd_net_),
            .in3(N__42857),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15570_3_lut_LC_13_11_4 .C_ON=1'b0;
    defparam \c0.i15570_3_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15570_3_lut_LC_13_11_4 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \c0.i15570_3_lut_LC_13_11_4  (
            .in0(N__47602),
            .in1(N__36890),
            .in2(_gnd_net_),
            .in3(N__43529),
            .lcout(\c0.n18247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15535_3_lut_LC_13_11_5 .C_ON=1'b0;
    defparam \c0.i15535_3_lut_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15535_3_lut_LC_13_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15535_3_lut_LC_13_11_5  (
            .in0(N__47610),
            .in1(N__39756),
            .in2(_gnd_net_),
            .in3(N__37277),
            .lcout(),
            .ltout(\c0.n18238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5__2203_LC_13_11_6 .C_ON=1'b0;
    defparam \c0.data_out_6__5__2203_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5__2203_LC_13_11_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_6__5__2203_LC_13_11_6  (
            .in0(N__47063),
            .in1(N__38789),
            .in2(N__36810),
            .in3(N__47356),
            .lcout(\c0.data_out_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49807),
            .ce(N__43424),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4__2204_LC_13_11_7 .C_ON=1'b0;
    defparam \c0.data_out_6__4__2204_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4__2204_LC_13_11_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__4__2204_LC_13_11_7  (
            .in0(N__47355),
            .in1(N__38864),
            .in2(N__40023),
            .in3(N__47066),
            .lcout(\c0.data_out_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49807),
            .ce(N__43424),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__1__2183_LC_13_12_0 .C_ON=1'b0;
    defparam \c0.data_out_9__1__2183_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__1__2183_LC_13_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__1__2183_LC_13_12_0  (
            .in0(N__36626),
            .in1(N__36786),
            .in2(N__36684),
            .in3(N__36769),
            .lcout(\c0.data_out_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49795),
            .ce(N__46844),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_592_LC_13_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_592_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_592_LC_13_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_592_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__36735),
            .in2(_gnd_net_),
            .in3(N__36717),
            .lcout(\c0.n17745 ),
            .ltout(\c0.n17745_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__7__2169_LC_13_12_2 .C_ON=1'b0;
    defparam \c0.data_out_10__7__2169_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__7__2169_LC_13_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__7__2169_LC_13_12_2  (
            .in0(N__36675),
            .in1(N__37005),
            .in2(N__36666),
            .in3(N__42605),
            .lcout(\c0.data_out_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49795),
            .ce(N__46844),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_13_12_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_13_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_13_12_3  (
            .in0(N__36933),
            .in1(N__36625),
            .in2(_gnd_net_),
            .in3(N__42858),
            .lcout(\c0.n8_adj_2219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15544_2_lut_LC_13_12_4 .C_ON=1'b0;
    defparam \c0.i15544_2_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15544_2_lut_LC_13_12_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i15544_2_lut_LC_13_12_4  (
            .in0(N__42859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36591),
            .lcout(\c0.n18376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__5__2211_LC_13_13_4 .C_ON=1'b0;
    defparam \c0.data_out_5__5__2211_LC_13_13_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__5__2211_LC_13_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__5__2211_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__39305),
            .in2(_gnd_net_),
            .in3(N__47380),
            .lcout(\c0.data_out_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(N__43413),
            .sr(N__43478));
    defparam \c0.i3_4_lut_adj_539_LC_13_13_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_539_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_539_LC_13_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_539_LC_13_13_5  (
            .in0(N__37092),
            .in1(N__37070),
            .in2(N__37036),
            .in3(N__37469),
            .lcout(\c0.n17730 ),
            .ltout(\c0.n17730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_544_LC_13_13_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_544_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_544_LC_13_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_544_LC_13_13_6  (
            .in0(N__37004),
            .in1(N__36989),
            .in2(N__36972),
            .in3(N__36969),
            .lcout(),
            .ltout(\c0.n14_adj_2363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_546_LC_13_13_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_546_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_546_LC_13_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_3_lut_adj_546_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__42536),
            .in2(N__36954),
            .in3(N__36951),
            .lcout(\c0.n17877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_443_LC_13_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_443_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_443_LC_13_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_443_LC_13_14_2  (
            .in0(N__39741),
            .in1(N__43528),
            .in2(_gnd_net_),
            .in3(N__37275),
            .lcout(\c0.n17816 ),
            .ltout(\c0.n17816_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_13_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_13_14_3  (
            .in0(N__36942),
            .in1(N__40322),
            .in2(N__36912),
            .in3(N__36908),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_13_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_13_14_5  (
            .in0(N__37276),
            .in1(N__39742),
            .in2(N__37503),
            .in3(N__42929),
            .lcout(\c0.n17786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__1__2199_LC_13_14_7 .C_ON=1'b0;
    defparam \c0.data_out_7__1__2199_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1__2199_LC_13_14_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_7__1__2199_LC_13_14_7  (
            .in0(N__47365),
            .in1(N__47140),
            .in2(N__38595),
            .in3(N__36870),
            .lcout(\c0.data_out_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49767),
            .ce(N__47885),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_572_LC_13_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_572_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_572_LC_13_15_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_572_LC_13_15_0  (
            .in0(N__47736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36829),
            .lcout(\c0.n17829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0__2208_LC_13_15_1 .C_ON=1'b0;
    defparam \c0.data_out_6__0__2208_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0__2208_LC_13_15_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_6__0__2208_LC_13_15_1  (
            .in0(N__39111),
            .in1(N__43382),
            .in2(N__47809),
            .in3(N__37536),
            .lcout(data_out_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49754),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_13_15_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_13_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_13_15_3  (
            .in0(N__39821),
            .in1(N__37313),
            .in2(_gnd_net_),
            .in3(N__42489),
            .lcout(\c0.n10680 ),
            .ltout(\c0.n10680_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15682_4_lut_LC_13_15_4 .C_ON=1'b0;
    defparam \c0.i15682_4_lut_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15682_4_lut_LC_13_15_4 .LUT_INIT=16'b0100100010000100;
    LogicCell40 \c0.i15682_4_lut_LC_13_15_4  (
            .in0(N__37494),
            .in1(N__47660),
            .in2(N__37488),
            .in3(N__37482),
            .lcout(\c0.n18250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_513_LC_13_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_513_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_513_LC_13_15_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_513_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__37441),
            .in2(_gnd_net_),
            .in3(N__37403),
            .lcout(\c0.n17771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1__2215_LC_13_16_0 .C_ON=1'b0;
    defparam \c0.data_out_5__1__2215_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1__2215_LC_13_16_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.data_out_5__1__2215_LC_13_16_0  (
            .in0(N__47139),
            .in1(N__47688),
            .in2(N__39453),
            .in3(N__47402),
            .lcout(data_out_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49742),
            .ce(N__43396),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__4__2212_LC_13_17_3 .C_ON=1'b0;
    defparam \c0.data_out_5__4__2212_LC_13_17_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__4__2212_LC_13_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__4__2212_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__39381),
            .in2(_gnd_net_),
            .in3(N__47398),
            .lcout(\c0.data_out_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49728),
            .ce(N__43383),
            .sr(N__43462));
    defparam \c0.i1_3_lut_4_lut_adj_505_LC_14_1_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_505_LC_14_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_505_LC_14_1_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_505_LC_14_1_0  (
            .in0(N__37220),
            .in1(N__46233),
            .in2(N__42275),
            .in3(N__37187),
            .lcout(\c0.n17880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15894_LC_14_1_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15894_LC_14_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15894_LC_14_1_2 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15894_LC_14_1_2  (
            .in0(N__50819),
            .in1(N__46165),
            .in2(N__48703),
            .in3(N__41323),
            .lcout(),
            .ltout(\c0.n18759_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18759_bdd_4_lut_LC_14_1_3 .C_ON=1'b0;
    defparam \c0.n18759_bdd_4_lut_LC_14_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18759_bdd_4_lut_LC_14_1_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n18759_bdd_4_lut_LC_14_1_3  (
            .in0(N__37140),
            .in1(N__40589),
            .in2(N__37692),
            .in3(N__48678),
            .lcout(\c0.n18762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_14_1_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_14_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_14_1_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_14_1_4  (
            .in0(N__40590),
            .in1(N__41229),
            .in2(N__37689),
            .in3(N__41189),
            .lcout(\c0.n10778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i121_LC_14_1_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i121_LC_14_1_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i121_LC_14_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i121_LC_14_1_5  (
            .in0(N__46234),
            .in1(N__38715),
            .in2(_gnd_net_),
            .in3(N__50473),
            .lcout(data_out_frame2_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49887),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15938_LC_14_1_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15938_LC_14_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15938_LC_14_1_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15938_LC_14_1_6  (
            .in0(N__40941),
            .in1(N__40198),
            .in2(N__48704),
            .in3(N__46166),
            .lcout(\c0.n18813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_429_LC_14_1_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_429_LC_14_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_429_LC_14_1_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_429_LC_14_1_7  (
            .in0(N__40199),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40942),
            .lcout(\c0.n10920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_431_LC_14_2_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_431_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_431_LC_14_2_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_431_LC_14_2_0  (
            .in0(N__46303),
            .in1(N__42265),
            .in2(N__45861),
            .in3(N__41766),
            .lcout(\c0.n17783 ),
            .ltout(\c0.n17783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_14_2_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_14_2_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_14_2_1  (
            .in0(N__37821),
            .in1(N__43675),
            .in2(N__37644),
            .in3(N__37641),
            .lcout(),
            .ltout(\c0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i153_LC_14_2_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i153_LC_14_2_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i153_LC_14_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i153_LC_14_2_2  (
            .in0(N__37626),
            .in1(N__44709),
            .in2(N__37605),
            .in3(N__40173),
            .lcout(\c0.data_out_frame2_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__50474),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_751_LC_14_2_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_751_LC_14_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_751_LC_14_2_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_751_LC_14_2_3  (
            .in0(N__41565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41035),
            .lcout(),
            .ltout(\c0.n10813_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_687_LC_14_2_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_687_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_687_LC_14_2_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_687_LC_14_2_4  (
            .in0(N__37587),
            .in1(N__46487),
            .in2(N__37563),
            .in3(N__37560),
            .lcout(),
            .ltout(\c0.n15_adj_2414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i162_LC_14_2_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i162_LC_14_2_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i162_LC_14_2_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i162_LC_14_2_5  (
            .in0(N__37908),
            .in1(N__41109),
            .in2(N__37902),
            .in3(N__40550),
            .lcout(\c0.data_out_frame2_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__50474),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_739_LC_14_3_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_739_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_739_LC_14_3_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_739_LC_14_3_0  (
            .in0(N__45540),
            .in1(N__41882),
            .in2(N__40629),
            .in3(N__37754),
            .lcout(),
            .ltout(\c0.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i160_LC_14_3_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i160_LC_14_3_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i160_LC_14_3_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i160_LC_14_3_1  (
            .in0(N__40164),
            .in1(N__37887),
            .in2(N__37875),
            .in3(N__40671),
            .lcout(\c0.data_out_frame2_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49880),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_725_LC_14_3_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_725_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_725_LC_14_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_725_LC_14_3_2  (
            .in0(N__45078),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40475),
            .lcout(\c0.n6_adj_2430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_433_LC_14_3_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_433_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_433_LC_14_3_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_433_LC_14_3_3  (
            .in0(N__41817),
            .in1(N__37860),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17777 ),
            .ltout(\c0.n17777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_726_LC_14_3_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_726_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_726_LC_14_3_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_726_LC_14_3_4  (
            .in0(N__50672),
            .in1(N__37812),
            .in2(N__37806),
            .in3(N__44513),
            .lcout(\c0.n10617 ),
            .ltout(\c0.n10617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_731_LC_14_3_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_731_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_731_LC_14_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_731_LC_14_3_5  (
            .in0(_gnd_net_),
            .in1(N__37803),
            .in2(N__37764),
            .in3(N__41577),
            .lcout(\c0.n17765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_723_LC_14_3_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_723_LC_14_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_723_LC_14_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_723_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(N__37742),
            .in2(_gnd_net_),
            .in3(N__44375),
            .lcout(\c0.n17853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i60_LC_14_4_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i60_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i60_LC_14_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i60_LC_14_4_0  (
            .in0(N__41454),
            .in1(N__45107),
            .in2(_gnd_net_),
            .in3(N__50356),
            .lcout(data_out_frame2_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i95_LC_14_4_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i95_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i95_LC_14_4_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i95_LC_14_4_1  (
            .in0(N__50360),
            .in1(N__39278),
            .in2(_gnd_net_),
            .in3(N__41322),
            .lcout(data_out_frame2_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i118_LC_14_4_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i118_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i118_LC_14_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i118_LC_14_4_2  (
            .in0(N__38839),
            .in1(N__43603),
            .in2(_gnd_net_),
            .in3(N__50354),
            .lcout(data_out_frame2_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i80_LC_14_4_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i80_LC_14_4_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i80_LC_14_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i80_LC_14_4_3  (
            .in0(N__50359),
            .in1(N__40097),
            .in2(_gnd_net_),
            .in3(N__41149),
            .lcout(data_out_frame2_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i75_LC_14_4_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i75_LC_14_4_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i75_LC_14_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i75_LC_14_4_4  (
            .in0(N__39424),
            .in1(N__46594),
            .in2(_gnd_net_),
            .in3(N__50357),
            .lcout(data_out_frame2_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i79_LC_14_4_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i79_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i79_LC_14_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i79_LC_14_4_5  (
            .in0(N__50358),
            .in1(N__40147),
            .in2(_gnd_net_),
            .in3(N__40576),
            .lcout(data_out_frame2_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i119_LC_14_4_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i119_LC_14_4_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i119_LC_14_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i119_LC_14_4_6  (
            .in0(N__39704),
            .in1(N__43699),
            .in2(_gnd_net_),
            .in3(N__50355),
            .lcout(data_out_frame2_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15819_LC_14_4_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15819_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15819_LC_14_4_7 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15819_LC_14_4_7  (
            .in0(N__43602),
            .in1(N__46161),
            .in2(N__48691),
            .in3(N__45410),
            .lcout(\c0.n18681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i0_LC_14_5_0.C_ON=1'b1;
    defparam rand_data_2481__i0_LC_14_5_0.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i0_LC_14_5_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i0_LC_14_5_0 (
            .in0(_gnd_net_),
            .in1(N__38369),
            .in2(_gnd_net_),
            .in3(N__37914),
            .lcout(rand_data_0),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(n16547),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i1_LC_14_5_1.C_ON=1'b1;
    defparam rand_data_2481__i1_LC_14_5_1.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i1_LC_14_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i1_LC_14_5_1 (
            .in0(_gnd_net_),
            .in1(N__38309),
            .in2(_gnd_net_),
            .in3(N__37911),
            .lcout(rand_data_1),
            .ltout(),
            .carryin(n16547),
            .carryout(n16548),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i2_LC_14_5_2.C_ON=1'b1;
    defparam rand_data_2481__i2_LC_14_5_2.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i2_LC_14_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i2_LC_14_5_2 (
            .in0(_gnd_net_),
            .in1(N__38251),
            .in2(_gnd_net_),
            .in3(N__37956),
            .lcout(rand_data_2),
            .ltout(),
            .carryin(n16548),
            .carryout(n16549),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i3_LC_14_5_3.C_ON=1'b1;
    defparam rand_data_2481__i3_LC_14_5_3.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i3_LC_14_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i3_LC_14_5_3 (
            .in0(_gnd_net_),
            .in1(N__38164),
            .in2(_gnd_net_),
            .in3(N__37953),
            .lcout(rand_data_3),
            .ltout(),
            .carryin(n16549),
            .carryout(n16550),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i4_LC_14_5_4.C_ON=1'b1;
    defparam rand_data_2481__i4_LC_14_5_4.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i4_LC_14_5_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i4_LC_14_5_4 (
            .in0(_gnd_net_),
            .in1(N__38082),
            .in2(_gnd_net_),
            .in3(N__37950),
            .lcout(rand_data_4),
            .ltout(),
            .carryin(n16550),
            .carryout(n16551),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i5_LC_14_5_5.C_ON=1'b1;
    defparam rand_data_2481__i5_LC_14_5_5.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i5_LC_14_5_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i5_LC_14_5_5 (
            .in0(_gnd_net_),
            .in1(N__44203),
            .in2(_gnd_net_),
            .in3(N__37947),
            .lcout(rand_data_5),
            .ltout(),
            .carryin(n16551),
            .carryout(n16552),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i6_LC_14_5_6.C_ON=1'b1;
    defparam rand_data_2481__i6_LC_14_5_6.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i6_LC_14_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i6_LC_14_5_6 (
            .in0(_gnd_net_),
            .in1(N__41258),
            .in2(_gnd_net_),
            .in3(N__37944),
            .lcout(rand_data_6),
            .ltout(),
            .carryin(n16552),
            .carryout(n16553),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i7_LC_14_5_7.C_ON=1'b1;
    defparam rand_data_2481__i7_LC_14_5_7.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i7_LC_14_5_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i7_LC_14_5_7 (
            .in0(_gnd_net_),
            .in1(N__42080),
            .in2(_gnd_net_),
            .in3(N__37941),
            .lcout(rand_data_7),
            .ltout(),
            .carryin(n16553),
            .carryout(n16554),
            .clk(N__49871),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i8_LC_14_6_0.C_ON=1'b1;
    defparam rand_data_2481__i8_LC_14_6_0.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i8_LC_14_6_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i8_LC_14_6_0 (
            .in0(_gnd_net_),
            .in1(N__38693),
            .in2(_gnd_net_),
            .in3(N__37938),
            .lcout(rand_data_8),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(n16555),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i9_LC_14_6_1.C_ON=1'b1;
    defparam rand_data_2481__i9_LC_14_6_1.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i9_LC_14_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i9_LC_14_6_1 (
            .in0(_gnd_net_),
            .in1(N__38626),
            .in2(_gnd_net_),
            .in3(N__37935),
            .lcout(rand_data_9),
            .ltout(),
            .carryin(n16555),
            .carryout(n16556),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i10_LC_14_6_2.C_ON=1'b1;
    defparam rand_data_2481__i10_LC_14_6_2.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i10_LC_14_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i10_LC_14_6_2 (
            .in0(_gnd_net_),
            .in1(N__38542),
            .in2(_gnd_net_),
            .in3(N__37932),
            .lcout(rand_data_10),
            .ltout(),
            .carryin(n16556),
            .carryout(n16557),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i11_LC_14_6_3.C_ON=1'b1;
    defparam rand_data_2481__i11_LC_14_6_3.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i11_LC_14_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i11_LC_14_6_3 (
            .in0(_gnd_net_),
            .in1(N__41446),
            .in2(_gnd_net_),
            .in3(N__37983),
            .lcout(rand_data_11),
            .ltout(),
            .carryin(n16557),
            .carryout(n16558),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i12_LC_14_6_4.C_ON=1'b1;
    defparam rand_data_2481__i12_LC_14_6_4.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i12_LC_14_6_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i12_LC_14_6_4 (
            .in0(_gnd_net_),
            .in1(N__50504),
            .in2(_gnd_net_),
            .in3(N__37980),
            .lcout(rand_data_12),
            .ltout(),
            .carryin(n16558),
            .carryout(n16559),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i13_LC_14_6_5.C_ON=1'b1;
    defparam rand_data_2481__i13_LC_14_6_5.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i13_LC_14_6_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i13_LC_14_6_5 (
            .in0(_gnd_net_),
            .in1(N__38441),
            .in2(_gnd_net_),
            .in3(N__37977),
            .lcout(rand_data_13),
            .ltout(),
            .carryin(n16559),
            .carryout(n16560),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i14_LC_14_6_6.C_ON=1'b1;
    defparam rand_data_2481__i14_LC_14_6_6.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i14_LC_14_6_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i14_LC_14_6_6 (
            .in0(_gnd_net_),
            .in1(N__39265),
            .in2(_gnd_net_),
            .in3(N__37974),
            .lcout(rand_data_14),
            .ltout(),
            .carryin(n16560),
            .carryout(n16561),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i15_LC_14_6_7.C_ON=1'b1;
    defparam rand_data_2481__i15_LC_14_6_7.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i15_LC_14_6_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i15_LC_14_6_7 (
            .in0(_gnd_net_),
            .in1(N__39207),
            .in2(_gnd_net_),
            .in3(N__37971),
            .lcout(rand_data_15),
            .ltout(),
            .carryin(n16561),
            .carryout(n16562),
            .clk(N__49863),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i16_LC_14_7_0.C_ON=1'b1;
    defparam rand_data_2481__i16_LC_14_7_0.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i16_LC_14_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i16_LC_14_7_0 (
            .in0(_gnd_net_),
            .in1(N__39135),
            .in2(_gnd_net_),
            .in3(N__37968),
            .lcout(rand_data_16),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(n16563),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i17_LC_14_7_1.C_ON=1'b1;
    defparam rand_data_2481__i17_LC_14_7_1.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i17_LC_14_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i17_LC_14_7_1 (
            .in0(_gnd_net_),
            .in1(N__39055),
            .in2(_gnd_net_),
            .in3(N__37965),
            .lcout(rand_data_17),
            .ltout(),
            .carryin(n16563),
            .carryout(n16564),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i18_LC_14_7_2.C_ON=1'b1;
    defparam rand_data_2481__i18_LC_14_7_2.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i18_LC_14_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i18_LC_14_7_2 (
            .in0(_gnd_net_),
            .in1(N__40869),
            .in2(_gnd_net_),
            .in3(N__37962),
            .lcout(rand_data_18),
            .ltout(),
            .carryin(n16564),
            .carryout(n16565),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i19_LC_14_7_3.C_ON=1'b1;
    defparam rand_data_2481__i19_LC_14_7_3.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i19_LC_14_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i19_LC_14_7_3 (
            .in0(_gnd_net_),
            .in1(N__38960),
            .in2(_gnd_net_),
            .in3(N__37959),
            .lcout(rand_data_19),
            .ltout(),
            .carryin(n16565),
            .carryout(n16566),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i20_LC_14_7_4.C_ON=1'b1;
    defparam rand_data_2481__i20_LC_14_7_4.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i20_LC_14_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i20_LC_14_7_4 (
            .in0(_gnd_net_),
            .in1(N__38891),
            .in2(_gnd_net_),
            .in3(N__38010),
            .lcout(rand_data_20),
            .ltout(),
            .carryin(n16566),
            .carryout(n16567),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i21_LC_14_7_5.C_ON=1'b1;
    defparam rand_data_2481__i21_LC_14_7_5.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i21_LC_14_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i21_LC_14_7_5 (
            .in0(_gnd_net_),
            .in1(N__38816),
            .in2(_gnd_net_),
            .in3(N__38007),
            .lcout(rand_data_21),
            .ltout(),
            .carryin(n16567),
            .carryout(n16568),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i22_LC_14_7_6.C_ON=1'b1;
    defparam rand_data_2481__i22_LC_14_7_6.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i22_LC_14_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i22_LC_14_7_6 (
            .in0(_gnd_net_),
            .in1(N__39680),
            .in2(_gnd_net_),
            .in3(N__38004),
            .lcout(rand_data_22),
            .ltout(),
            .carryin(n16568),
            .carryout(n16569),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i23_LC_14_7_7.C_ON=1'b1;
    defparam rand_data_2481__i23_LC_14_7_7.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i23_LC_14_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i23_LC_14_7_7 (
            .in0(_gnd_net_),
            .in1(N__39602),
            .in2(_gnd_net_),
            .in3(N__38001),
            .lcout(rand_data_23),
            .ltout(),
            .carryin(n16569),
            .carryout(n16570),
            .clk(N__49857),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i24_LC_14_8_0.C_ON=1'b1;
    defparam rand_data_2481__i24_LC_14_8_0.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i24_LC_14_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i24_LC_14_8_0 (
            .in0(_gnd_net_),
            .in1(N__39539),
            .in2(_gnd_net_),
            .in3(N__37998),
            .lcout(rand_data_24),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(n16571),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i25_LC_14_8_1.C_ON=1'b1;
    defparam rand_data_2481__i25_LC_14_8_1.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i25_LC_14_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i25_LC_14_8_1 (
            .in0(_gnd_net_),
            .in1(N__39477),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(rand_data_25),
            .ltout(),
            .carryin(n16571),
            .carryout(n16572),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i26_LC_14_8_2.C_ON=1'b1;
    defparam rand_data_2481__i26_LC_14_8_2.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i26_LC_14_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i26_LC_14_8_2 (
            .in0(_gnd_net_),
            .in1(N__39411),
            .in2(_gnd_net_),
            .in3(N__37992),
            .lcout(rand_data_26),
            .ltout(),
            .carryin(n16572),
            .carryout(n16573),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i27_LC_14_8_3.C_ON=1'b1;
    defparam rand_data_2481__i27_LC_14_8_3.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i27_LC_14_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i27_LC_14_8_3 (
            .in0(_gnd_net_),
            .in1(N__42128),
            .in2(_gnd_net_),
            .in3(N__37989),
            .lcout(rand_data_27),
            .ltout(),
            .carryin(n16573),
            .carryout(n16574),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i28_LC_14_8_4.C_ON=1'b1;
    defparam rand_data_2481__i28_LC_14_8_4.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i28_LC_14_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i28_LC_14_8_4 (
            .in0(_gnd_net_),
            .in1(N__41478),
            .in2(_gnd_net_),
            .in3(N__37986),
            .lcout(rand_data_28),
            .ltout(),
            .carryin(n16574),
            .carryout(n16575),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i29_LC_14_8_5.C_ON=1'b1;
    defparam rand_data_2481__i29_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i29_LC_14_8_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i29_LC_14_8_5 (
            .in0(_gnd_net_),
            .in1(N__39325),
            .in2(_gnd_net_),
            .in3(N__38409),
            .lcout(rand_data_29),
            .ltout(),
            .carryin(n16575),
            .carryout(n16576),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i30_LC_14_8_6.C_ON=1'b1;
    defparam rand_data_2481__i30_LC_14_8_6.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i30_LC_14_8_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i30_LC_14_8_6 (
            .in0(_gnd_net_),
            .in1(N__40125),
            .in2(_gnd_net_),
            .in3(N__38406),
            .lcout(rand_data_30),
            .ltout(),
            .carryin(n16576),
            .carryout(n16577),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2481__i31_LC_14_8_7.C_ON=1'b0;
    defparam rand_data_2481__i31_LC_14_8_7.SEQ_MODE=4'b1000;
    defparam rand_data_2481__i31_LC_14_8_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2481__i31_LC_14_8_7 (
            .in0(_gnd_net_),
            .in1(N__40076),
            .in2(_gnd_net_),
            .in3(N__38403),
            .lcout(rand_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49850),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i0_LC_14_9_0.C_ON=1'b1;
    defparam rand_setpoint_2482__i0_LC_14_9_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i0_LC_14_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i0_LC_14_9_0 (
            .in0(_gnd_net_),
            .in1(N__38381),
            .in2(N__50945),
            .in3(_gnd_net_),
            .lcout(rand_setpoint_0),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(n16578),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i1_LC_14_9_1.C_ON=1'b1;
    defparam rand_setpoint_2482__i1_LC_14_9_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i1_LC_14_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i1_LC_14_9_1 (
            .in0(_gnd_net_),
            .in1(N__38316),
            .in2(N__40010),
            .in3(N__38280),
            .lcout(rand_setpoint_1),
            .ltout(),
            .carryin(n16578),
            .carryout(n16579),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i2_LC_14_9_2.C_ON=1'b1;
    defparam rand_setpoint_2482__i2_LC_14_9_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i2_LC_14_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i2_LC_14_9_2 (
            .in0(_gnd_net_),
            .in1(N__38261),
            .in2(N__38207),
            .in3(N__38190),
            .lcout(rand_setpoint_2),
            .ltout(),
            .carryin(n16579),
            .carryout(n16580),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i3_LC_14_9_3.C_ON=1'b1;
    defparam rand_setpoint_2482__i3_LC_14_9_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i3_LC_14_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i3_LC_14_9_3 (
            .in0(_gnd_net_),
            .in1(N__38175),
            .in2(N__38129),
            .in3(N__38112),
            .lcout(rand_setpoint_3),
            .ltout(),
            .carryin(n16580),
            .carryout(n16581),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i4_LC_14_9_4.C_ON=1'b1;
    defparam rand_setpoint_2482__i4_LC_14_9_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i4_LC_14_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i4_LC_14_9_4 (
            .in0(_gnd_net_),
            .in1(N__38048),
            .in2(N__38090),
            .in3(N__38037),
            .lcout(rand_setpoint_4),
            .ltout(),
            .carryin(n16581),
            .carryout(n16582),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i5_LC_14_9_5.C_ON=1'b1;
    defparam rand_setpoint_2482__i5_LC_14_9_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i5_LC_14_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i5_LC_14_9_5 (
            .in0(_gnd_net_),
            .in1(N__38024),
            .in2(N__44228),
            .in3(N__38013),
            .lcout(rand_setpoint_5),
            .ltout(),
            .carryin(n16582),
            .carryout(n16583),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i6_LC_14_9_6.C_ON=1'b1;
    defparam rand_setpoint_2482__i6_LC_14_9_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i6_LC_14_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i6_LC_14_9_6 (
            .in0(_gnd_net_),
            .in1(N__38762),
            .in2(N__41280),
            .in3(N__38751),
            .lcout(rand_setpoint_6),
            .ltout(),
            .carryin(n16583),
            .carryout(n16584),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i7_LC_14_9_7.C_ON=1'b1;
    defparam rand_setpoint_2482__i7_LC_14_9_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i7_LC_14_9_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i7_LC_14_9_7 (
            .in0(_gnd_net_),
            .in1(N__38738),
            .in2(N__42097),
            .in3(N__38727),
            .lcout(rand_setpoint_7),
            .ltout(),
            .carryin(n16584),
            .carryout(n16585),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i8_LC_14_10_0.C_ON=1'b1;
    defparam rand_setpoint_2482__i8_LC_14_10_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i8_LC_14_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i8_LC_14_10_0 (
            .in0(_gnd_net_),
            .in1(N__38702),
            .in2(N__43169),
            .in3(N__38664),
            .lcout(rand_setpoint_8),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(n16586),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i9_LC_14_10_1.C_ON=1'b1;
    defparam rand_setpoint_2482__i9_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i9_LC_14_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i9_LC_14_10_1 (
            .in0(_gnd_net_),
            .in1(N__38649),
            .in2(N__38588),
            .in3(N__38571),
            .lcout(rand_setpoint_9),
            .ltout(),
            .carryin(n16586),
            .carryout(n16587),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i10_LC_14_10_2.C_ON=1'b1;
    defparam rand_setpoint_2482__i10_LC_14_10_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i10_LC_14_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i10_LC_14_10_2 (
            .in0(_gnd_net_),
            .in1(N__38552),
            .in2(N__38508),
            .in3(N__38493),
            .lcout(rand_setpoint_10),
            .ltout(),
            .carryin(n16587),
            .carryout(n16588),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i11_LC_14_10_3.C_ON=1'b1;
    defparam rand_setpoint_2482__i11_LC_14_10_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i11_LC_14_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i11_LC_14_10_3 (
            .in0(_gnd_net_),
            .in1(N__41453),
            .in2(N__42888),
            .in3(N__38490),
            .lcout(rand_setpoint_11),
            .ltout(),
            .carryin(n16588),
            .carryout(n16589),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i12_LC_14_10_4.C_ON=1'b1;
    defparam rand_setpoint_2482__i12_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i12_LC_14_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i12_LC_14_10_4 (
            .in0(_gnd_net_),
            .in1(N__50523),
            .in2(N__38480),
            .in3(N__38463),
            .lcout(rand_setpoint_12),
            .ltout(),
            .carryin(n16589),
            .carryout(n16590),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i13_LC_14_10_5.C_ON=1'b1;
    defparam rand_setpoint_2482__i13_LC_14_10_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i13_LC_14_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i13_LC_14_10_5 (
            .in0(_gnd_net_),
            .in1(N__38449),
            .in2(N__40040),
            .in3(N__38412),
            .lcout(rand_setpoint_13),
            .ltout(),
            .carryin(n16590),
            .carryout(n16591),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i14_LC_14_10_6.C_ON=1'b1;
    defparam rand_setpoint_2482__i14_LC_14_10_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i14_LC_14_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i14_LC_14_10_6 (
            .in0(_gnd_net_),
            .in1(N__39283),
            .in2(N__47915),
            .in3(N__39237),
            .lcout(rand_setpoint_14),
            .ltout(),
            .carryin(n16591),
            .carryout(n16592),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i15_LC_14_10_7.C_ON=1'b1;
    defparam rand_setpoint_2482__i15_LC_14_10_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i15_LC_14_10_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i15_LC_14_10_7 (
            .in0(_gnd_net_),
            .in1(N__39173),
            .in2(N__39230),
            .in3(N__39162),
            .lcout(rand_setpoint_15),
            .ltout(),
            .carryin(n16592),
            .carryout(n16593),
            .clk(N__49831),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i16_LC_14_11_0.C_ON=1'b1;
    defparam rand_setpoint_2482__i16_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i16_LC_14_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i16_LC_14_11_0 (
            .in0(_gnd_net_),
            .in1(N__39148),
            .in2(N__39107),
            .in3(N__39090),
            .lcout(rand_setpoint_16),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(n16594),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i17_LC_14_11_1.C_ON=1'b1;
    defparam rand_setpoint_2482__i17_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i17_LC_14_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i17_LC_14_11_1 (
            .in0(_gnd_net_),
            .in1(N__39070),
            .in2(N__39026),
            .in3(N__39009),
            .lcout(rand_setpoint_17),
            .ltout(),
            .carryin(n16594),
            .carryout(n16595),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i18_LC_14_11_2.C_ON=1'b1;
    defparam rand_setpoint_2482__i18_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i18_LC_14_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i18_LC_14_11_2 (
            .in0(_gnd_net_),
            .in1(N__40876),
            .in2(N__39002),
            .in3(N__38985),
            .lcout(rand_setpoint_18),
            .ltout(),
            .carryin(n16595),
            .carryout(n16596),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i19_LC_14_11_3.C_ON=1'b1;
    defparam rand_setpoint_2482__i19_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i19_LC_14_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i19_LC_14_11_3 (
            .in0(_gnd_net_),
            .in1(N__38979),
            .in2(N__38927),
            .in3(N__38910),
            .lcout(rand_setpoint_19),
            .ltout(),
            .carryin(n16596),
            .carryout(n16597),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i20_LC_14_11_4.C_ON=1'b1;
    defparam rand_setpoint_2482__i20_LC_14_11_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i20_LC_14_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i20_LC_14_11_4 (
            .in0(_gnd_net_),
            .in1(N__38906),
            .in2(N__38865),
            .in3(N__38850),
            .lcout(rand_setpoint_20),
            .ltout(),
            .carryin(n16597),
            .carryout(n16598),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i21_LC_14_11_5.C_ON=1'b1;
    defparam rand_setpoint_2482__i21_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i21_LC_14_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i21_LC_14_11_5 (
            .in0(_gnd_net_),
            .in1(N__38838),
            .in2(N__38790),
            .in3(N__38775),
            .lcout(rand_setpoint_21),
            .ltout(),
            .carryin(n16598),
            .carryout(n16599),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i22_LC_14_11_6.C_ON=1'b1;
    defparam rand_setpoint_2482__i22_LC_14_11_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i22_LC_14_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i22_LC_14_11_6 (
            .in0(_gnd_net_),
            .in1(N__39699),
            .in2(N__39653),
            .in3(N__39636),
            .lcout(rand_setpoint_22),
            .ltout(),
            .carryin(n16599),
            .carryout(n16600),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i23_LC_14_11_7.C_ON=1'b1;
    defparam rand_setpoint_2482__i23_LC_14_11_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i23_LC_14_11_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i23_LC_14_11_7 (
            .in0(_gnd_net_),
            .in1(N__39624),
            .in2(N__39575),
            .in3(N__39558),
            .lcout(rand_setpoint_23),
            .ltout(),
            .carryin(n16600),
            .carryout(n16601),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i24_LC_14_12_0.C_ON=1'b1;
    defparam rand_setpoint_2482__i24_LC_14_12_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i24_LC_14_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i24_LC_14_12_0 (
            .in0(_gnd_net_),
            .in1(N__39553),
            .in2(N__42513),
            .in3(N__39513),
            .lcout(rand_setpoint_24),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(n16602),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i25_LC_14_12_1.C_ON=1'b1;
    defparam rand_setpoint_2482__i25_LC_14_12_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i25_LC_14_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i25_LC_14_12_1 (
            .in0(_gnd_net_),
            .in1(N__39492),
            .in2(N__39446),
            .in3(N__39429),
            .lcout(rand_setpoint_25),
            .ltout(),
            .carryin(n16602),
            .carryout(n16603),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i26_LC_14_12_2.C_ON=1'b1;
    defparam rand_setpoint_2482__i26_LC_14_12_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i26_LC_14_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i26_LC_14_12_2 (
            .in0(_gnd_net_),
            .in1(N__39415),
            .in2(N__39854),
            .in3(N__39387),
            .lcout(rand_setpoint_26),
            .ltout(),
            .carryin(n16603),
            .carryout(n16604),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i27_LC_14_12_3.C_ON=1'b1;
    defparam rand_setpoint_2482__i27_LC_14_12_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i27_LC_14_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i27_LC_14_12_3 (
            .in0(_gnd_net_),
            .in1(N__42138),
            .in2(N__39773),
            .in3(N__39384),
            .lcout(rand_setpoint_27),
            .ltout(),
            .carryin(n16604),
            .carryout(n16605),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i28_LC_14_12_4.C_ON=1'b1;
    defparam rand_setpoint_2482__i28_LC_14_12_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i28_LC_14_12_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i28_LC_14_12_4 (
            .in0(_gnd_net_),
            .in1(N__41499),
            .in2(N__39374),
            .in3(N__39357),
            .lcout(rand_setpoint_28),
            .ltout(),
            .carryin(n16605),
            .carryout(n16606),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i29_LC_14_12_5.C_ON=1'b1;
    defparam rand_setpoint_2482__i29_LC_14_12_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i29_LC_14_12_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i29_LC_14_12_5 (
            .in0(_gnd_net_),
            .in1(N__39342),
            .in2(N__39306),
            .in3(N__39291),
            .lcout(rand_setpoint_29),
            .ltout(),
            .carryin(n16606),
            .carryout(n16607),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i30_LC_14_12_6.C_ON=1'b1;
    defparam rand_setpoint_2482__i30_LC_14_12_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i30_LC_14_12_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2482__i30_LC_14_12_6 (
            .in0(_gnd_net_),
            .in1(N__40146),
            .in2(N__39791),
            .in3(N__40101),
            .lcout(rand_setpoint_30),
            .ltout(),
            .carryin(n16607),
            .carryout(n16608),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2482__i31_LC_14_12_7.C_ON=1'b0;
    defparam rand_setpoint_2482__i31_LC_14_12_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2482__i31_LC_14_12_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rand_setpoint_2482__i31_LC_14_12_7 (
            .in0(N__40092),
            .in1(N__43545),
            .in2(_gnd_net_),
            .in3(N__40044),
            .lcout(rand_setpoint_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49808),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5__2195_LC_14_13_2 .C_ON=1'b0;
    defparam \c0.data_out_7__5__2195_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5__2195_LC_14_13_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__5__2195_LC_14_13_2  (
            .in0(N__39931),
            .in1(N__40041),
            .in2(N__47799),
            .in3(N__47886),
            .lcout(\c0.data_out_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15534_3_lut_LC_14_13_3 .C_ON=1'b0;
    defparam \c0.i15534_3_lut_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15534_3_lut_LC_14_13_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15534_3_lut_LC_14_13_3  (
            .in0(N__47661),
            .in1(N__39743),
            .in2(_gnd_net_),
            .in3(N__39822),
            .lcout(\c0.n18234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__1__2191_LC_14_13_4 .C_ON=1'b0;
    defparam \c0.data_out_8__1__2191_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__1__2191_LC_14_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__1__2191_LC_14_13_4  (
            .in0(N__46814),
            .in1(N__40011),
            .in2(_gnd_net_),
            .in3(N__39972),
            .lcout(\c0.data_out_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49796),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_562_LC_14_13_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_562_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_562_LC_14_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_562_LC_14_13_6  (
            .in0(N__39930),
            .in1(N__47735),
            .in2(_gnd_net_),
            .in3(N__39909),
            .lcout(\c0.n10533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2__2214_LC_14_14_1 .C_ON=1'b0;
    defparam \c0.data_out_5__2__2214_LC_14_14_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__2__2214_LC_14_14_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.data_out_5__2__2214_LC_14_14_1  (
            .in0(N__47407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39855),
            .lcout(\c0.data_out_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49783),
            .ce(N__43418),
            .sr(N__43477));
    defparam \c0.data_out_5__6__2210_LC_14_14_2 .C_ON=1'b0;
    defparam \c0.data_out_5__6__2210_LC_14_14_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__6__2210_LC_14_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__6__2210_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__39792),
            .in2(_gnd_net_),
            .in3(N__47409),
            .lcout(\c0.data_out_7__2__N_447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49783),
            .ce(N__43418),
            .sr(N__43477));
    defparam \c0.data_out_5__3__2213_LC_14_14_4 .C_ON=1'b0;
    defparam \c0.data_out_5__3__2213_LC_14_14_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__3__2213_LC_14_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__3__2213_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__39774),
            .in2(_gnd_net_),
            .in3(N__47408),
            .lcout(\c0.data_out_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49783),
            .ce(N__43418),
            .sr(N__43477));
    defparam \c0.data_out_10__4__2172_LC_14_15_0 .C_ON=1'b0;
    defparam \c0.data_out_10__4__2172_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__4__2172_LC_14_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_10__4__2172_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__40341),
            .in2(_gnd_net_),
            .in3(N__40323),
            .lcout(\c0.data_out_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49768),
            .ce(N__46857),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__0__2232_LC_14_16_0 .C_ON=1'b0;
    defparam \c0.data_out_3__0__2232_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0__2232_LC_14_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_3__0__2232_LC_14_16_0  (
            .in0(N__40245),
            .in1(N__40281),
            .in2(_gnd_net_),
            .in3(N__43395),
            .lcout(data_out_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_14_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_14_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_14_16_4  (
            .in0(N__40244),
            .in1(N__40226),
            .in2(_gnd_net_),
            .in3(N__42862),
            .lcout(\c0.n2_adj_2221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__0__2240_LC_14_16_5 .C_ON=1'b0;
    defparam \c0.data_out_2__0__2240_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__0__2240_LC_14_16_5 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_2__0__2240_LC_14_16_5  (
            .in0(N__40227),
            .in1(N__43394),
            .in2(_gnd_net_),
            .in3(N__47141),
            .lcout(data_out_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_15_1_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_15_1_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_15_1_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_15_1_0  (
            .in0(N__46164),
            .in1(N__40218),
            .in2(N__48702),
            .in3(N__41568),
            .lcout(\c0.n6_adj_2227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15874_LC_15_1_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15874_LC_15_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15874_LC_15_1_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15874_LC_15_1_1  (
            .in0(N__41763),
            .in1(N__43708),
            .in2(N__48700),
            .in3(N__46163),
            .lcout(\c0.n18705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_810_LC_15_1_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_810_LC_15_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_810_LC_15_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_810_LC_15_1_2  (
            .in0(N__45305),
            .in1(N__40949),
            .in2(_gnd_net_),
            .in3(N__40203),
            .lcout(\c0.n17899 ),
            .ltout(\c0.n17899_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_738_LC_15_1_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_738_LC_15_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_738_LC_15_1_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_738_LC_15_1_3  (
            .in0(N__41864),
            .in1(N__44010),
            .in2(N__40167),
            .in3(N__42180),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_796_LC_15_1_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_796_LC_15_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_796_LC_15_1_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_796_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(N__40840),
            .in2(_gnd_net_),
            .in3(N__44324),
            .lcout(\c0.n17736 ),
            .ltout(\c0.n17736_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_541_LC_15_1_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_541_LC_15_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_541_LC_15_1_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_541_LC_15_1_5  (
            .in0(N__41863),
            .in1(N__41218),
            .in2(N__40611),
            .in3(N__40587),
            .lcout(\c0.n17914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18813_bdd_4_lut_LC_15_1_6 .C_ON=1'b0;
    defparam \c0.n18813_bdd_4_lut_LC_15_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18813_bdd_4_lut_LC_15_1_6 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \c0.n18813_bdd_4_lut_LC_15_1_6  (
            .in0(N__42231),
            .in1(N__44268),
            .in2(N__48701),
            .in3(N__40608),
            .lcout(\c0.n18816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_501_LC_15_1_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_501_LC_15_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_501_LC_15_1_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_501_LC_15_1_7  (
            .in0(N__44325),
            .in1(_gnd_net_),
            .in2(N__40845),
            .in3(N__40588),
            .lcout(\c0.n10725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_683_LC_15_2_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_683_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_683_LC_15_2_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_683_LC_15_2_0  (
            .in0(N__40549),
            .in1(N__41883),
            .in2(N__40509),
            .in3(N__46308),
            .lcout(),
            .ltout(\c0.n17_adj_2413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i163_LC_15_2_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i163_LC_15_2_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i163_LC_15_2_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i163_LC_15_2_1  (
            .in0(N__43979),
            .in1(N__40491),
            .in2(N__40479),
            .in3(N__40371),
            .lcout(\c0.data_out_frame2_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49888),
            .ce(N__50462),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_681_LC_15_2_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_681_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_681_LC_15_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_681_LC_15_2_2  (
            .in0(N__40476),
            .in1(N__45267),
            .in2(N__40436),
            .in3(N__40407),
            .lcout(\c0.n17862 ),
            .ltout(\c0.n17862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_676_LC_15_2_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_676_LC_15_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_676_LC_15_2_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_676_LC_15_2_3  (
            .in0(N__40905),
            .in1(N__45536),
            .in2(N__40365),
            .in3(N__40362),
            .lcout(),
            .ltout(\c0.n12_adj_2410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i164_LC_15_2_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i164_LC_15_2_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i164_LC_15_2_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i164_LC_15_2_4  (
            .in0(N__41679),
            .in1(N__50553),
            .in2(N__40344),
            .in3(N__43776),
            .lcout(\c0.data_out_frame2_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49888),
            .ce(N__50462),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_719_LC_15_2_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_719_LC_15_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_719_LC_15_2_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_719_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__40992),
            .in2(_gnd_net_),
            .in3(N__40950),
            .lcout(\c0.n17889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_790_LC_15_3_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_790_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_790_LC_15_3_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_790_LC_15_3_0  (
            .in0(N__44099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41145),
            .lcout(\c0.n17868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i51_LC_15_3_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i51_LC_15_3_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i51_LC_15_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i51_LC_15_3_1  (
            .in0(N__40892),
            .in1(N__40839),
            .in2(_gnd_net_),
            .in3(N__50436),
            .lcout(data_out_frame2_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49885),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18645_bdd_4_lut_LC_15_3_2 .C_ON=1'b0;
    defparam \c0.n18645_bdd_4_lut_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18645_bdd_4_lut_LC_15_3_2 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.n18645_bdd_4_lut_LC_15_3_2  (
            .in0(N__43761),
            .in1(N__48686),
            .in2(N__46595),
            .in3(N__40815),
            .lcout(\c0.n18648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_770_LC_15_3_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_770_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_770_LC_15_3_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_770_LC_15_3_3  (
            .in0(N__45814),
            .in1(N__41331),
            .in2(N__44535),
            .in3(N__40787),
            .lcout(\c0.n18_adj_2441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18663_bdd_4_lut_LC_15_3_4 .C_ON=1'b0;
    defparam \c0.n18663_bdd_4_lut_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18663_bdd_4_lut_LC_15_3_4 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18663_bdd_4_lut_LC_15_3_4  (
            .in0(N__40786),
            .in1(N__41376),
            .in2(N__44581),
            .in3(N__48685),
            .lcout(\c0.n18666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_520_LC_15_3_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_520_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_520_LC_15_3_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_520_LC_15_3_5  (
            .in0(N__43610),
            .in1(_gnd_net_),
            .in2(N__43679),
            .in3(N__40752),
            .lcout(\c0.n17917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_740_LC_15_3_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_740_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_740_LC_15_3_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_740_LC_15_3_6  (
            .in0(N__40707),
            .in1(N__40688),
            .in2(N__41523),
            .in3(N__44523),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_15_4_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_15_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_15_4_0  (
            .in0(N__46191),
            .in1(N__40665),
            .in2(_gnd_net_),
            .in3(N__44690),
            .lcout(\c0.n5_adj_2439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15804_LC_15_4_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15804_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15804_LC_15_4_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15804_LC_15_4_1  (
            .in0(N__45625),
            .in1(N__41414),
            .in2(N__48693),
            .in3(N__46192),
            .lcout(\c0.n18663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_769_LC_15_4_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_769_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_769_LC_15_4_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_769_LC_15_4_2  (
            .in0(N__41370),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45015),
            .lcout(\c0.n10911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_772_LC_15_4_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_772_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_772_LC_15_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_772_LC_15_4_3  (
            .in0(N__50571),
            .in1(N__45244),
            .in2(_gnd_net_),
            .in3(N__41312),
            .lcout(\c0.n17810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i103_LC_15_4_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i103_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i103_LC_15_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i103_LC_15_4_4  (
            .in0(N__41262),
            .in1(N__43579),
            .in2(_gnd_net_),
            .in3(N__50446),
            .lcout(data_out_frame2_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i77_LC_15_4_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i77_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i77_LC_15_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i77_LC_15_4_5  (
            .in0(N__50447),
            .in1(N__41507),
            .in2(_gnd_net_),
            .in3(N__41217),
            .lcout(data_out_frame2_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_812_LC_15_4_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_812_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_812_LC_15_4_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_812_LC_15_4_6  (
            .in0(N__41185),
            .in1(N__44053),
            .in2(N__41150),
            .in3(N__44614),
            .lcout(\c0.n10703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i93_LC_15_4_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i93_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i93_LC_15_4_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i93_LC_15_4_7  (
            .in0(N__50448),
            .in1(_gnd_net_),
            .in2(N__50581),
            .in3(N__50525),
            .lcout(data_out_frame2_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_542_LC_15_5_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_542_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_542_LC_15_5_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_542_LC_15_5_0  (
            .in0(N__46590),
            .in1(N__46707),
            .in2(N__41121),
            .in3(N__43575),
            .lcout(\c0.n14_adj_2362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_522_LC_15_5_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_522_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_522_LC_15_5_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_522_LC_15_5_1  (
            .in0(N__46411),
            .in1(N__41567),
            .in2(N__41094),
            .in3(N__41037),
            .lcout(\c0.n17892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_728_LC_15_5_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_728_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_728_LC_15_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_728_LC_15_5_2  (
            .in0(N__46589),
            .in1(N__41901),
            .in2(_gnd_net_),
            .in3(N__41765),
            .lcout(\c0.n17789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_15_5_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_15_5_3 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_15_5_3  (
            .in0(N__41859),
            .in1(N__48609),
            .in2(N__41826),
            .in3(N__46193),
            .lcout(\c0.n6_adj_2218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_646_LC_15_5_4 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_646_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_646_LC_15_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_646_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(N__41816),
            .in2(_gnd_net_),
            .in3(N__41764),
            .lcout(\c0.n18_adj_2393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_730_LC_15_5_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_730_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_730_LC_15_5_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_730_LC_15_5_5  (
            .in0(N__41723),
            .in1(N__41670),
            .in2(N__41625),
            .in3(N__50821),
            .lcout(\c0.n10_adj_2431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_15_5_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_15_5_6 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_15_5_6  (
            .in0(N__46194),
            .in1(N__44067),
            .in2(N__48684),
            .in3(N__43855),
            .lcout(\c0.n6_adj_2360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_766_LC_15_5_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_766_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_766_LC_15_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_766_LC_15_5_7  (
            .in0(_gnd_net_),
            .in1(N__41566),
            .in2(_gnd_net_),
            .in3(N__50881),
            .lcout(\c0.n17865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i109_LC_15_6_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i109_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i109_LC_15_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i109_LC_15_6_0  (
            .in0(N__41500),
            .in1(N__42969),
            .in2(_gnd_net_),
            .in3(N__50453),
            .lcout(data_out_frame2_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i140_LC_15_6_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i140_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i140_LC_15_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i140_LC_15_6_1  (
            .in0(N__50454),
            .in1(N__41447),
            .in2(_gnd_net_),
            .in3(N__41973),
            .lcout(data_out_frame2_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_696_LC_15_6_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_696_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_696_LC_15_6_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_696_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__42230),
            .in2(_gnd_net_),
            .in3(N__41954),
            .lcout(\c0.n17902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_679_LC_15_6_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_679_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_679_LC_15_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_679_LC_15_6_3  (
            .in0(N__42201),
            .in1(N__44754),
            .in2(_gnd_net_),
            .in3(N__50820),
            .lcout(\c0.n10583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18705_bdd_4_lut_LC_15_6_4 .C_ON=1'b0;
    defparam \c0.n18705_bdd_4_lut_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18705_bdd_4_lut_LC_15_6_4 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18705_bdd_4_lut_LC_15_6_4  (
            .in0(N__48607),
            .in1(N__42192),
            .in2(N__43584),
            .in3(N__42173),
            .lcout(\c0.n18708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i76_LC_15_6_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i76_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i76_LC_15_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i76_LC_15_6_5  (
            .in0(N__50455),
            .in1(N__42149),
            .in2(_gnd_net_),
            .in3(N__44571),
            .lcout(data_out_frame2_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i104_LC_15_6_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i104_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i104_LC_15_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i104_LC_15_6_6  (
            .in0(N__42087),
            .in1(N__44267),
            .in2(_gnd_net_),
            .in3(N__50452),
            .lcout(data_out_frame2_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18657_bdd_4_lut_LC_15_6_7 .C_ON=1'b0;
    defparam \c0.n18657_bdd_4_lut_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18657_bdd_4_lut_LC_15_6_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18657_bdd_4_lut_LC_15_6_7  (
            .in0(N__42053),
            .in1(N__48608),
            .in2(N__43821),
            .in3(N__42015),
            .lcout(\c0.n18660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15794_LC_15_7_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15794_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15794_LC_15_7_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15794_LC_15_7_0  (
            .in0(N__42003),
            .in1(N__48618),
            .in2(N__41985),
            .in3(N__46159),
            .lcout(),
            .ltout(\c0.n18651_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18651_bdd_4_lut_LC_15_7_1 .C_ON=1'b0;
    defparam \c0.n18651_bdd_4_lut_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18651_bdd_4_lut_LC_15_7_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18651_bdd_4_lut_LC_15_7_1  (
            .in0(N__48619),
            .in1(N__41972),
            .in2(N__41961),
            .in3(N__41958),
            .lcout(),
            .ltout(\c0.n18654_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_15_7_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_15_7_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_15_7_2  (
            .in0(N__48076),
            .in1(N__41916),
            .in2(N__41904),
            .in3(N__48139),
            .lcout(\c0.n22_adj_2259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15859_LC_15_7_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15859_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15859_LC_15_7_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15859_LC_15_7_3  (
            .in0(N__42438),
            .in1(N__49097),
            .in2(N__42429),
            .in3(N__48077),
            .lcout(),
            .ltout(\c0.n18735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18735_bdd_4_lut_LC_15_7_4 .C_ON=1'b0;
    defparam \c0.n18735_bdd_4_lut_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18735_bdd_4_lut_LC_15_7_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18735_bdd_4_lut_LC_15_7_4  (
            .in0(N__49098),
            .in1(N__42417),
            .in2(N__42408),
            .in3(N__42405),
            .lcout(),
            .ltout(\c0.n18738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_15_7_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_15_7_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_15_7_5  (
            .in0(N__42396),
            .in1(N__49099),
            .in2(N__42390),
            .in3(N__48950),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49864),
            .ce(N__48828),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15833_LC_15_8_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15833_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15833_LC_15_8_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15833_LC_15_8_0  (
            .in0(N__46150),
            .in1(N__42372),
            .in2(N__43881),
            .in3(N__48402),
            .lcout(\c0.n18699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15943_LC_15_8_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15943_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15943_LC_15_8_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15943_LC_15_8_1  (
            .in0(N__42354),
            .in1(N__49094),
            .in2(N__42345),
            .in3(N__48079),
            .lcout(),
            .ltout(\c0.n18777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18777_bdd_4_lut_LC_15_8_2 .C_ON=1'b0;
    defparam \c0.n18777_bdd_4_lut_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18777_bdd_4_lut_LC_15_8_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18777_bdd_4_lut_LC_15_8_2  (
            .in0(N__49095),
            .in1(N__42327),
            .in2(N__42315),
            .in3(N__42312),
            .lcout(\c0.n18780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18699_bdd_4_lut_LC_15_8_3 .C_ON=1'b0;
    defparam \c0.n18699_bdd_4_lut_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18699_bdd_4_lut_LC_15_8_3 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18699_bdd_4_lut_LC_15_8_3  (
            .in0(N__48403),
            .in1(N__42303),
            .in2(N__42297),
            .in3(N__42276),
            .lcout(),
            .ltout(\c0.n18702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_15_8_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_15_8_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_15_8_4  (
            .in0(N__48080),
            .in1(N__44469),
            .in2(N__42234),
            .in3(N__48138),
            .lcout(),
            .ltout(\c0.n22_adj_2240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_15_8_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_15_8_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_15_8_5  (
            .in0(N__43002),
            .in1(N__49096),
            .in2(N__42996),
            .in3(N__48949),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49858),
            .ce(N__48824),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15899_LC_15_9_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15899_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15899_LC_15_9_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15899_LC_15_9_0  (
            .in0(N__48620),
            .in1(N__46080),
            .in2(N__44439),
            .in3(N__45013),
            .lcout(),
            .ltout(\c0.n18783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18783_bdd_4_lut_LC_15_9_1 .C_ON=1'b0;
    defparam \c0.n18783_bdd_4_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18783_bdd_4_lut_LC_15_9_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n18783_bdd_4_lut_LC_15_9_1  (
            .in0(N__45201),
            .in1(N__48621),
            .in2(N__42981),
            .in3(N__42976),
            .lcout(\c0.n18161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11016_2_lut_LC_15_9_4 .C_ON=1'b0;
    defparam \c0.i11016_2_lut_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11016_2_lut_LC_15_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i11016_2_lut_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__47399),
            .in2(_gnd_net_),
            .in3(N__47129),
            .lcout(n2732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15645_2_lut_LC_15_11_3 .C_ON=1'b0;
    defparam \c0.i15645_2_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15645_2_lut_LC_15_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15645_2_lut_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__42933),
            .in2(_gnd_net_),
            .in3(N__42863),
            .lcout(\c0.n18311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15532_2_lut_LC_15_11_4 .C_ON=1'b0;
    defparam \c0.i15532_2_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15532_2_lut_LC_15_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15532_2_lut_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__42887),
            .in2(_gnd_net_),
            .in3(N__47404),
            .lcout(\c0.n18201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_15_11_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_15_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_15_11_6  (
            .in0(N__42864),
            .in1(N__42524),
            .in2(_gnd_net_),
            .in3(N__42604),
            .lcout(\c0.n5_adj_2217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__3__2197_LC_15_12_7 .C_ON=1'b0;
    defparam \c0.data_out_7__3__2197_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3__2197_LC_15_12_7 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \c0.data_out_7__3__2197_LC_15_12_7  (
            .in0(N__47671),
            .in1(N__47130),
            .in2(N__42549),
            .in3(N__43514),
            .lcout(\c0.data_out_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49820),
            .ce(N__47893),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__0__2216_LC_15_13_0 .C_ON=1'b0;
    defparam \c0.data_out_5__0__2216_LC_15_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__0__2216_LC_15_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__0__2216_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__42512),
            .in2(_gnd_net_),
            .in3(N__47405),
            .lcout(\c0.data_out_6__1__N_537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49809),
            .ce(N__43417),
            .sr(N__43479));
    defparam \c0.data_out_5__7__2209_LC_15_13_3 .C_ON=1'b0;
    defparam \c0.data_out_5__7__2209_LC_15_13_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__7__2209_LC_15_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.data_out_5__7__2209_LC_15_13_3  (
            .in0(N__47406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43544),
            .lcout(\c0.data_out_7__3__N_441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49809),
            .ce(N__43417),
            .sr(N__43479));
    defparam \c0.data_out_1__1__2247_LC_15_14_4 .C_ON=1'b0;
    defparam \c0.data_out_1__1__2247_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__1__2247_LC_15_14_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \c0.data_out_1__1__2247_LC_15_14_4  (
            .in0(N__47676),
            .in1(N__47410),
            .in2(_gnd_net_),
            .in3(N__47144),
            .lcout(\c0.data_out_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49797),
            .ce(N__43419),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0__2200_LC_15_15_4 .C_ON=1'b0;
    defparam \c0.data_out_7__0__2200_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0__2200_LC_15_15_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__0__2200_LC_15_15_4  (
            .in0(N__43185),
            .in1(N__47411),
            .in2(N__43176),
            .in3(N__47145),
            .lcout(\c0.data_out_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49784),
            .ce(N__47884),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15884_LC_16_1_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15884_LC_16_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15884_LC_16_1_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15884_LC_16_1_1  (
            .in0(N__43122),
            .in1(N__49108),
            .in2(N__43113),
            .in3(N__48071),
            .lcout(),
            .ltout(\c0.n18765_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18765_bdd_4_lut_LC_16_1_2 .C_ON=1'b0;
    defparam \c0.n18765_bdd_4_lut_LC_16_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18765_bdd_4_lut_LC_16_1_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18765_bdd_4_lut_LC_16_1_2  (
            .in0(N__49109),
            .in1(N__43101),
            .in2(N__43089),
            .in3(N__43086),
            .lcout(),
            .ltout(\c0.n18768_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_16_1_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_16_1_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_16_1_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_16_1_3  (
            .in0(N__43989),
            .in1(N__49110),
            .in2(N__43077),
            .in3(N__48951),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49892),
            .ce(N__48811),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15779_LC_16_1_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15779_LC_16_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15779_LC_16_1_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15779_LC_16_1_4  (
            .in0(N__43056),
            .in1(N__48679),
            .in2(N__43038),
            .in3(N__46184),
            .lcout(),
            .ltout(\c0.n18633_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18633_bdd_4_lut_LC_16_1_5 .C_ON=1'b0;
    defparam \c0.n18633_bdd_4_lut_LC_16_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18633_bdd_4_lut_LC_16_1_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18633_bdd_4_lut_LC_16_1_5  (
            .in0(N__48680),
            .in1(N__43026),
            .in2(N__43005),
            .in3(N__46654),
            .lcout(),
            .ltout(\c0.n18636_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_16_1_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_16_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_16_1_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_16_1_6  (
            .in0(N__48070),
            .in1(N__43998),
            .in2(N__43992),
            .in3(N__48169),
            .lcout(\c0.n22_adj_2268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_753_LC_16_2_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_753_LC_16_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_753_LC_16_2_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_753_LC_16_2_1  (
            .in0(N__50763),
            .in1(N__43583),
            .in2(N__43983),
            .in3(N__43959),
            .lcout(),
            .ltout(\c0.n20_adj_2438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i159_LC_16_2_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i159_LC_16_2_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i159_LC_16_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i159_LC_16_2_2  (
            .in0(N__43911),
            .in1(N__43767),
            .in2(N__43902),
            .in3(N__43899),
            .lcout(\c0.data_out_frame2_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(N__50475),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_750_LC_16_2_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_750_LC_16_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_750_LC_16_2_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_750_LC_16_2_3  (
            .in0(N__43866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43820),
            .lcout(\c0.n10905 ),
            .ltout(\c0.n10905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_16_2_4 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_16_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_16_2_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_2_lut_3_lut_4_lut_LC_16_2_4  (
            .in0(N__44150),
            .in1(N__44284),
            .in2(N__43770),
            .in3(N__46486),
            .lcout(\c0.n16_adj_2391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_801_LC_16_2_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_801_LC_16_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_801_LC_16_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_801_LC_16_2_5  (
            .in0(N__43710),
            .in1(N__43760),
            .in2(_gnd_net_),
            .in3(N__45790),
            .lcout(\c0.n17920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_427_LC_16_2_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_427_LC_16_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_427_LC_16_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_427_LC_16_2_6  (
            .in0(N__45791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43709),
            .lcout(\c0.n10788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_756_LC_16_3_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_756_LC_16_3_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_756_LC_16_3_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_756_LC_16_3_0  (
            .in0(N__43680),
            .in1(N__43614),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_767_LC_16_3_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_767_LC_16_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_767_LC_16_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_767_LC_16_3_1  (
            .in0(_gnd_net_),
            .in1(N__43574),
            .in2(_gnd_net_),
            .in3(N__48221),
            .lcout(\c0.n10929 ),
            .ltout(\c0.n10929_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_734_LC_16_3_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_734_LC_16_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_734_LC_16_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_734_LC_16_3_2  (
            .in0(_gnd_net_),
            .in1(N__44857),
            .in2(N__44526),
            .in3(N__44928),
            .lcout(\c0.n17823 ),
            .ltout(\c0.n17823_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_656_LC_16_3_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_656_LC_16_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_656_LC_16_3_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_656_LC_16_3_3  (
            .in0(N__44433),
            .in1(N__44517),
            .in2(N__44502),
            .in3(N__46485),
            .lcout(),
            .ltout(\c0.n17_adj_2401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i167_LC_16_3_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i167_LC_16_3_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i167_LC_16_3_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i167_LC_16_3_4  (
            .in0(N__44499),
            .in1(N__46545),
            .in2(N__44493),
            .in3(N__44489),
            .lcout(\c0.data_out_frame2_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(N__50466),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_660_LC_16_3_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_660_LC_16_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_660_LC_16_3_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_660_LC_16_3_5  (
            .in0(N__44453),
            .in1(N__44582),
            .in2(N__44438),
            .in3(N__44388),
            .lcout(\c0.n18_adj_2402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_649_LC_16_3_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_649_LC_16_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_649_LC_16_3_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_649_LC_16_3_6  (
            .in0(N__44376),
            .in1(N__44331),
            .in2(N__44285),
            .in3(N__44858),
            .lcout(\c0.n22_adj_2395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i102_LC_16_4_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i102_LC_16_4_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i102_LC_16_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i102_LC_16_4_0  (
            .in0(N__44140),
            .in1(N__44230),
            .in2(_gnd_net_),
            .in3(N__50449),
            .lcout(data_out_frame2_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_16_4_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_16_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_16_4_1  (
            .in0(N__45115),
            .in1(N__44103),
            .in2(_gnd_net_),
            .in3(N__46196),
            .lcout(\c0.n5_adj_2381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_735_LC_16_4_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_735_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_735_LC_16_4_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_735_LC_16_4_2  (
            .in0(N__44900),
            .in1(N__46416),
            .in2(N__44061),
            .in3(N__45117),
            .lcout(\c0.n30_adj_2434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_667_LC_16_4_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_667_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_667_LC_16_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_667_LC_16_4_3  (
            .in0(N__45116),
            .in1(N__45093),
            .in2(_gnd_net_),
            .in3(N__45045),
            .lcout(\c0.n17871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_733_LC_16_4_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_733_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_733_LC_16_4_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_733_LC_16_4_4  (
            .in0(N__46353),
            .in1(N__45014),
            .in2(N__44971),
            .in3(N__45546),
            .lcout(\c0.n10710 ),
            .ltout(\c0.n10710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_662_LC_16_4_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_662_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_662_LC_16_4_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_662_LC_16_4_5  (
            .in0(N__44718),
            .in1(N__45287),
            .in2(N__44922),
            .in3(N__44919),
            .lcout(\c0.n20_adj_2404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_16_4_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_16_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_16_4_6  (
            .in0(N__46195),
            .in1(N__44901),
            .in2(_gnd_net_),
            .in3(N__44859),
            .lcout(\c0.n5_adj_2386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_764_LC_16_4_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_764_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_764_LC_16_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_764_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(N__44811),
            .in2(_gnd_net_),
            .in3(N__44753),
            .lcout(\c0.n10877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_16_5_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_16_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_16_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_711_LC_16_5_0  (
            .in0(N__45668),
            .in1(N__45621),
            .in2(_gnd_net_),
            .in3(N__45683),
            .lcout(),
            .ltout(\c0.n10593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_16_5_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_16_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__45380),
            .in2(N__44712),
            .in3(N__44697),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_729_LC_16_5_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_729_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_729_LC_16_5_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_729_LC_16_5_2  (
            .in0(N__44696),
            .in1(N__44661),
            .in2(N__44625),
            .in3(N__44564),
            .lcout(\c0.n17751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_534_LC_16_5_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_534_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_534_LC_16_5_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_534_LC_16_5_3  (
            .in0(N__45682),
            .in1(N__45667),
            .in2(N__45626),
            .in3(N__45576),
            .lcout(\c0.n17798 ),
            .ltout(\c0.n17798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_648_LC_16_5_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_648_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_648_LC_16_5_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_648_LC_16_5_4  (
            .in0(N__45523),
            .in1(N__45507),
            .in2(N__45489),
            .in3(N__45482),
            .lcout(),
            .ltout(\c0.n24_adj_2394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_651_LC_16_5_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_651_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_651_LC_16_5_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_651_LC_16_5_5  (
            .in0(N__45468),
            .in1(N__45462),
            .in2(N__45417),
            .in3(N__45414),
            .lcout(),
            .ltout(\c0.n26_adj_2396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i168_LC_16_5_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i168_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i168_LC_16_5_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i168_LC_16_5_6  (
            .in0(N__45381),
            .in1(N__45369),
            .in2(N__45360),
            .in3(N__45353),
            .lcout(\c0.data_out_frame2_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49882),
            .ce(N__50469),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_668_LC_16_6_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_668_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_668_LC_16_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_668_LC_16_6_2  (
            .in0(N__46656),
            .in1(_gnd_net_),
            .in2(N__50552),
            .in3(N__45315),
            .lcout(),
            .ltout(\c0.n14_adj_2406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i165_LC_16_6_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i165_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i165_LC_16_6_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i165_LC_16_6_3  (
            .in0(N__45288),
            .in1(N__46662),
            .in2(N__45270),
            .in3(N__45123),
            .lcout(\c0.data_out_frame2_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__50468),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_670_LC_16_6_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_670_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_670_LC_16_6_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_670_LC_16_6_4  (
            .in0(N__45263),
            .in1(N__45249),
            .in2(N__45207),
            .in3(N__45147),
            .lcout(\c0.n15_adj_2407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_685_LC_16_6_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_685_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_685_LC_16_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_685_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__46715),
            .in2(_gnd_net_),
            .in3(N__46604),
            .lcout(\c0.n17856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_654_LC_16_6_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_654_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_654_LC_16_6_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_654_LC_16_6_6  (
            .in0(N__46655),
            .in1(N__46536),
            .in2(N__46608),
            .in3(N__46563),
            .lcout(\c0.n16_adj_2399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15988_LC_16_7_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15988_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15988_LC_16_7_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15988_LC_16_7_0  (
            .in0(N__48694),
            .in1(N__46533),
            .in2(N__46488),
            .in3(N__46157),
            .lcout(),
            .ltout(\c0.n18891_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18891_bdd_4_lut_LC_16_7_1 .C_ON=1'b0;
    defparam \c0.n18891_bdd_4_lut_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18891_bdd_4_lut_LC_16_7_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18891_bdd_4_lut_LC_16_7_1  (
            .in0(N__48692),
            .in1(N__46410),
            .in2(N__46356),
            .in3(N__46352),
            .lcout(\c0.n18060 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_16_7_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_16_7_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_16_7_2  (
            .in0(N__48695),
            .in1(N__46304),
            .in2(N__46263),
            .in3(N__46158),
            .lcout(),
            .ltout(\c0.n18897_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18897_bdd_4_lut_LC_16_7_3 .C_ON=1'b0;
    defparam \c0.n18897_bdd_4_lut_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18897_bdd_4_lut_LC_16_7_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n18897_bdd_4_lut_LC_16_7_3  (
            .in0(N__45857),
            .in1(N__48696),
            .in2(N__45819),
            .in3(N__45816),
            .lcout(),
            .ltout(\c0.n18057_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15854_LC_16_7_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15854_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15854_LC_16_7_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15854_LC_16_7_4  (
            .in0(N__45732),
            .in1(N__49111),
            .in2(N__45726),
            .in3(N__48081),
            .lcout(),
            .ltout(\c0.n18723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18723_bdd_4_lut_LC_16_7_5 .C_ON=1'b0;
    defparam \c0.n18723_bdd_4_lut_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18723_bdd_4_lut_LC_16_7_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18723_bdd_4_lut_LC_16_7_5  (
            .in0(N__49112),
            .in1(N__45723),
            .in2(N__45714),
            .in3(N__45711),
            .lcout(),
            .ltout(\c0.n18726_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_16_7_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_16_7_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_16_7_6  (
            .in0(N__49200),
            .in1(N__49113),
            .in2(N__49182),
            .in3(N__48948),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49873),
            .ce(N__48816),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15889_LC_16_8_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15889_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15889_LC_16_8_3 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15889_LC_16_8_3  (
            .in0(N__49170),
            .in1(N__48078),
            .in2(N__49158),
            .in3(N__49114),
            .lcout(),
            .ltout(\c0.n18771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18771_bdd_4_lut_LC_16_8_4 .C_ON=1'b0;
    defparam \c0.n18771_bdd_4_lut_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18771_bdd_4_lut_LC_16_8_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18771_bdd_4_lut_LC_16_8_4  (
            .in0(N__49115),
            .in1(N__49149),
            .in2(N__49131),
            .in3(N__49128),
            .lcout(),
            .ltout(\c0.n18774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_16_8_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_16_8_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_16_8_5  (
            .in0(N__47925),
            .in1(N__49116),
            .in2(N__48954),
            .in3(N__48947),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49865),
            .ce(N__48823),
            .sr(_gnd_net_));
    defparam \c0.n18669_bdd_4_lut_LC_16_9_3 .C_ON=1'b0;
    defparam \c0.n18669_bdd_4_lut_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18669_bdd_4_lut_LC_16_9_3 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \c0.n18669_bdd_4_lut_LC_16_9_3  (
            .in0(N__48717),
            .in1(N__48705),
            .in2(N__49914),
            .in3(N__48222),
            .lcout(),
            .ltout(\c0.n18672_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_9_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_9_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_9_4  (
            .in0(N__48180),
            .in1(N__48157),
            .in2(N__48084),
            .in3(N__48075),
            .lcout(\c0.n22_adj_2243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6__2194_LC_16_12_5 .C_ON=1'b0;
    defparam \c0.data_out_7__6__2194_LC_16_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6__2194_LC_16_12_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_7__6__2194_LC_16_12_5  (
            .in0(N__47919),
            .in1(N__47894),
            .in2(N__47791),
            .in3(N__47723),
            .lcout(\c0.data_out_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15718_2_lut_3_lut_LC_16_13_3 .C_ON=1'b0;
    defparam \c0.i15718_2_lut_3_lut_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15718_2_lut_3_lut_LC_16_13_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.i15718_2_lut_3_lut_LC_16_13_3  (
            .in0(N__47633),
            .in1(N__47403),
            .in2(_gnd_net_),
            .in3(N__47143),
            .lcout(data_out_10__7__N_110),
            .ltout(data_out_10__7__N_110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__0__2192_LC_16_13_4 .C_ON=1'b0;
    defparam \c0.data_out_8__0__2192_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__0__2192_LC_16_13_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_out_8__0__2192_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__50949),
            .in2(N__50928),
            .in3(N__50910),
            .lcout(data_out_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49821),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_752_LC_17_2_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_752_LC_17_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_752_LC_17_2_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_752_LC_17_2_3  (
            .in0(N__50757),
            .in1(N__50886),
            .in2(N__50832),
            .in3(N__50822),
            .lcout(\c0.n18_adj_2437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_674_LC_17_4_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_674_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_674_LC_17_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_674_LC_17_4_2  (
            .in0(_gnd_net_),
            .in1(N__50756),
            .in2(_gnd_net_),
            .in3(N__50712),
            .lcout(),
            .ltout(\c0.n6_adj_2409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_675_LC_17_4_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_675_LC_17_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_675_LC_17_4_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_675_LC_17_4_3  (
            .in0(N__50676),
            .in1(N__50625),
            .in2(N__50589),
            .in3(N__50585),
            .lcout(\c0.n17905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i141_LC_17_4_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i141_LC_17_4_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i141_LC_17_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i141_LC_17_4_4  (
            .in0(N__50524),
            .in1(N__49907),
            .in2(_gnd_net_),
            .in3(N__50450),
            .lcout(data_out_frame2_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
