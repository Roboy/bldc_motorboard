-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 21:12:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : inout std_logic;
    PIN_5 : inout std_logic;
    PIN_4 : inout std_logic;
    PIN_3 : out std_logic;
    PIN_24 : out std_logic;
    PIN_23 : out std_logic;
    PIN_22 : out std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : out std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : inout std_logic;
    PIN_11 : inout std_logic;
    PIN_10 : inout std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__51094\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50699\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n4_adj_2271_cascade_\ : std_logic;
signal \c0.n2_adj_2341\ : std_logic;
signal \c0.n2_adj_2341_cascade_\ : std_logic;
signal \c0.n10425\ : std_logic;
signal \c0.n10465\ : std_logic;
signal \n10429_cascade_\ : std_logic;
signal n12965 : std_logic;
signal n242 : std_logic;
signal \n12965_cascade_\ : std_logic;
signal n10429 : std_logic;
signal n8_adj_2541 : std_logic;
signal n18_adj_2539 : std_logic;
signal \n21_adj_2538_cascade_\ : std_logic;
signal n15_adj_2540 : std_logic;
signal \c0.n17263\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n17265\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n17267\ : std_logic;
signal \c0.n17269\ : std_logic;
signal \c0.n17303\ : std_logic;
signal \c0.n17271\ : std_logic;
signal \c0.n17713_cascade_\ : std_logic;
signal \c0.n8_adj_2234\ : std_logic;
signal \c0.n17281\ : std_logic;
signal \c0.n17259\ : std_logic;
signal \c0.n17261\ : std_logic;
signal \c0.n13900\ : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n8_adj_2257\ : std_logic;
signal \c0.n8_adj_2258\ : std_logic;
signal \c0.n39_cascade_\ : std_logic;
signal \c0.n48_adj_2383_cascade_\ : std_logic;
signal \c0.n40\ : std_logic;
signal \c0.n41\ : std_logic;
signal \c0.n43_adj_2384\ : std_logic;
signal \c0.n3_adj_2281\ : std_logic;
signal \c0.n3_adj_2322\ : std_logic;
signal \c0.n3_adj_2311\ : std_logic;
signal \c0.n3_adj_2307\ : std_logic;
signal \c0.n42\ : std_logic;
signal \c0.n3_adj_2299\ : std_logic;
signal \c0.n3_adj_2293\ : std_logic;
signal \c0.n3_adj_2297\ : std_logic;
signal \c0.n3_adj_2326\ : std_logic;
signal \c0.n3_adj_2313\ : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n49_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.n50_adj_2353\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.n17275\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n8_adj_2252\ : std_logic;
signal \c0.n8_adj_2246\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.n17277\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.n17283\ : std_logic;
signal \n17694_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n17279\ : std_logic;
signal \FRAME_MATCHER_state_31_N_1406_0_cascade_\ : std_logic;
signal \n1166_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.n10497_cascade_\ : std_logic;
signal \c0.n17713\ : std_logic;
signal \c0.n17239\ : std_logic;
signal n15 : std_logic;
signal n1437 : std_logic;
signal n8_adj_2498 : std_logic;
signal \c0.n6_adj_2265_cascade_\ : std_logic;
signal \c0.n18907\ : std_logic;
signal \n13_adj_2469_cascade_\ : std_logic;
signal n7 : std_logic;
signal \c0.n3_adj_2301\ : std_logic;
signal \c0.n232_cascade_\ : std_logic;
signal \c0.n6_adj_2364\ : std_logic;
signal n237 : std_logic;
signal \n237_cascade_\ : std_logic;
signal n22_adj_2465 : std_logic;
signal \c0.n3_adj_2309\ : std_logic;
signal \c0.n10353_cascade_\ : std_logic;
signal \c0.n3_adj_2345\ : std_logic;
signal \c0.n3_adj_2343\ : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.n3_adj_2295\ : std_logic;
signal \c0.n3_adj_2291\ : std_logic;
signal \c0.n3_adj_2289\ : std_logic;
signal \c0.n3_adj_2283\ : std_logic;
signal \c0.n3_adj_2279\ : std_logic;
signal \c0.n3_adj_2303\ : std_logic;
signal \PIN_2_c_1\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.n8_adj_2245\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.n17293\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n8_adj_2247\ : std_logic;
signal \c0.n10497\ : std_logic;
signal \c0.n2_adj_2315\ : std_logic;
signal \c0.n8_adj_2273_cascade_\ : std_logic;
signal \c0.n8_adj_2273\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n17273\ : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n17299\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.n46_adj_2356\ : std_logic;
signal \c0.n56\ : std_logic;
signal \c0.n10513_cascade_\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1275\ : std_logic;
signal \c0.n6033_cascade_\ : std_logic;
signal \c0.n2126_cascade_\ : std_logic;
signal \c0.n27\ : std_logic;
signal \c0.n23_cascade_\ : std_logic;
signal \c0.n30_cascade_\ : std_logic;
signal \c0.n50_cascade_\ : std_logic;
signal n13849 : std_logic;
signal \c0.n19_adj_2351\ : std_logic;
signal \c0.n10346\ : std_logic;
signal \c0.n17_cascade_\ : std_logic;
signal \c0.n25_adj_2352\ : std_logic;
signal \c0.n17962_cascade_\ : std_logic;
signal \c0.n4_adj_2226\ : std_logic;
signal \c0.n9575_cascade_\ : std_logic;
signal n12999 : std_logic;
signal \c0.n232\ : std_logic;
signal \n12999_cascade_\ : std_logic;
signal n18 : std_logic;
signal \c0.n9575\ : std_logic;
signal n12966 : std_logic;
signal n15118 : std_logic;
signal \FRAME_MATCHER_i_31__N_1273\ : std_logic;
signal \c0.n16685_cascade_\ : std_logic;
signal \c0.n6_adj_2267\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1270\ : std_logic;
signal \c0.n7528\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.n3_adj_2332\ : std_logic;
signal \c0.n3_adj_2330\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_0\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \c0.n27_adj_2426\ : std_logic;
signal \c0.n16486\ : std_logic;
signal \c0.n115\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n16487\ : std_logic;
signal \c0.n16488\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_4\ : std_logic;
signal \c0.n16489\ : std_logic;
signal \c0.n16490\ : std_logic;
signal \c0.n16491\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_7\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_7\ : std_logic;
signal \c0.n16492\ : std_logic;
signal \c0.n16493\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_8\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_9\ : std_logic;
signal \c0.n16494\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_10\ : std_logic;
signal \c0.n16495\ : std_logic;
signal \c0.n16496\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_12\ : std_logic;
signal \c0.n16497\ : std_logic;
signal \c0.n16498\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_14\ : std_logic;
signal \c0.n16499\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_15\ : std_logic;
signal \c0.n16500\ : std_logic;
signal \c0.n16501\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_16\ : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_16\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_17\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_17\ : std_logic;
signal \c0.n16502\ : std_logic;
signal \c0.n16503\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_19\ : std_logic;
signal \c0.n16504\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_20\ : std_logic;
signal \c0.n16505\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_21\ : std_logic;
signal \c0.n16506\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_22\ : std_logic;
signal \c0.n16507\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_23\ : std_logic;
signal \c0.n16508\ : std_logic;
signal \c0.n16509\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_24\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_25\ : std_logic;
signal \c0.n16510\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_26\ : std_logic;
signal \c0.n16511\ : std_logic;
signal \c0.n16512\ : std_logic;
signal \c0.n16513\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_29\ : std_logic;
signal \c0.n16514\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_30\ : std_logic;
signal \c0.n16515\ : std_logic;
signal \c0.n16516\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_31\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_9\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal \c0.n3_adj_2328\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_6\ : std_logic;
signal \c0.n3_adj_2334\ : std_logic;
signal \control.n18909\ : std_logic;
signal \c0.n8_adj_2254\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.n8_adj_2250\ : std_logic;
signal \c0.n4_adj_2271\ : std_logic;
signal \c0.n8_adj_2249\ : std_logic;
signal \c0.n4_adj_2349\ : std_logic;
signal \c0.n8_adj_2244\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.n30_adj_2355_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n51\ : std_logic;
signal \c0.n10613_cascade_\ : std_logic;
signal \c0.n22_adj_2346\ : std_logic;
signal data_in_frame_5_6 : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.n2126\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal \c0.n2137_adj_2237\ : std_logic;
signal \c0.n2137_adj_2237_cascade_\ : std_logic;
signal data_in_frame_2_0 : std_logic;
signal data_in_frame_2_5 : std_logic;
signal \n16802_cascade_\ : std_logic;
signal \c0.n10569_cascade_\ : std_logic;
signal data_in_frame_0_1 : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \n11058_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_3\ : std_logic;
signal \c0.n1502\ : std_logic;
signal \c0.n1502_cascade_\ : std_logic;
signal \c0.n10522\ : std_logic;
signal \c0.n4_adj_2266\ : std_logic;
signal \c0.n13033_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_30\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_29\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_28\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_19\ : std_logic;
signal \FRAME_MATCHER_i_31\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_31\ : std_logic;
signal \n63_adj_2534_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_18\ : std_logic;
signal \c0.n63_adj_2262_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_5\ : std_logic;
signal \c0.n3_adj_2336\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \c0.n10_adj_2378\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_4\ : std_logic;
signal \c0.n7199\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \c0.n10353\ : std_logic;
signal \c0.n3_adj_2338\ : std_logic;
signal n63 : std_logic;
signal \c0.n63_adj_2262\ : std_logic;
signal n63_adj_2534 : std_logic;
signal \c0.n113\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_6\ : std_logic;
signal \c0.n109\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_11\ : std_logic;
signal \c0.n3_adj_2324\ : std_logic;
signal \c0.n26_adj_2379_cascade_\ : std_logic;
signal \c0.n44_adj_2382\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_12\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_27\ : std_logic;
signal \c0.n13033\ : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_26\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_27\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \c0.n3_adj_2287\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_3\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.n3_adj_2340\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_28\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \c0.n3_adj_2285\ : std_logic;
signal n18043 : std_logic;
signal n18044 : std_logic;
signal \LED_c\ : std_logic;
signal \PIN_3_c_2\ : std_logic;
signal \c0.n4_adj_2225\ : std_logic;
signal tx2_o : std_logic;
signal tx2_enable : std_logic;
signal \c0.n4_adj_2216\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal data_in_frame_2_2 : std_logic;
signal \c0.n18_adj_2417\ : std_logic;
signal data_in_frame_2_1 : std_logic;
signal \c0.n21_adj_2421\ : std_logic;
signal \c0.n24_adj_2418\ : std_logic;
signal \c0.n23_adj_2420_cascade_\ : std_logic;
signal \n16797_cascade_\ : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.rx.n129_cascade_\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal data_in_frame_6_1 : std_logic;
signal data_in_frame_6_7 : std_logic;
signal \c0.n17813\ : std_logic;
signal \c0.n10761\ : std_logic;
signal data_in_frame_0_0 : std_logic;
signal \c0.n10761_cascade_\ : std_logic;
signal \c0.data_in_frame_1_5\ : std_logic;
signal \c0.n17733_cascade_\ : std_logic;
signal data_in_frame_6_0 : std_logic;
signal \c0.n17735\ : std_logic;
signal \c0.data_in_frame_1_6\ : std_logic;
signal \c0.n17733\ : std_logic;
signal \c0.n10569\ : std_logic;
signal data_in_frame_6_3 : std_logic;
signal \c0.n17734_cascade_\ : std_logic;
signal \c0.data_in_frame_1_7\ : std_logic;
signal \c0.n19_adj_2400\ : std_logic;
signal \c0.n18_adj_2398\ : std_logic;
signal \c0.n18000_cascade_\ : std_logic;
signal data_in_frame_5_2 : std_logic;
signal \c0.FRAME_MATCHER_i_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal \c0.rx.n12963\ : std_logic;
signal \n120_cascade_\ : std_logic;
signal data_in_frame_2_3 : std_logic;
signal data_in_frame_0_4 : std_logic;
signal data_in_frame_0_5 : std_logic;
signal data_in_frame_2_6 : std_logic;
signal \c0.n15_adj_2416\ : std_logic;
signal \c0.n2138\ : std_logic;
signal \c0.n22_adj_2419\ : std_logic;
signal data_in_frame_5_7 : std_logic;
signal data_in_frame_2_7 : std_logic;
signal \c0.rx.n17702_cascade_\ : std_logic;
signal \c0.rx.n17702\ : std_logic;
signal \c0.rx.n17704_cascade_\ : std_logic;
signal n11058 : std_logic;
signal n16802 : std_logic;
signal \c0.n18002_cascade_\ : std_logic;
signal \c0.n10498\ : std_logic;
signal \c0.rx.n10988_cascade_\ : std_logic;
signal \c0.rx.n12624_cascade_\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n20_adj_2371_cascade_\ : std_logic;
signal \c0.n10516\ : std_logic;
signal \c0.n10516_cascade_\ : std_logic;
signal \c0.n10367\ : std_logic;
signal data_in_0_5 : std_logic;
signal \c0.n10367_cascade_\ : std_logic;
signal \c0.n15_adj_2389\ : std_logic;
signal data_in_1_4 : std_logic;
signal data_in_0_4 : std_logic;
signal data_in_3_4 : std_logic;
signal \c0.n14_adj_2388\ : std_logic;
signal \c0.n18631\ : std_logic;
signal data_in_1_5 : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.n18_adj_2370\ : std_logic;
signal \c0.n13_adj_2380\ : std_logic;
signal \c0.rx.n10988\ : std_logic;
signal \c0.n18006_cascade_\ : std_logic;
signal \c0.n14_adj_2375\ : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_2_5 : std_logic;
signal rx_data_7 : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \c0.rx.n16532\ : std_logic;
signal \c0.rx.n16533\ : std_logic;
signal \c0.rx.n16534\ : std_logic;
signal \c0.rx.n16535\ : std_logic;
signal \c0.rx.n16536\ : std_logic;
signal \c0.rx.n16537\ : std_logic;
signal \c0.rx.n16538\ : std_logic;
signal \c0.rx.n12819\ : std_logic;
signal \c0.n18225_cascade_\ : std_logic;
signal \c0.rx.n5\ : std_logic;
signal \c0.rx.n57\ : std_logic;
signal \c0.rx.n15905_cascade_\ : std_logic;
signal \c0.rx.n6_cascade_\ : std_logic;
signal \c0.rx.n12\ : std_logic;
signal \c0.rx.n12_cascade_\ : std_logic;
signal \c0.rx.n11082\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \c0.n3_adj_2305\ : std_logic;
signal n1166 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.n3_adj_2317\ : std_logic;
signal n26 : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal n25 : std_logic;
signal n16609 : std_logic;
signal n24 : std_logic;
signal n16610 : std_logic;
signal n23 : std_logic;
signal n16611 : std_logic;
signal n22_adj_2481 : std_logic;
signal n16612 : std_logic;
signal n21 : std_logic;
signal n16613 : std_logic;
signal n20 : std_logic;
signal n16614 : std_logic;
signal n19 : std_logic;
signal n16615 : std_logic;
signal n16616 : std_logic;
signal n18_adj_2480 : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal n17 : std_logic;
signal n16617 : std_logic;
signal n16 : std_logic;
signal n16618 : std_logic;
signal n15_adj_2479 : std_logic;
signal n16619 : std_logic;
signal n14_adj_2478 : std_logic;
signal n16620 : std_logic;
signal n13 : std_logic;
signal n16621 : std_logic;
signal n12 : std_logic;
signal n16622 : std_logic;
signal n11 : std_logic;
signal n16623 : std_logic;
signal n16624 : std_logic;
signal n10_adj_2467 : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal n9 : std_logic;
signal n16625 : std_logic;
signal n8 : std_logic;
signal n16626 : std_logic;
signal n7_adj_2476 : std_logic;
signal n16627 : std_logic;
signal n6 : std_logic;
signal n16628 : std_logic;
signal blink_counter_21 : std_logic;
signal n16629 : std_logic;
signal blink_counter_22 : std_logic;
signal n16630 : std_logic;
signal blink_counter_23 : std_logic;
signal n16631 : std_logic;
signal n16632 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal n16633 : std_logic;
signal blink_counter_25 : std_logic;
signal \control.n11\ : std_logic;
signal \PIN_1_c_0\ : std_logic;
signal \c0.n13808_cascade_\ : std_logic;
signal \c0.n14064_cascade_\ : std_logic;
signal \c0.n4_adj_2203\ : std_logic;
signal \c0.n4_adj_2201\ : std_logic;
signal n17694 : std_logic;
signal \c0.n43\ : std_logic;
signal \c0.n4_adj_2199\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \c0.n18253\ : std_logic;
signal \c0.n16479\ : std_logic;
signal \c0.n18314\ : std_logic;
signal \c0.n16480\ : std_logic;
signal \c0.n18315\ : std_logic;
signal \c0.n16481\ : std_logic;
signal \c0.n16482\ : std_logic;
signal \c0.byte_transmit_counter2_5\ : std_logic;
signal \c0.n18316\ : std_logic;
signal \c0.n16483\ : std_logic;
signal \c0.byte_transmit_counter2_6\ : std_logic;
signal \c0.n18317\ : std_logic;
signal \c0.n16484\ : std_logic;
signal \c0.byte_transmit_counter2_7\ : std_logic;
signal \c0.tx2_transmit_N_1996\ : std_logic;
signal \c0.n16485\ : std_logic;
signal \c0.n18318\ : std_logic;
signal \c0.n18100_cascade_\ : std_logic;
signal \c0.n18103_cascade_\ : std_logic;
signal \c0.n2122\ : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.n16994\ : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal data_in_frame_6_6 : std_logic;
signal data_in_frame_5_1 : std_logic;
signal data_in_frame_6_2 : std_logic;
signal n16797 : std_logic;
signal data_in_frame_5_4 : std_logic;
signal n158 : std_logic;
signal n12600 : std_logic;
signal rx_data_3 : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal \c0.rx.n129\ : std_logic;
signal data_in_frame_5_3 : std_logic;
signal \c0.data_in_frame_1_2\ : std_logic;
signal data_in_frame_5_5 : std_logic;
signal \c0.data_in_frame_1_3\ : std_logic;
signal \c0.n16981_cascade_\ : std_logic;
signal \c0.n20_adj_2397\ : std_logic;
signal \c0.n20_adj_2350\ : std_logic;
signal \c0.n2128\ : std_logic;
signal data_in_frame_6_4 : std_logic;
signal data_in_frame_5_0 : std_logic;
signal \c0.n2128_cascade_\ : std_logic;
signal \c0.n22_adj_2392\ : std_logic;
signal data_in_frame_0_2 : std_logic;
signal data_in_frame_0_3 : std_logic;
signal \c0.n2120\ : std_logic;
signal \c0.n2124\ : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal \c0.n2120_cascade_\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.n19_adj_2415\ : std_logic;
signal \c0.data_in_frame_1_0\ : std_logic;
signal \c0.data_in_frame_1_1\ : std_logic;
signal data_in_frame_0_7 : std_logic;
signal \c0.data_in_frame_1_4\ : std_logic;
signal \c0.n17721_cascade_\ : std_logic;
signal data_in_frame_0_6 : std_logic;
signal \c0.n10_adj_2390\ : std_logic;
signal rx_data_4 : std_logic;
signal n120 : std_logic;
signal data_in_frame_2_4 : std_logic;
signal \c0.rx.n18729_cascade_\ : std_logic;
signal \c0.rx.n18732_cascade_\ : std_logic;
signal \c0.rx.n11\ : std_logic;
signal n12582 : std_logic;
signal n135_adj_2463 : std_logic;
signal \n4_adj_2471_cascade_\ : std_logic;
signal data_in_1_0 : std_logic;
signal \c0.rx.n110\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.rx.r_SM_Main_2_N_2088_2_cascade_\ : std_logic;
signal \c0.rx.n161\ : std_logic;
signal rx_data_0 : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_3_6 : std_logic;
signal \c0.n8_adj_2385\ : std_logic;
signal \c0.n15_adj_2372\ : std_logic;
signal data_in_1_2 : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.rx.r_Bit_Index_0\ : std_logic;
signal n151 : std_logic;
signal \n151_cascade_\ : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.n18008\ : std_logic;
signal \c0.n8_adj_2369_cascade_\ : std_logic;
signal \c0.n10493\ : std_logic;
signal data_in_2_6 : std_logic;
signal data_in_1_6 : std_logic;
signal \c0.rx.n18304\ : std_logic;
signal rx_data_5 : std_logic;
signal data_in_3_5 : std_logic;
signal rx_data_1 : std_logic;
signal data_in_3_0 : std_logic;
signal data_in_2_0 : std_logic;
signal data_in_1_7 : std_logic;
signal \c0.n13693\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2088_2\ : std_logic;
signal \c0.rx.n11041_cascade_\ : std_logic;
signal \c0.rx.r_Bit_Index_2\ : std_logic;
signal \c0.rx.n167\ : std_logic;
signal n12527 : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_3_7 : std_logic;
signal \c0.n6_adj_2368\ : std_logic;
signal data_in_1_3 : std_logic;
signal data_in_0_3 : std_logic;
signal data_in_0_1 : std_logic;
signal \c0.rx.n18196\ : std_logic;
signal \c0.rx.n18194\ : std_logic;
signal \c0.rx.n12552_cascade_\ : std_logic;
signal rx_data_6 : std_logic;
signal \c0.rx.r_Bit_Index_1\ : std_logic;
signal \c0.rx.r_SM_Main_2\ : std_logic;
signal n164_adj_2464 : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.n17990_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.n18024_cascade_\ : std_logic;
signal \c0.rx.n12828\ : std_logic;
signal \c0.rx.n12828_cascade_\ : std_logic;
signal \c0.rx.n18303\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.n15902\ : std_logic;
signal \c0.rx.r_Clock_Count_0\ : std_logic;
signal \c0.rx.n18211\ : std_logic;
signal \c0.rx.r_SM_Main_1\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal \c0.rx.r_SM_Main_0\ : std_logic;
signal \c0.rx.n4\ : std_logic;
signal \c0.tx.n54_cascade_\ : std_logic;
signal \c0.tx.n10\ : std_logic;
signal \c0.tx.n54\ : std_logic;
signal \c0.tx.n47_cascade_\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n16524\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n16525\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n16526\ : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal \c0.tx.n16527\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal \c0.tx.n16528\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal \c0.tx.n16529\ : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal \c0.tx.n16530\ : std_logic;
signal \c0.tx.n16531\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_8\ : std_logic;
signal \c0.tx.n11297\ : std_logic;
signal \control.n8\ : std_logic;
signal \control.PHASES_5_N_2152_1_cascade_\ : std_logic;
signal \control.n10356\ : std_logic;
signal \c0.n18801_cascade_\ : std_logic;
signal \c0.n18804\ : std_logic;
signal \c0.n18843\ : std_logic;
signal \c0.n18846_cascade_\ : std_logic;
signal \c0.n22_adj_2239\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal \c0.n18675_cascade_\ : std_logic;
signal \c0.n18678_cascade_\ : std_logic;
signal \c0.n18741_cascade_\ : std_logic;
signal \c0.n22_adj_2242\ : std_logic;
signal \c0.n18744_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal \n17689_cascade_\ : std_logic;
signal \c0.n18684\ : std_logic;
signal \c0.n18072\ : std_logic;
signal \c0.tx2.n14_cascade_\ : std_logic;
signal \c0.n18284_cascade_\ : std_logic;
signal \c0.n27_adj_2405\ : std_logic;
signal \c0.n29_adj_2408\ : std_logic;
signal \c0.n12704_cascade_\ : std_logic;
signal \c0.n18287\ : std_logic;
signal n612 : std_logic;
signal \c0.n18289_cascade_\ : std_logic;
signal \c0.n18831\ : std_logic;
signal \c0.n18079_cascade_\ : std_logic;
signal \c0.n17725\ : std_logic;
signal \c0.n16863\ : std_logic;
signal \c0.n16982\ : std_logic;
signal \c0.n17722\ : std_logic;
signal \c0.n28_adj_2403\ : std_logic;
signal \c0.n6033\ : std_logic;
signal \c0.n18085_cascade_\ : std_logic;
signal \c0.n4494\ : std_logic;
signal \c0.n28\ : std_logic;
signal \c0.n12704\ : std_logic;
signal \c0.n18082\ : std_logic;
signal \c0.n18270\ : std_logic;
signal \c0.n6035\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \c0.tx2.n16539\ : std_logic;
signal \c0.tx2.n16540\ : std_logic;
signal \c0.tx2.n16541\ : std_logic;
signal \c0.tx2.n16542\ : std_logic;
signal \c0.tx2.n16543\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \c0.tx2.n16544\ : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \c0.tx2.n16545\ : std_logic;
signal \c0.tx2.n16546\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \c0.tx2.r_Clock_Count_8\ : std_logic;
signal \c0.tx2.n11312\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \c0.n16517\ : std_logic;
signal \c0.n16518\ : std_logic;
signal \c0.n16519\ : std_logic;
signal \c0.n16520\ : std_logic;
signal \c0.n16521\ : std_logic;
signal \c0.n16522\ : std_logic;
signal \c0.n16523\ : std_logic;
signal \c0.n18254\ : std_logic;
signal \c0.n4_adj_2231\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.n73\ : std_logic;
signal \c0.n44\ : std_logic;
signal tx_enable : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal data_in_1_1 : std_logic;
signal \n3_adj_2525_cascade_\ : std_logic;
signal tx_o : std_logic;
signal \c0.tx.n17697\ : std_logic;
signal data_out_1_7 : std_logic;
signal \c0.tx.n11030_cascade_\ : std_logic;
signal \c0.tx.n18041\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_2062\ : std_logic;
signal n18750 : std_logic;
signal \n10_adj_2532_cascade_\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.tx.n17984\ : std_logic;
signal \n10_adj_2537_cascade_\ : std_logic;
signal \n10_adj_2535_cascade_\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \c0.n18188\ : std_logic;
signal n5155 : std_logic;
signal \c0.n18354\ : std_logic;
signal n18756 : std_logic;
signal \c0.data_out_3_6\ : std_logic;
signal data_out_3_7 : std_logic;
signal data_out_2_7 : std_logic;
signal \c0.n2_adj_2229\ : std_logic;
signal \n2837_cascade_\ : std_logic;
signal data_out_0_5 : std_logic;
signal \control.n12_cascade_\ : std_logic;
signal \control.n10\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \control.n9_adj_2459\ : std_logic;
signal \control.n16647\ : std_logic;
signal \control.pwm_delay_2\ : std_logic;
signal \control.n16648\ : std_logic;
signal \control.pwm_delay_3\ : std_logic;
signal \control.n16649\ : std_logic;
signal \control.pwm_delay_4\ : std_logic;
signal \control.n16650\ : std_logic;
signal \control.pwm_delay_5\ : std_logic;
signal \control.n16651\ : std_logic;
signal \control.pwm_delay_6\ : std_logic;
signal \control.n16652\ : std_logic;
signal \control.pwm_delay_7\ : std_logic;
signal \control.n16653\ : std_logic;
signal \control.n16654\ : std_logic;
signal \control.pwm_delay_8\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \control.n16655\ : std_logic;
signal \c0.n18888_cascade_\ : std_logic;
signal \c0.n18789_cascade_\ : std_logic;
signal \c0.n18792_cascade_\ : std_logic;
signal \c0.n22_adj_2270\ : std_logic;
signal \c0.n18885\ : std_logic;
signal \c0.n10861_cascade_\ : std_logic;
signal \c0.n18798\ : std_logic;
signal \c0.n10893_cascade_\ : std_logic;
signal data_out_frame2_17_1 : std_logic;
signal \c0.n5_adj_2435_cascade_\ : std_logic;
signal \c0.n6_adj_2223\ : std_logic;
signal \c0.n18687_cascade_\ : std_logic;
signal \c0.n18690\ : std_logic;
signal \c0.n5_adj_2197\ : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n6_adj_2354\ : std_logic;
signal \c0.n18855\ : std_logic;
signal tx2_active : std_logic;
signal \c0.n14064\ : std_logic;
signal \c0.n12359_cascade_\ : std_logic;
signal \c0.n6_adj_2443_cascade_\ : std_logic;
signal \c0.n10513\ : std_logic;
signal \c0.FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n10958\ : std_logic;
signal \c0.r_SM_Main_2_N_2034_0_adj_2213\ : std_logic;
signal n6707 : std_logic;
signal \c0.tx2.n12769\ : std_logic;
signal \r_SM_Main_2_N_2031_1\ : std_logic;
signal \r_SM_Main_2_N_2031_1_cascade_\ : std_logic;
signal \n18014_cascade_\ : std_logic;
signal \c0.n18362\ : std_logic;
signal \c0.n12359\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1272\ : std_logic;
signal \c0.n4_adj_2204\ : std_logic;
signal \c0.tx2.n13800\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal n3 : std_logic;
signal \c0.tx2.n18164\ : std_logic;
signal \c0.tx2.n18163\ : std_logic;
signal \c0.tx2.n18062\ : std_logic;
signal \c0.tx2.n18717_cascade_\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_2062\ : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal \c0.tx2.n10\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal \c0.tx2.n10_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.n12775\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.n18061\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal n11096 : std_logic;
signal \c0.n18260_cascade_\ : std_logic;
signal \c0.n130\ : std_logic;
signal \c0.n3465\ : std_logic;
signal \c0.n4806\ : std_logic;
signal byte_transmit_counter_6 : std_logic;
signal \tx_transmit_N_1947_6\ : std_logic;
signal \tx_transmit_N_1947_4\ : std_logic;
signal \c0.n4_cascade_\ : std_logic;
signal \n5341_cascade_\ : std_logic;
signal \tx_transmit_N_1947_7\ : std_logic;
signal byte_transmit_counter_7 : std_logic;
signal \c0.tx_transmit_N_1947_5\ : std_logic;
signal n10973 : std_logic;
signal n5341 : std_logic;
signal \c0.byte_transmit_counter_5\ : std_logic;
signal \c0.n17998\ : std_logic;
signal \c0.tx.n17938\ : std_logic;
signal n10_adj_2536 : std_logic;
signal \n5440_cascade_\ : std_logic;
signal n18016 : std_logic;
signal \n18016_cascade_\ : std_logic;
signal \c0.n8_adj_2207\ : std_logic;
signal \c0.tx.n13802\ : std_logic;
signal \c0.tx.n13802_cascade_\ : std_logic;
signal \c0.tx.n6796_cascade_\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal \c0.tx.n18167\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \c0.tx.n18711\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.tx.n18040\ : std_logic;
signal \c0.n8_adj_2205\ : std_logic;
signal \c0.tx.r_SM_Main_2\ : std_logic;
signal \c0.tx.r_SM_Main_0\ : std_logic;
signal \c0.tx.r_SM_Main_1\ : std_logic;
signal \c0.tx.r_SM_Main_2_N_2031_1\ : std_logic;
signal n18012 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.tx.n18166\ : std_logic;
signal \c0.n5_adj_2241\ : std_logic;
signal \c0.n18753\ : std_logic;
signal \c0.n2\ : std_logic;
signal \c0.n18189\ : std_logic;
signal \n18876_cascade_\ : std_logic;
signal n10_adj_2531 : std_logic;
signal \c0.n5_adj_2196_cascade_\ : std_logic;
signal \c0.n18873\ : std_logic;
signal \n5_cascade_\ : std_logic;
signal \c0.n8_adj_2209\ : std_logic;
signal n10_adj_2533 : std_logic;
signal \n10_adj_2528_cascade_\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal data_out_3_5 : std_logic;
signal data_out_1_6 : std_logic;
signal \c0.data_out_0_6\ : std_logic;
signal \c0.n1_adj_2272\ : std_logic;
signal data_out_2_5 : std_logic;
signal \c0.n18335\ : std_logic;
signal \c0.data_out_2_3\ : std_logic;
signal \c0.n19_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_1\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.n18266\ : std_logic;
signal \c0.n18360\ : std_logic;
signal \c0.n18256\ : std_logic;
signal \c0.n14_adj_2359_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_0\ : std_logic;
signal \c0.n15_adj_2429\ : std_logic;
signal \c0.n17847\ : std_logic;
signal \c0.n10867_cascade_\ : std_logic;
signal \c0.n17739_cascade_\ : std_logic;
signal data_out_frame2_17_0 : std_logic;
signal \c0.n18840\ : std_logic;
signal \c0.n18795\ : std_logic;
signal data_out_frame2_18_7 : std_logic;
signal data_out_frame2_5_1 : std_logic;
signal \c0.n18837\ : std_logic;
signal data_out_frame2_18_1 : std_logic;
signal data_out_frame2_17_7 : std_logic;
signal \c0.n17727\ : std_logic;
signal data_out_frame2_7_1 : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \c0.n16634\ : std_logic;
signal \c0.n16635\ : std_logic;
signal \c0.n16636\ : std_logic;
signal \c0.n16637\ : std_logic;
signal \c0.n16638\ : std_logic;
signal \c0.n16639\ : std_logic;
signal \c0.n16640\ : std_logic;
signal \c0.n16641\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \c0.n16642\ : std_logic;
signal \c0.n16643\ : std_logic;
signal \c0.n16644\ : std_logic;
signal \c0.n16645\ : std_logic;
signal \c0.n16646\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal n26_adj_2466 : std_logic;
signal \c0.n18019\ : std_logic;
signal n129 : std_logic;
signal \c0.r_SM_Main_2_N_2034_0\ : std_logic;
signal \n129_cascade_\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal \c0.n1707\ : std_logic;
signal \c0.delay_counter_11\ : std_logic;
signal \c0.delay_counter_12\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.n24\ : std_logic;
signal n12227 : std_logic;
signal \n574_cascade_\ : std_logic;
signal \c0.n98\ : std_logic;
signal \c0.n18230\ : std_logic;
signal \n17978_cascade_\ : std_logic;
signal \UART_TRANSMITTER_state_7_N_1223_1\ : std_logic;
signal n18202 : std_logic;
signal n574 : std_logic;
signal n4 : std_logic;
signal n22_adj_2522 : std_logic;
signal \c0.n18226\ : std_logic;
signal n21_adj_2524 : std_logic;
signal n6_adj_2470 : std_logic;
signal n18368 : std_logic;
signal \c0.n18861_cascade_\ : std_logic;
signal \c0.n18377\ : std_logic;
signal \n18864_cascade_\ : std_logic;
signal \n10_adj_2529_cascade_\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal n10_adj_2499 : std_logic;
signal \c0.n10550_cascade_\ : std_logic;
signal \c0.n10524\ : std_logic;
signal \c0.n10550\ : std_logic;
signal \c0.n10746\ : std_logic;
signal \c0.n6_adj_2361\ : std_logic;
signal \c0.n10746_cascade_\ : std_logic;
signal \n17758_cascade_\ : std_logic;
signal \c0.n10734\ : std_logic;
signal \c0.n8_adj_2232\ : std_logic;
signal n10_adj_2461 : std_logic;
signal data_out_8_7 : std_logic;
signal \c0.n17742_cascade_\ : std_logic;
signal \c0.n17742\ : std_logic;
signal \c0.n10558\ : std_logic;
signal \c0.data_out_9_5\ : std_logic;
signal \c0.n6_adj_2365_cascade_\ : std_logic;
signal \c0.n5_adj_2220\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n18265\ : std_logic;
signal n9667 : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \c0.n1_cascade_\ : std_logic;
signal n22 : std_logic;
signal \c0.n18849\ : std_logic;
signal \n18852_cascade_\ : std_logic;
signal n10 : std_logic;
signal \c0.n18264\ : std_logic;
signal \c0.n8\ : std_logic;
signal n10_adj_2527 : std_logic;
signal \c0.n18322\ : std_logic;
signal data_out_0_1 : std_logic;
signal \n11017_cascade_\ : std_logic;
signal data_out_0_0 : std_logic;
signal data_out_3_4 : std_logic;
signal \control.PHASES_5_N_2152_1\ : std_logic;
signal \control.pwm_delay_9\ : std_logic;
signal \control.n18\ : std_logic;
signal \control.n17926\ : std_logic;
signal \control.PHASES_5__N_2160_cascade_\ : std_logic;
signal \control.n5\ : std_logic;
signal \control.n17950\ : std_logic;
signal \control.n9\ : std_logic;
signal \c0.n18639_cascade_\ : std_logic;
signal \c0.n10700_cascade_\ : std_logic;
signal \c0.n21\ : std_logic;
signal \c0.n17804\ : std_logic;
signal \c0.n17874\ : std_logic;
signal \c0.n17908\ : std_logic;
signal \c0.n18_adj_2423\ : std_logic;
signal \c0.n17908_cascade_\ : std_logic;
signal \c0.n28_adj_2425\ : std_logic;
signal \c0.n30_adj_2424_cascade_\ : std_logic;
signal \c0.n29_adj_2427\ : std_logic;
signal data_out_frame2_17_5 : std_logic;
signal data_out_frame2_12_1 : std_logic;
signal \c0.n10829_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_1\ : std_logic;
signal \c0.n14161\ : std_logic;
signal \c0.FRAME_MATCHER_state_2\ : std_logic;
signal \c0.n50\ : std_logic;
signal \n11114_cascade_\ : std_logic;
signal data_out_frame2_18_0 : std_logic;
signal data_out_frame2_6_7 : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.delay_counter_13\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.n18810\ : std_logic;
signal \c0.tx_transmit_N_1947_0\ : std_logic;
signal \c0.tx_transmit_N_1947_1\ : std_logic;
signal \c0.tx_transmit_N_1947_2\ : std_logic;
signal \c0.n155\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.n22\ : std_logic;
signal n25_adj_2468 : std_logic;
signal \c0.n18807\ : std_logic;
signal \c0.n5_adj_2436\ : std_logic;
signal \r_Bit_Index_0_adj_2519\ : std_logic;
signal \r_Bit_Index_1_adj_2518\ : std_logic;
signal \tx_transmit_N_1947_3\ : std_logic;
signal \c0.n85\ : std_logic;
signal \c0.n14068\ : std_logic;
signal \c0.n18259\ : std_logic;
signal n18014 : std_logic;
signal n4_adj_2472 : std_logic;
signal n11545 : std_logic;
signal \r_Bit_Index_2_adj_2517\ : std_logic;
signal \c0.n17715\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \c0.n18\ : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_3_3 : std_logic;
signal rx_data_ready : std_logic;
signal data_in_2_3 : std_logic;
signal \c0.n18365\ : std_logic;
signal data_out_frame2_18_5 : std_logic;
signal n1 : std_logic;
signal n24_adj_2523 : std_logic;
signal n18_adj_2526 : std_logic;
signal \c0.n17761_cascade_\ : std_logic;
signal n9_adj_2477 : std_logic;
signal \c0.n17761\ : std_logic;
signal \c0.n18747\ : std_logic;
signal \c0.n17807_cascade_\ : std_logic;
signal data_out_9_2 : std_logic;
signal \c0.n6_adj_2318_cascade_\ : std_logic;
signal \c0.data_out_9_0\ : std_logic;
signal \c0.data_out_9_6\ : std_logic;
signal \c0.n6_adj_2367\ : std_logic;
signal \c0.n17850\ : std_logic;
signal \c0.n10749\ : std_logic;
signal \c0.data_out_9__2__N_367_cascade_\ : std_logic;
signal \c0.n15_adj_2319_cascade_\ : std_logic;
signal \c0.n14_adj_2320\ : std_logic;
signal \c0.data_out_10_2\ : std_logic;
signal \c0.n17826\ : std_logic;
signal \c0.data_out_9_7\ : std_logic;
signal \c0.n17774\ : std_logic;
signal \c0.n17774_cascade_\ : std_logic;
signal \c0.data_out_10_3\ : std_logic;
signal \c0.data_out_10_5\ : std_logic;
signal \c0.n6_adj_2314\ : std_logic;
signal \c0.n17883\ : std_logic;
signal \c0.n10801_cascade_\ : std_logic;
signal \c0.data_out_10_0\ : std_logic;
signal \c0.n17768\ : std_logic;
signal \c0.n10_adj_2366_cascade_\ : std_logic;
signal \c0.data_out_10_1\ : std_logic;
signal \c0.data_out_6_1\ : std_logic;
signal \c0.n17819\ : std_logic;
signal \c0.n6_adj_2277\ : std_logic;
signal \c0.data_out_9_4\ : std_logic;
signal \c0.n8_adj_2211_cascade_\ : std_logic;
signal \c0.n18222_cascade_\ : std_logic;
signal \c0.n18693_cascade_\ : std_logic;
signal n18696 : std_logic;
signal \c0.data_out_6_2\ : std_logic;
signal \c0.n5_adj_2347\ : std_logic;
signal byte_transmit_counter_1 : std_logic;
signal \c0.n18191\ : std_logic;
signal \c0.n18867_cascade_\ : std_logic;
signal byte_transmit_counter_2 : std_logic;
signal n10_adj_2505 : std_logic;
signal \n18870_cascade_\ : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal n10_adj_2530 : std_logic;
signal \c0.n5_adj_2214\ : std_logic;
signal \c0.data_out_1_4\ : std_logic;
signal \c0.n18190\ : std_logic;
signal \c0.n2_adj_2348\ : std_logic;
signal \c0.n18334\ : std_logic;
signal \c0.data_out_7_4\ : std_logic;
signal data_out_3_2 : std_logic;
signal \c0.data_out_1_2\ : std_logic;
signal \c0.n18223\ : std_logic;
signal data_out_2_2 : std_logic;
signal \PIN_24_c_3\ : std_logic;
signal \control.n6\ : std_logic;
signal \control.n17251\ : std_logic;
signal \PIN_23_c_4\ : std_logic;
signal \control.n6_adj_2460\ : std_logic;
signal \control.n10490\ : std_logic;
signal hall3 : std_logic;
signal hall2 : std_logic;
signal hall1 : std_logic;
signal \control.PHASES_5__N_2160\ : std_logic;
signal \control.PHASES_5_N_2130_5\ : std_logic;
signal \c0.n17748\ : std_logic;
signal data_out_frame2_15_1 : std_logic;
signal \c0.n10829\ : std_logic;
signal \c0.n10890_cascade_\ : std_logic;
signal \c0.n17_adj_2449\ : std_logic;
signal \c0.n16_adj_2448_cascade_\ : std_logic;
signal \c0.n17911\ : std_logic;
signal \c0.n15_adj_2445\ : std_logic;
signal \c0.n14_adj_2444_cascade_\ : std_logic;
signal data_out_frame2_16_1 : std_logic;
signal \c0.data_out_frame2_20_5\ : std_logic;
signal \c0.n16_adj_2358\ : std_logic;
signal \c0.n10720_cascade_\ : std_logic;
signal data_out_frame2_10_2 : std_logic;
signal \c0.n10819\ : std_logic;
signal \c0.n17886\ : std_logic;
signal \c0.n20_adj_2442\ : std_logic;
signal \c0.n16_cascade_\ : std_logic;
signal \c0.n17795\ : std_logic;
signal \c0.data_out_frame2_19_5\ : std_logic;
signal \c0.n10839\ : std_logic;
signal \c0.n10890\ : std_logic;
signal data_out_frame2_10_5 : std_logic;
signal \c0.n10816\ : std_logic;
signal \c0.n12_adj_2446_cascade_\ : std_logic;
signal data_out_frame2_6_4 : std_logic;
signal \c0.n10864\ : std_logic;
signal \c0.n10_adj_2440\ : std_logic;
signal \c0.n6_adj_2357\ : std_logic;
signal \c0.n18879_cascade_\ : std_logic;
signal \c0.n10852\ : std_logic;
signal \c0.n10867\ : std_logic;
signal data_out_frame2_8_5 : std_logic;
signal \c0.n14_adj_2447\ : std_logic;
signal \c0.data_out_frame2_19_4\ : std_logic;
signal data_out_frame2_15_3 : std_logic;
signal \c0.n6_adj_2422_cascade_\ : std_logic;
signal data_out_frame2_18_4 : std_logic;
signal \c0.n10870_cascade_\ : std_logic;
signal \c0.n27_adj_2428\ : std_logic;
signal \c0.n5_adj_2274\ : std_logic;
signal data_out_8_2 : std_logic;
signal \c0.n11056\ : std_logic;
signal \c0.n18199_cascade_\ : std_logic;
signal \c0.n17832\ : std_logic;
signal \c0.n18242_cascade_\ : std_logic;
signal \c0.data_out_6_6\ : std_logic;
signal \c0.n5\ : std_logic;
signal \c0.n18247\ : std_logic;
signal \c0.n18238_cascade_\ : std_logic;
signal \c0.data_out_6_4\ : std_logic;
signal \c0.n6_adj_2276\ : std_logic;
signal \c0.data_out_6_7\ : std_logic;
signal \c0.data_out_6_5\ : std_logic;
signal data_out_8_4 : std_logic;
signal \c0.n17745\ : std_logic;
signal \c0.n10542\ : std_logic;
signal \c0.n17745_cascade_\ : std_logic;
signal \c0.data_out_10_7\ : std_logic;
signal data_out_8_3 : std_logic;
signal \c0.n8_adj_2219\ : std_logic;
signal data_out_0_3 : std_logic;
signal \c0.n18376\ : std_logic;
signal data_out_10_6 : std_logic;
signal \c0.data_out_7_2\ : std_logic;
signal \c0.data_out_9_1\ : std_logic;
signal \c0.n17730\ : std_logic;
signal \c0.n17835\ : std_logic;
signal \c0.n17844\ : std_logic;
signal \c0.n17730_cascade_\ : std_logic;
signal n17758 : std_logic;
signal \c0.n14_adj_2363_cascade_\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.data_out_9_3\ : std_logic;
signal \c0.n17816_cascade_\ : std_logic;
signal \c0.n17877\ : std_logic;
signal \c0.n12\ : std_logic;
signal \c0.n17786\ : std_logic;
signal \c0.n18184\ : std_logic;
signal \c0.data_out_7_1\ : std_logic;
signal \c0.n10537\ : std_logic;
signal data_out_6_0 : std_logic;
signal \c0.n10680\ : std_logic;
signal \c0.n17816\ : std_logic;
signal \c0.n10680_cascade_\ : std_logic;
signal \c0.data_out_5_5\ : std_logic;
signal data_out_8_6 : std_logic;
signal data_out_8_5 : std_logic;
signal \c0.n17771\ : std_logic;
signal data_out_5_1 : std_logic;
signal \c0.data_out_5_4\ : std_logic;
signal data_out_frame2_13_2 : std_logic;
signal data_out_frame2_16_0 : std_logic;
signal data_out_frame2_8_6 : std_logic;
signal \c0.n18759_cascade_\ : std_logic;
signal data_out_frame2_6_0 : std_logic;
signal \c0.n10920\ : std_logic;
signal \c0.n17783_cascade_\ : std_logic;
signal \c0.n10849\ : std_logic;
signal \c0.n17859\ : std_logic;
signal \c0.n15_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_0\ : std_logic;
signal \c0.n10688\ : std_logic;
signal \c0.n10813_cascade_\ : std_logic;
signal \c0.n10577\ : std_logic;
signal \c0.n17783\ : std_logic;
signal \c0.n15_adj_2414_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_1\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.n32_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_7\ : std_logic;
signal \c0.data_out_frame2_0_7\ : std_logic;
signal \c0.n17777\ : std_logic;
signal \c0.n6_adj_2430\ : std_logic;
signal \c0.n17777_cascade_\ : std_logic;
signal data_out_frame2_5_5 : std_logic;
signal \c0.n10617_cascade_\ : std_logic;
signal \c0.n17765\ : std_logic;
signal \c0.data_out_frame2_0_4\ : std_logic;
signal \c0.n18681\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal n16547 : std_logic;
signal n16548 : std_logic;
signal n16549 : std_logic;
signal n16550 : std_logic;
signal n16551 : std_logic;
signal n16552 : std_logic;
signal n16553 : std_logic;
signal n16554 : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal n16555 : std_logic;
signal n16556 : std_logic;
signal n16557 : std_logic;
signal n16558 : std_logic;
signal n16559 : std_logic;
signal n16560 : std_logic;
signal n16561 : std_logic;
signal n16562 : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal n16563 : std_logic;
signal n16564 : std_logic;
signal n16565 : std_logic;
signal n16566 : std_logic;
signal n16567 : std_logic;
signal n16568 : std_logic;
signal n16569 : std_logic;
signal n16570 : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal n16571 : std_logic;
signal n16572 : std_logic;
signal n16573 : std_logic;
signal n16574 : std_logic;
signal n16575 : std_logic;
signal n16576 : std_logic;
signal n16577 : std_logic;
signal rand_data_0 : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal rand_data_1 : std_logic;
signal n16578 : std_logic;
signal rand_data_2 : std_logic;
signal rand_setpoint_2 : std_logic;
signal n16579 : std_logic;
signal rand_data_3 : std_logic;
signal rand_setpoint_3 : std_logic;
signal n16580 : std_logic;
signal rand_data_4 : std_logic;
signal rand_setpoint_4 : std_logic;
signal n16581 : std_logic;
signal rand_setpoint_5 : std_logic;
signal n16582 : std_logic;
signal rand_setpoint_6 : std_logic;
signal n16583 : std_logic;
signal rand_setpoint_7 : std_logic;
signal n16584 : std_logic;
signal n16585 : std_logic;
signal rand_data_8 : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal rand_data_9 : std_logic;
signal rand_setpoint_9 : std_logic;
signal n16586 : std_logic;
signal rand_data_10 : std_logic;
signal rand_setpoint_10 : std_logic;
signal n16587 : std_logic;
signal n16588 : std_logic;
signal rand_setpoint_12 : std_logic;
signal n16589 : std_logic;
signal rand_data_13 : std_logic;
signal n16590 : std_logic;
signal rand_data_14 : std_logic;
signal n16591 : std_logic;
signal rand_data_15 : std_logic;
signal rand_setpoint_15 : std_logic;
signal n16592 : std_logic;
signal n16593 : std_logic;
signal rand_data_16 : std_logic;
signal rand_setpoint_16 : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal rand_data_17 : std_logic;
signal rand_setpoint_17 : std_logic;
signal n16594 : std_logic;
signal rand_setpoint_18 : std_logic;
signal n16595 : std_logic;
signal rand_data_19 : std_logic;
signal rand_setpoint_19 : std_logic;
signal n16596 : std_logic;
signal rand_data_20 : std_logic;
signal rand_setpoint_20 : std_logic;
signal n16597 : std_logic;
signal rand_data_21 : std_logic;
signal rand_setpoint_21 : std_logic;
signal n16598 : std_logic;
signal rand_data_22 : std_logic;
signal rand_setpoint_22 : std_logic;
signal n16599 : std_logic;
signal rand_data_23 : std_logic;
signal rand_setpoint_23 : std_logic;
signal n16600 : std_logic;
signal n16601 : std_logic;
signal rand_data_24 : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal rand_data_25 : std_logic;
signal rand_setpoint_25 : std_logic;
signal n16602 : std_logic;
signal rand_data_26 : std_logic;
signal n16603 : std_logic;
signal n16604 : std_logic;
signal rand_setpoint_28 : std_logic;
signal n16605 : std_logic;
signal rand_data_29 : std_logic;
signal rand_setpoint_29 : std_logic;
signal n16606 : std_logic;
signal rand_data_30 : std_logic;
signal n16607 : std_logic;
signal rand_data_31 : std_logic;
signal n16608 : std_logic;
signal rand_setpoint_13 : std_logic;
signal \c0.n18234\ : std_logic;
signal rand_setpoint_1 : std_logic;
signal \c0.data_out_8_1\ : std_logic;
signal \c0.data_out_7_5\ : std_logic;
signal \c0.data_out_7_7\ : std_logic;
signal \c0.n10533\ : std_logic;
signal rand_setpoint_26 : std_logic;
signal \c0.data_out_5_2\ : std_logic;
signal rand_setpoint_30 : std_logic;
signal rand_setpoint_27 : std_logic;
signal \c0.data_out_5_3\ : std_logic;
signal \c0.n17718\ : std_logic;
signal \c0.n17829\ : std_logic;
signal \c0.data_out_10_4\ : std_logic;
signal n2837 : std_logic;
signal data_out_3_0 : std_logic;
signal \c0.n2_adj_2221\ : std_logic;
signal data_out_2_0 : std_logic;
signal \c0.n5_adj_2433\ : std_logic;
signal data_out_frame2_14_7 : std_logic;
signal \c0.n17899\ : std_logic;
signal \c0.n17899_cascade_\ : std_logic;
signal \c0.n34\ : std_logic;
signal \c0.n17736\ : std_logic;
signal \c0.n17736_cascade_\ : std_logic;
signal \c0.n18813\ : std_logic;
signal \c0.n18816\ : std_logic;
signal data_out_frame2_9_6 : std_logic;
signal \c0.n10725\ : std_logic;
signal data_out_frame2_7_0 : std_logic;
signal \c0.n10700\ : std_logic;
signal \c0.n16_adj_2412\ : std_logic;
signal \c0.n17_adj_2413_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_1\ : std_logic;
signal \c0.n10782\ : std_logic;
signal data_out_frame2_14_1 : std_logic;
signal \c0.n17862\ : std_logic;
signal \c0.n17862_cascade_\ : std_logic;
signal \c0.n17841\ : std_logic;
signal \c0.n12_adj_2410_cascade_\ : std_logic;
signal data_out_frame2_16_7 : std_logic;
signal data_out_frame2_15_7 : std_logic;
signal \c0.n17889\ : std_logic;
signal rand_data_18 : std_logic;
signal data_out_frame2_6_2 : std_logic;
signal \c0.n18645\ : std_logic;
signal \c0.n18_adj_2441\ : std_logic;
signal data_out_frame2_8_3 : std_logic;
signal data_out_frame2_10_1 : std_logic;
signal \c0.n17838\ : std_logic;
signal \c0.n17792\ : std_logic;
signal \c0.n33\ : std_logic;
signal data_out_frame2_6_6 : std_logic;
signal data_out_frame2_10_3 : std_logic;
signal \c0.n18663\ : std_logic;
signal data_out_frame2_5_0 : std_logic;
signal \c0.n10911\ : std_logic;
signal data_out_frame2_11_6 : std_logic;
signal rand_data_6 : std_logic;
signal data_out_frame2_9_4 : std_logic;
signal data_out_frame2_7_7 : std_logic;
signal data_out_frame2_9_7 : std_logic;
signal \c0.n10617\ : std_logic;
signal \c0.n14_adj_2362\ : std_logic;
signal data_out_frame2_12_2 : std_logic;
signal data_out_frame2_10_4 : std_logic;
signal \c0.n17880\ : std_logic;
signal \c0.n17789\ : std_logic;
signal data_out_frame2_5_6 : std_logic;
signal \c0.n5_adj_2439\ : std_logic;
signal \c0.data_out_frame2_0_6\ : std_logic;
signal data_out_frame2_15_6 : std_logic;
signal data_out_frame2_13_1 : std_logic;
signal data_out_frame2_8_7 : std_logic;
signal \c0.data_out_frame2_0_0\ : std_logic;
signal \c0.n10_adj_2431\ : std_logic;
signal data_out_frame2_5_2 : std_logic;
signal \c0.n17865\ : std_logic;
signal rand_data_28 : std_logic;
signal rand_data_11 : std_logic;
signal data_out_frame2_13_7 : std_logic;
signal \c0.n10_adj_2411\ : std_logic;
signal \c0.n18705\ : std_logic;
signal data_out_frame2_13_6 : std_logic;
signal rand_data_27 : std_logic;
signal rand_data_7 : std_logic;
signal data_out_frame2_13_3 : std_logic;
signal \c0.n18657\ : std_logic;
signal data_out_frame2_18_3 : std_logic;
signal \c0.data_out_frame2_19_3\ : std_logic;
signal data_out_frame2_17_3 : std_logic;
signal \c0.n18651_cascade_\ : std_logic;
signal data_out_frame2_16_3 : std_logic;
signal \c0.data_out_frame2_20_3\ : std_logic;
signal \c0.n18654_cascade_\ : std_logic;
signal \c0.n18666\ : std_logic;
signal \c0.n18660\ : std_logic;
signal \c0.n18371\ : std_logic;
signal \c0.n18735_cascade_\ : std_logic;
signal \c0.n6_adj_2360\ : std_logic;
signal \c0.n22_adj_2259\ : std_logic;
signal \c0.n18738_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal data_out_frame2_18_6 : std_logic;
signal \c0.n18708\ : std_logic;
signal \c0.n18762\ : std_logic;
signal \c0.n18308\ : std_logic;
signal \c0.n18777_cascade_\ : std_logic;
signal \c0.n6_adj_2218\ : std_logic;
signal \c0.n18699\ : std_logic;
signal data_out_frame2_17_6 : std_logic;
signal data_out_frame2_16_6 : std_logic;
signal \c0.n18702_cascade_\ : std_logic;
signal \c0.n18780\ : std_logic;
signal \c0.n22_adj_2240_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal \c0.n18783_cascade_\ : std_logic;
signal data_out_frame2_13_4 : std_logic;
signal \c0.data_out_7__2__N_447\ : std_logic;
signal \c0.n18311\ : std_logic;
signal rand_setpoint_11 : std_logic;
signal byte_transmit_counter_0 : std_logic;
signal \c0.data_out_6_3\ : std_logic;
signal \c0.n5_adj_2217\ : std_logic;
signal \c0.n18201\ : std_logic;
signal \c0.data_out_7_3\ : std_logic;
signal rand_setpoint_24 : std_logic;
signal \c0.data_out_6__1__N_537\ : std_logic;
signal rand_setpoint_31 : std_logic;
signal \c0.data_out_7__3__N_441\ : std_logic;
signal \c0.n11277\ : std_logic;
signal \c0.data_out_1_1\ : std_logic;
signal n11017 : std_logic;
signal \c0.n18250\ : std_logic;
signal rand_setpoint_8 : std_logic;
signal \c0.data_out_7_0\ : std_logic;
signal \c0.n18648\ : std_logic;
signal \c0.n18642\ : std_logic;
signal \c0.n18221\ : std_logic;
signal \c0.n18765_cascade_\ : std_logic;
signal \c0.n6_adj_2227\ : std_logic;
signal \c0.n18768_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal data_out_frame2_18_2 : std_logic;
signal \c0.data_out_frame2_19_2\ : std_logic;
signal data_out_frame2_17_2 : std_logic;
signal \c0.n18633_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_2\ : std_logic;
signal \c0.n18636_cascade_\ : std_logic;
signal \c0.n22_adj_2268\ : std_logic;
signal \c0.n17892\ : std_logic;
signal data_out_frame2_9_1 : std_logic;
signal \c0.n10893\ : std_logic;
signal \c0.n20_adj_2438_cascade_\ : std_logic;
signal \c0.n17755\ : std_logic;
signal \c0.data_out_frame2_19_6\ : std_logic;
signal data_out_frame2_5_3 : std_logic;
signal data_out_frame2_12_3 : std_logic;
signal \c0.n10905\ : std_logic;
signal \c0.n10905_cascade_\ : std_logic;
signal \c0.n16_adj_2391\ : std_logic;
signal data_out_frame2_8_2 : std_logic;
signal data_out_frame2_14_6 : std_logic;
signal data_out_frame2_11_7 : std_logic;
signal data_out_frame2_14_5 : std_logic;
signal data_out_frame2_12_6 : std_logic;
signal \c0.n10929\ : std_logic;
signal \c0.n10929_cascade_\ : std_logic;
signal \c0.n17823\ : std_logic;
signal \c0.n17853\ : std_logic;
signal \c0.n17823_cascade_\ : std_logic;
signal \c0.n17895\ : std_logic;
signal \c0.n17_adj_2401_cascade_\ : std_logic;
signal \c0.n17914\ : std_logic;
signal \c0.data_out_frame2_20_6\ : std_logic;
signal \c0.n10703\ : std_logic;
signal data_out_frame2_14_4 : std_logic;
signal \c0.n10825\ : std_logic;
signal \c0.data_out_frame2_0_5\ : std_logic;
signal data_out_frame2_8_1 : std_logic;
signal data_out_frame2_12_7 : std_logic;
signal rand_data_5 : std_logic;
signal data_out_frame2_12_5 : std_logic;
signal data_out_frame2_6_3 : std_logic;
signal \c0.n5_adj_2381\ : std_logic;
signal data_out_frame2_6_1 : std_logic;
signal \c0.n30_adj_2434\ : std_logic;
signal data_out_frame2_7_3 : std_logic;
signal \c0.data_out_frame2_0_3\ : std_logic;
signal data_out_frame2_14_3 : std_logic;
signal data_out_frame2_15_4 : std_logic;
signal data_out_frame2_7_4 : std_logic;
signal \c0.n10710\ : std_logic;
signal \c0.n10710_cascade_\ : std_logic;
signal \c0.n18_adj_2402\ : std_logic;
signal \c0.n20_adj_2404\ : std_logic;
signal data_out_frame2_6_5 : std_logic;
signal data_out_frame2_7_5 : std_logic;
signal \c0.n5_adj_2386\ : std_logic;
signal data_out_frame2_13_5 : std_logic;
signal data_out_frame2_10_7 : std_logic;
signal \c0.n10877\ : std_logic;
signal \c0.n10593_cascade_\ : std_logic;
signal \c0.n14\ : std_logic;
signal data_out_frame2_7_6 : std_logic;
signal data_out_frame2_5_7 : std_logic;
signal data_out_frame2_9_5 : std_logic;
signal data_out_frame2_9_3 : std_logic;
signal \c0.n17810\ : std_logic;
signal data_out_frame2_11_2 : std_logic;
signal data_out_frame2_11_3 : std_logic;
signal data_out_frame2_11_1 : std_logic;
signal \c0.n17798\ : std_logic;
signal \c0.n17751\ : std_logic;
signal \c0.n17868\ : std_logic;
signal \c0.n17798_cascade_\ : std_logic;
signal \c0.n17902\ : std_logic;
signal \c0.n18_adj_2393\ : std_logic;
signal data_out_frame2_16_5 : std_logic;
signal \c0.n24_adj_2394_cascade_\ : std_logic;
signal data_out_frame2_15_5 : std_logic;
signal \c0.n17920\ : std_logic;
signal \c0.n22_adj_2395\ : std_logic;
signal \c0.n26_adj_2396_cascade_\ : std_logic;
signal \c0.n17917\ : std_logic;
signal \c0.data_out_frame2_20_7\ : std_logic;
signal \c0.n10778\ : std_logic;
signal \c0.n17871\ : std_logic;
signal \c0.n14_adj_2406_cascade_\ : std_logic;
signal \c0.n10583\ : std_logic;
signal data_out_frame2_11_5 : std_logic;
signal data_out_frame2_12_4 : std_logic;
signal \c0.n17780\ : std_logic;
signal \c0.n15_adj_2407\ : std_logic;
signal data_out_frame2_5_4 : std_logic;
signal \c0.n17856\ : std_logic;
signal data_out_frame2_16_2 : std_logic;
signal data_out_frame2_9_2 : std_logic;
signal \c0.n10887\ : std_logic;
signal \c0.n16_adj_2399\ : std_logic;
signal data_out_frame2_10_0 : std_logic;
signal data_out_frame2_11_0 : std_logic;
signal data_out_frame2_9_0 : std_logic;
signal \c0.n18891_cascade_\ : std_logic;
signal data_out_frame2_8_0 : std_logic;
signal data_out_frame2_14_0 : std_logic;
signal data_out_frame2_15_0 : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal data_out_frame2_13_0 : std_logic;
signal \c0.n18897_cascade_\ : std_logic;
signal data_out_frame2_12_0 : std_logic;
signal \c0.n18060\ : std_logic;
signal \c0.n18057_cascade_\ : std_logic;
signal \c0.n18374\ : std_logic;
signal \c0.n18723_cascade_\ : std_logic;
signal \c0.n6_adj_2275\ : std_logic;
signal \c0.n22_adj_2373\ : std_logic;
signal \c0.n18726_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal \c0.n18160\ : std_logic;
signal \c0.n18161\ : std_logic;
signal \c0.n18067\ : std_logic;
signal \c0.n18771_cascade_\ : std_logic;
signal \c0.n18068\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.n18774_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.tx2.n9639\ : std_logic;
signal \c0.n18669\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal data_out_frame2_16_4 : std_logic;
signal \c0.data_out_frame2_20_4\ : std_logic;
signal \c0.n7263\ : std_logic;
signal \c0.n18672_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n22_adj_2243\ : std_logic;
signal rand_setpoint_14 : std_logic;
signal \c0.n11016\ : std_logic;
signal n2732 : std_logic;
signal \c0.data_out_7_6\ : std_logic;
signal \UART_TRANSMITTER_state_2\ : std_logic;
signal \UART_TRANSMITTER_state_0\ : std_logic;
signal \UART_TRANSMITTER_state_1\ : std_logic;
signal \data_out_10__7__N_110\ : std_logic;
signal rand_setpoint_0 : std_logic;
signal \data_out_10__7__N_110_cascade_\ : std_logic;
signal data_out_8_0 : std_logic;
signal data_out_frame2_8_4 : std_logic;
signal \c0.n10788\ : std_logic;
signal data_out_frame2_10_6 : std_logic;
signal \c0.n18_adj_2437\ : std_logic;
signal data_out_frame2_7_2 : std_logic;
signal data_out_frame2_15_2 : std_logic;
signal \c0.data_out_frame2_0_2\ : std_logic;
signal data_out_frame2_14_2 : std_logic;
signal \c0.n6_adj_2409_cascade_\ : std_logic;
signal data_out_frame2_11_4 : std_logic;
signal \c0.n17905\ : std_logic;
signal rand_data_12 : std_logic;
signal n11114 : std_logic;
signal data_out_frame2_17_4 : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_22_wire\ : std_logic;
signal \PIN_23_wire\ : std_logic;
signal \PIN_24_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    PIN_1 <= \PIN_1_wire\;
    PIN_22 <= \PIN_22_wire\;
    PIN_23 <= \PIN_23_wire\;
    PIN_24 <= \PIN_24_wire\;
    PIN_2 <= \PIN_2_wire\;
    PIN_3 <= \PIN_3_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51094\,
            DIN => \N__51093\,
            DOUT => \N__51092\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51094\,
            PADOUT => \N__51093\,
            PADIN => \N__51092\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22809\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51085\,
            DIN => \N__51084\,
            DOUT => \N__51083\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51085\,
            PADOUT => \N__51084\,
            PADIN => \N__51083\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24903\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51076\,
            DIN => \N__51075\,
            DOUT => \N__51074\,
            PACKAGEPIN => \PIN_22_wire\
        );

    \PIN_22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51076\,
            PADOUT => \N__51075\,
            PADIN => \N__51074\,
            CLOCKENABLE => \N__32793\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35292\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__49893\,
            OUTPUTENABLE => '0'
        );

    \PIN_23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51067\,
            DIN => \N__51066\,
            DOUT => \N__51065\,
            PACKAGEPIN => \PIN_23_wire\
        );

    \PIN_23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51067\,
            PADOUT => \N__51066\,
            PADIN => \N__51065\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35742\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51058\,
            DIN => \N__51057\,
            DOUT => \N__51056\,
            PACKAGEPIN => \PIN_24_wire\
        );

    \PIN_24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51058\,
            PADOUT => \N__51057\,
            PADIN => \N__51056\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35778\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51049\,
            DIN => \N__51048\,
            DOUT => \N__51047\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51049\,
            PADOUT => \N__51048\,
            PADIN => \N__51047\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__18558\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51040\,
            DIN => \N__51039\,
            DOUT => \N__51038\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51040\,
            PADOUT => \N__51039\,
            PADIN => \N__51038\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22797\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51031\,
            DIN => \N__51030\,
            DOUT => \N__51029\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51031\,
            PADOUT => \N__51030\,
            PADIN => \N__51029\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51022\,
            DIN => \N__51021\,
            DOUT => \N__51020\,
            PACKAGEPIN => PIN_4
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51022\,
            PADOUT => \N__51021\,
            PADIN => \N__51020\,
            CLOCKENABLE => 'H',
            DIN0 => hall1,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51013\,
            DIN => \N__51012\,
            DOUT => \N__51011\,
            PACKAGEPIN => PIN_5
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51013\,
            PADOUT => \N__51012\,
            PADIN => \N__51011\,
            CLOCKENABLE => 'H',
            DIN0 => hall2,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51004\,
            DIN => \N__51003\,
            DOUT => \N__51002\,
            PACKAGEPIN => PIN_6
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51004\,
            PADOUT => \N__51003\,
            PADIN => \N__51002\,
            CLOCKENABLE => 'H',
            DIN0 => hall3,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50995\,
            DIN => \N__50994\,
            DOUT => \N__50993\,
            PACKAGEPIN => PIN_12
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50995\,
            PADOUT => \N__50994\,
            PADIN => \N__50993\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__49822\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50986\,
            DIN => \N__50985\,
            DOUT => \N__50984\,
            PACKAGEPIN => PIN_11
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50986\,
            PADOUT => \N__50985\,
            PADIN => \N__50984\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22769\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__22734\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50977\,
            DIN => \N__50976\,
            DOUT => \N__50975\,
            PACKAGEPIN => PIN_10
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50977\,
            PADOUT => \N__50976\,
            PADIN => \N__50975\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29367\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__29121\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50968\,
            DIN => \N__50967\,
            DOUT => \N__50966\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50968\,
            PADOUT => \N__50967\,
            PADIN => \N__50966\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__12716\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50946\
        );

    \I__12715\ : LocalMux
    port map (
            O => \N__50946\,
            I => \N__50942\
        );

    \I__12714\ : CascadeMux
    port map (
            O => \N__50945\,
            I => \N__50939\
        );

    \I__12713\ : Span4Mux_v
    port map (
            O => \N__50942\,
            I => \N__50936\
        );

    \I__12712\ : InMux
    port map (
            O => \N__50939\,
            I => \N__50933\
        );

    \I__12711\ : Odrv4
    port map (
            O => \N__50936\,
            I => rand_setpoint_0
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__50933\,
            I => rand_setpoint_0
        );

    \I__12709\ : CascadeMux
    port map (
            O => \N__50928\,
            I => \data_out_10__7__N_110_cascade_\
        );

    \I__12708\ : InMux
    port map (
            O => \N__50925\,
            I => \N__50918\
        );

    \I__12707\ : InMux
    port map (
            O => \N__50924\,
            I => \N__50918\
        );

    \I__12706\ : CascadeMux
    port map (
            O => \N__50923\,
            I => \N__50915\
        );

    \I__12705\ : LocalMux
    port map (
            O => \N__50918\,
            I => \N__50911\
        );

    \I__12704\ : InMux
    port map (
            O => \N__50915\,
            I => \N__50905\
        );

    \I__12703\ : InMux
    port map (
            O => \N__50914\,
            I => \N__50905\
        );

    \I__12702\ : Span4Mux_h
    port map (
            O => \N__50911\,
            I => \N__50902\
        );

    \I__12701\ : InMux
    port map (
            O => \N__50910\,
            I => \N__50899\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__50905\,
            I => \N__50896\
        );

    \I__12699\ : Span4Mux_h
    port map (
            O => \N__50902\,
            I => \N__50893\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__50899\,
            I => data_out_8_0
        );

    \I__12697\ : Odrv12
    port map (
            O => \N__50896\,
            I => data_out_8_0
        );

    \I__12696\ : Odrv4
    port map (
            O => \N__50893\,
            I => data_out_8_0
        );

    \I__12695\ : InMux
    port map (
            O => \N__50886\,
            I => \N__50882\
        );

    \I__12694\ : InMux
    port map (
            O => \N__50885\,
            I => \N__50878\
        );

    \I__12693\ : LocalMux
    port map (
            O => \N__50882\,
            I => \N__50875\
        );

    \I__12692\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50872\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__50878\,
            I => \N__50865\
        );

    \I__12690\ : Span4Mux_v
    port map (
            O => \N__50875\,
            I => \N__50860\
        );

    \I__12689\ : LocalMux
    port map (
            O => \N__50872\,
            I => \N__50860\
        );

    \I__12688\ : InMux
    port map (
            O => \N__50871\,
            I => \N__50857\
        );

    \I__12687\ : InMux
    port map (
            O => \N__50870\,
            I => \N__50854\
        );

    \I__12686\ : InMux
    port map (
            O => \N__50869\,
            I => \N__50851\
        );

    \I__12685\ : InMux
    port map (
            O => \N__50868\,
            I => \N__50848\
        );

    \I__12684\ : Span4Mux_v
    port map (
            O => \N__50865\,
            I => \N__50839\
        );

    \I__12683\ : Span4Mux_h
    port map (
            O => \N__50860\,
            I => \N__50839\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__50857\,
            I => \N__50839\
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__50854\,
            I => \N__50839\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__50851\,
            I => data_out_frame2_8_4
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__50848\,
            I => data_out_frame2_8_4
        );

    \I__12678\ : Odrv4
    port map (
            O => \N__50839\,
            I => data_out_frame2_8_4
        );

    \I__12677\ : CascadeMux
    port map (
            O => \N__50832\,
            I => \N__50829\
        );

    \I__12676\ : InMux
    port map (
            O => \N__50829\,
            I => \N__50826\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__50826\,
            I => \c0.n10788\
        );

    \I__12674\ : InMux
    port map (
            O => \N__50823\,
            I => \N__50816\
        );

    \I__12673\ : InMux
    port map (
            O => \N__50822\,
            I => \N__50813\
        );

    \I__12672\ : InMux
    port map (
            O => \N__50821\,
            I => \N__50810\
        );

    \I__12671\ : InMux
    port map (
            O => \N__50820\,
            I => \N__50807\
        );

    \I__12670\ : InMux
    port map (
            O => \N__50819\,
            I => \N__50804\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__50816\,
            I => \N__50801\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__50813\,
            I => \N__50798\
        );

    \I__12667\ : LocalMux
    port map (
            O => \N__50810\,
            I => \N__50793\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__50807\,
            I => \N__50793\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__50804\,
            I => \N__50790\
        );

    \I__12664\ : Span4Mux_s0_v
    port map (
            O => \N__50801\,
            I => \N__50786\
        );

    \I__12663\ : Span4Mux_h
    port map (
            O => \N__50798\,
            I => \N__50779\
        );

    \I__12662\ : Span4Mux_v
    port map (
            O => \N__50793\,
            I => \N__50779\
        );

    \I__12661\ : Span4Mux_s1_v
    port map (
            O => \N__50790\,
            I => \N__50779\
        );

    \I__12660\ : InMux
    port map (
            O => \N__50789\,
            I => \N__50776\
        );

    \I__12659\ : Span4Mux_v
    port map (
            O => \N__50786\,
            I => \N__50773\
        );

    \I__12658\ : Span4Mux_h
    port map (
            O => \N__50779\,
            I => \N__50770\
        );

    \I__12657\ : LocalMux
    port map (
            O => \N__50776\,
            I => data_out_frame2_10_6
        );

    \I__12656\ : Odrv4
    port map (
            O => \N__50773\,
            I => data_out_frame2_10_6
        );

    \I__12655\ : Odrv4
    port map (
            O => \N__50770\,
            I => data_out_frame2_10_6
        );

    \I__12654\ : InMux
    port map (
            O => \N__50763\,
            I => \N__50760\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__50760\,
            I => \c0.n18_adj_2437\
        );

    \I__12652\ : InMux
    port map (
            O => \N__50757\,
            I => \N__50753\
        );

    \I__12651\ : InMux
    port map (
            O => \N__50756\,
            I => \N__50750\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__50753\,
            I => \N__50747\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__50750\,
            I => \N__50744\
        );

    \I__12648\ : Span4Mux_s2_v
    port map (
            O => \N__50747\,
            I => \N__50739\
        );

    \I__12647\ : Span4Mux_h
    port map (
            O => \N__50744\,
            I => \N__50736\
        );

    \I__12646\ : CascadeMux
    port map (
            O => \N__50743\,
            I => \N__50733\
        );

    \I__12645\ : InMux
    port map (
            O => \N__50742\,
            I => \N__50730\
        );

    \I__12644\ : Span4Mux_h
    port map (
            O => \N__50739\,
            I => \N__50727\
        );

    \I__12643\ : Span4Mux_h
    port map (
            O => \N__50736\,
            I => \N__50724\
        );

    \I__12642\ : InMux
    port map (
            O => \N__50733\,
            I => \N__50721\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__50730\,
            I => data_out_frame2_7_2
        );

    \I__12640\ : Odrv4
    port map (
            O => \N__50727\,
            I => data_out_frame2_7_2
        );

    \I__12639\ : Odrv4
    port map (
            O => \N__50724\,
            I => data_out_frame2_7_2
        );

    \I__12638\ : LocalMux
    port map (
            O => \N__50721\,
            I => data_out_frame2_7_2
        );

    \I__12637\ : InMux
    port map (
            O => \N__50712\,
            I => \N__50707\
        );

    \I__12636\ : InMux
    port map (
            O => \N__50711\,
            I => \N__50704\
        );

    \I__12635\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50699\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__50707\,
            I => \N__50696\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__50704\,
            I => \N__50693\
        );

    \I__12632\ : InMux
    port map (
            O => \N__50703\,
            I => \N__50690\
        );

    \I__12631\ : InMux
    port map (
            O => \N__50702\,
            I => \N__50687\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__50699\,
            I => data_out_frame2_15_2
        );

    \I__12629\ : Odrv12
    port map (
            O => \N__50696\,
            I => data_out_frame2_15_2
        );

    \I__12628\ : Odrv4
    port map (
            O => \N__50693\,
            I => data_out_frame2_15_2
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__50690\,
            I => data_out_frame2_15_2
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__50687\,
            I => data_out_frame2_15_2
        );

    \I__12625\ : InMux
    port map (
            O => \N__50676\,
            I => \N__50673\
        );

    \I__12624\ : LocalMux
    port map (
            O => \N__50673\,
            I => \N__50668\
        );

    \I__12623\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50665\
        );

    \I__12622\ : InMux
    port map (
            O => \N__50671\,
            I => \N__50661\
        );

    \I__12621\ : Span4Mux_h
    port map (
            O => \N__50668\,
            I => \N__50656\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__50665\,
            I => \N__50656\
        );

    \I__12619\ : CascadeMux
    port map (
            O => \N__50664\,
            I => \N__50652\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__50661\,
            I => \N__50649\
        );

    \I__12617\ : Span4Mux_s3_v
    port map (
            O => \N__50656\,
            I => \N__50646\
        );

    \I__12616\ : InMux
    port map (
            O => \N__50655\,
            I => \N__50643\
        );

    \I__12615\ : InMux
    port map (
            O => \N__50652\,
            I => \N__50640\
        );

    \I__12614\ : Span4Mux_h
    port map (
            O => \N__50649\,
            I => \N__50637\
        );

    \I__12613\ : Span4Mux_h
    port map (
            O => \N__50646\,
            I => \N__50634\
        );

    \I__12612\ : LocalMux
    port map (
            O => \N__50643\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__50640\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__12610\ : Odrv4
    port map (
            O => \N__50637\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__12609\ : Odrv4
    port map (
            O => \N__50634\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__12608\ : InMux
    port map (
            O => \N__50625\,
            I => \N__50622\
        );

    \I__12607\ : LocalMux
    port map (
            O => \N__50622\,
            I => \N__50617\
        );

    \I__12606\ : CascadeMux
    port map (
            O => \N__50621\,
            I => \N__50614\
        );

    \I__12605\ : InMux
    port map (
            O => \N__50620\,
            I => \N__50610\
        );

    \I__12604\ : Span4Mux_h
    port map (
            O => \N__50617\,
            I => \N__50607\
        );

    \I__12603\ : InMux
    port map (
            O => \N__50614\,
            I => \N__50604\
        );

    \I__12602\ : InMux
    port map (
            O => \N__50613\,
            I => \N__50601\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__50610\,
            I => \N__50594\
        );

    \I__12600\ : Span4Mux_h
    port map (
            O => \N__50607\,
            I => \N__50594\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__50604\,
            I => \N__50594\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__50601\,
            I => data_out_frame2_14_2
        );

    \I__12597\ : Odrv4
    port map (
            O => \N__50594\,
            I => data_out_frame2_14_2
        );

    \I__12596\ : CascadeMux
    port map (
            O => \N__50589\,
            I => \c0.n6_adj_2409_cascade_\
        );

    \I__12595\ : InMux
    port map (
            O => \N__50586\,
            I => \N__50582\
        );

    \I__12594\ : InMux
    port map (
            O => \N__50585\,
            I => \N__50578\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__50582\,
            I => \N__50575\
        );

    \I__12592\ : CascadeMux
    port map (
            O => \N__50581\,
            I => \N__50572\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__50578\,
            I => \N__50568\
        );

    \I__12590\ : Span4Mux_h
    port map (
            O => \N__50575\,
            I => \N__50565\
        );

    \I__12589\ : InMux
    port map (
            O => \N__50572\,
            I => \N__50560\
        );

    \I__12588\ : InMux
    port map (
            O => \N__50571\,
            I => \N__50560\
        );

    \I__12587\ : Odrv4
    port map (
            O => \N__50568\,
            I => data_out_frame2_11_4
        );

    \I__12586\ : Odrv4
    port map (
            O => \N__50565\,
            I => data_out_frame2_11_4
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__50560\,
            I => data_out_frame2_11_4
        );

    \I__12584\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50549\
        );

    \I__12583\ : CascadeMux
    port map (
            O => \N__50552\,
            I => \N__50546\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__50549\,
            I => \N__50543\
        );

    \I__12581\ : InMux
    port map (
            O => \N__50546\,
            I => \N__50540\
        );

    \I__12580\ : Span4Mux_s3_v
    port map (
            O => \N__50543\,
            I => \N__50537\
        );

    \I__12579\ : LocalMux
    port map (
            O => \N__50540\,
            I => \N__50534\
        );

    \I__12578\ : Odrv4
    port map (
            O => \N__50537\,
            I => \c0.n17905\
        );

    \I__12577\ : Odrv4
    port map (
            O => \N__50534\,
            I => \c0.n17905\
        );

    \I__12576\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50526\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__50526\,
            I => \N__50520\
        );

    \I__12574\ : InMux
    port map (
            O => \N__50525\,
            I => \N__50517\
        );

    \I__12573\ : InMux
    port map (
            O => \N__50524\,
            I => \N__50514\
        );

    \I__12572\ : InMux
    port map (
            O => \N__50523\,
            I => \N__50511\
        );

    \I__12571\ : Span4Mux_h
    port map (
            O => \N__50520\,
            I => \N__50506\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__50517\,
            I => \N__50506\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__50514\,
            I => \N__50501\
        );

    \I__12568\ : LocalMux
    port map (
            O => \N__50511\,
            I => \N__50498\
        );

    \I__12567\ : Span4Mux_h
    port map (
            O => \N__50506\,
            I => \N__50495\
        );

    \I__12566\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50492\
        );

    \I__12565\ : InMux
    port map (
            O => \N__50504\,
            I => \N__50489\
        );

    \I__12564\ : Span4Mux_v
    port map (
            O => \N__50501\,
            I => \N__50484\
        );

    \I__12563\ : Span4Mux_v
    port map (
            O => \N__50498\,
            I => \N__50484\
        );

    \I__12562\ : Odrv4
    port map (
            O => \N__50495\,
            I => rand_data_12
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__50492\,
            I => rand_data_12
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__50489\,
            I => rand_data_12
        );

    \I__12559\ : Odrv4
    port map (
            O => \N__50484\,
            I => rand_data_12
        );

    \I__12558\ : CEMux
    port map (
            O => \N__50475\,
            I => \N__50470\
        );

    \I__12557\ : CEMux
    port map (
            O => \N__50474\,
            I => \N__50459\
        );

    \I__12556\ : InMux
    port map (
            O => \N__50473\,
            I => \N__50456\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__50470\,
            I => \N__50441\
        );

    \I__12554\ : CEMux
    port map (
            O => \N__50469\,
            I => \N__50438\
        );

    \I__12553\ : CEMux
    port map (
            O => \N__50468\,
            I => \N__50420\
        );

    \I__12552\ : CEMux
    port map (
            O => \N__50467\,
            I => \N__50416\
        );

    \I__12551\ : CEMux
    port map (
            O => \N__50466\,
            I => \N__50413\
        );

    \I__12550\ : InMux
    port map (
            O => \N__50465\,
            I => \N__50406\
        );

    \I__12549\ : InMux
    port map (
            O => \N__50464\,
            I => \N__50406\
        );

    \I__12548\ : InMux
    port map (
            O => \N__50463\,
            I => \N__50406\
        );

    \I__12547\ : CEMux
    port map (
            O => \N__50462\,
            I => \N__50395\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__50459\,
            I => \N__50392\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__50456\,
            I => \N__50389\
        );

    \I__12544\ : InMux
    port map (
            O => \N__50455\,
            I => \N__50380\
        );

    \I__12543\ : InMux
    port map (
            O => \N__50454\,
            I => \N__50380\
        );

    \I__12542\ : InMux
    port map (
            O => \N__50453\,
            I => \N__50380\
        );

    \I__12541\ : InMux
    port map (
            O => \N__50452\,
            I => \N__50380\
        );

    \I__12540\ : InMux
    port map (
            O => \N__50451\,
            I => \N__50377\
        );

    \I__12539\ : InMux
    port map (
            O => \N__50450\,
            I => \N__50374\
        );

    \I__12538\ : InMux
    port map (
            O => \N__50449\,
            I => \N__50371\
        );

    \I__12537\ : InMux
    port map (
            O => \N__50448\,
            I => \N__50364\
        );

    \I__12536\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50364\
        );

    \I__12535\ : InMux
    port map (
            O => \N__50446\,
            I => \N__50364\
        );

    \I__12534\ : InMux
    port map (
            O => \N__50445\,
            I => \N__50361\
        );

    \I__12533\ : CEMux
    port map (
            O => \N__50444\,
            I => \N__50351\
        );

    \I__12532\ : Span4Mux_s2_v
    port map (
            O => \N__50441\,
            I => \N__50345\
        );

    \I__12531\ : LocalMux
    port map (
            O => \N__50438\,
            I => \N__50345\
        );

    \I__12530\ : CEMux
    port map (
            O => \N__50437\,
            I => \N__50342\
        );

    \I__12529\ : InMux
    port map (
            O => \N__50436\,
            I => \N__50339\
        );

    \I__12528\ : InMux
    port map (
            O => \N__50435\,
            I => \N__50336\
        );

    \I__12527\ : InMux
    port map (
            O => \N__50434\,
            I => \N__50327\
        );

    \I__12526\ : InMux
    port map (
            O => \N__50433\,
            I => \N__50327\
        );

    \I__12525\ : InMux
    port map (
            O => \N__50432\,
            I => \N__50327\
        );

    \I__12524\ : InMux
    port map (
            O => \N__50431\,
            I => \N__50327\
        );

    \I__12523\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50324\
        );

    \I__12522\ : InMux
    port map (
            O => \N__50429\,
            I => \N__50317\
        );

    \I__12521\ : InMux
    port map (
            O => \N__50428\,
            I => \N__50317\
        );

    \I__12520\ : InMux
    port map (
            O => \N__50427\,
            I => \N__50317\
        );

    \I__12519\ : CEMux
    port map (
            O => \N__50426\,
            I => \N__50310\
        );

    \I__12518\ : InMux
    port map (
            O => \N__50425\,
            I => \N__50303\
        );

    \I__12517\ : InMux
    port map (
            O => \N__50424\,
            I => \N__50303\
        );

    \I__12516\ : InMux
    port map (
            O => \N__50423\,
            I => \N__50303\
        );

    \I__12515\ : LocalMux
    port map (
            O => \N__50420\,
            I => \N__50294\
        );

    \I__12514\ : CEMux
    port map (
            O => \N__50419\,
            I => \N__50291\
        );

    \I__12513\ : LocalMux
    port map (
            O => \N__50416\,
            I => \N__50288\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__50413\,
            I => \N__50285\
        );

    \I__12511\ : LocalMux
    port map (
            O => \N__50406\,
            I => \N__50282\
        );

    \I__12510\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50277\
        );

    \I__12509\ : InMux
    port map (
            O => \N__50404\,
            I => \N__50277\
        );

    \I__12508\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50264\
        );

    \I__12507\ : InMux
    port map (
            O => \N__50402\,
            I => \N__50264\
        );

    \I__12506\ : InMux
    port map (
            O => \N__50401\,
            I => \N__50264\
        );

    \I__12505\ : InMux
    port map (
            O => \N__50400\,
            I => \N__50264\
        );

    \I__12504\ : InMux
    port map (
            O => \N__50399\,
            I => \N__50264\
        );

    \I__12503\ : InMux
    port map (
            O => \N__50398\,
            I => \N__50264\
        );

    \I__12502\ : LocalMux
    port map (
            O => \N__50395\,
            I => \N__50237\
        );

    \I__12501\ : Span4Mux_s3_v
    port map (
            O => \N__50392\,
            I => \N__50234\
        );

    \I__12500\ : Span4Mux_s3_v
    port map (
            O => \N__50389\,
            I => \N__50229\
        );

    \I__12499\ : LocalMux
    port map (
            O => \N__50380\,
            I => \N__50229\
        );

    \I__12498\ : LocalMux
    port map (
            O => \N__50377\,
            I => \N__50226\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__50374\,
            I => \N__50219\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__50371\,
            I => \N__50219\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__50364\,
            I => \N__50219\
        );

    \I__12494\ : LocalMux
    port map (
            O => \N__50361\,
            I => \N__50216\
        );

    \I__12493\ : InMux
    port map (
            O => \N__50360\,
            I => \N__50201\
        );

    \I__12492\ : InMux
    port map (
            O => \N__50359\,
            I => \N__50201\
        );

    \I__12491\ : InMux
    port map (
            O => \N__50358\,
            I => \N__50201\
        );

    \I__12490\ : InMux
    port map (
            O => \N__50357\,
            I => \N__50201\
        );

    \I__12489\ : InMux
    port map (
            O => \N__50356\,
            I => \N__50201\
        );

    \I__12488\ : InMux
    port map (
            O => \N__50355\,
            I => \N__50201\
        );

    \I__12487\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50201\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__50351\,
            I => \N__50198\
        );

    \I__12485\ : CEMux
    port map (
            O => \N__50350\,
            I => \N__50195\
        );

    \I__12484\ : Span4Mux_v
    port map (
            O => \N__50345\,
            I => \N__50188\
        );

    \I__12483\ : LocalMux
    port map (
            O => \N__50342\,
            I => \N__50188\
        );

    \I__12482\ : LocalMux
    port map (
            O => \N__50339\,
            I => \N__50188\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__50336\,
            I => \N__50179\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__50327\,
            I => \N__50179\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__50324\,
            I => \N__50179\
        );

    \I__12478\ : LocalMux
    port map (
            O => \N__50317\,
            I => \N__50179\
        );

    \I__12477\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50170\
        );

    \I__12476\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50170\
        );

    \I__12475\ : InMux
    port map (
            O => \N__50314\,
            I => \N__50170\
        );

    \I__12474\ : InMux
    port map (
            O => \N__50313\,
            I => \N__50170\
        );

    \I__12473\ : LocalMux
    port map (
            O => \N__50310\,
            I => \N__50165\
        );

    \I__12472\ : LocalMux
    port map (
            O => \N__50303\,
            I => \N__50165\
        );

    \I__12471\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50152\
        );

    \I__12470\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50152\
        );

    \I__12469\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50152\
        );

    \I__12468\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50152\
        );

    \I__12467\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50152\
        );

    \I__12466\ : InMux
    port map (
            O => \N__50297\,
            I => \N__50152\
        );

    \I__12465\ : Span4Mux_v
    port map (
            O => \N__50294\,
            I => \N__50115\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__50291\,
            I => \N__50112\
        );

    \I__12463\ : Span4Mux_s3_v
    port map (
            O => \N__50288\,
            I => \N__50109\
        );

    \I__12462\ : Span4Mux_h
    port map (
            O => \N__50285\,
            I => \N__50100\
        );

    \I__12461\ : Span4Mux_v
    port map (
            O => \N__50282\,
            I => \N__50100\
        );

    \I__12460\ : LocalMux
    port map (
            O => \N__50277\,
            I => \N__50100\
        );

    \I__12459\ : LocalMux
    port map (
            O => \N__50264\,
            I => \N__50100\
        );

    \I__12458\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50091\
        );

    \I__12457\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50091\
        );

    \I__12456\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50091\
        );

    \I__12455\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50091\
        );

    \I__12454\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50076\
        );

    \I__12453\ : InMux
    port map (
            O => \N__50258\,
            I => \N__50076\
        );

    \I__12452\ : InMux
    port map (
            O => \N__50257\,
            I => \N__50076\
        );

    \I__12451\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50076\
        );

    \I__12450\ : InMux
    port map (
            O => \N__50255\,
            I => \N__50076\
        );

    \I__12449\ : InMux
    port map (
            O => \N__50254\,
            I => \N__50076\
        );

    \I__12448\ : InMux
    port map (
            O => \N__50253\,
            I => \N__50076\
        );

    \I__12447\ : InMux
    port map (
            O => \N__50252\,
            I => \N__50059\
        );

    \I__12446\ : InMux
    port map (
            O => \N__50251\,
            I => \N__50059\
        );

    \I__12445\ : InMux
    port map (
            O => \N__50250\,
            I => \N__50059\
        );

    \I__12444\ : InMux
    port map (
            O => \N__50249\,
            I => \N__50059\
        );

    \I__12443\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50059\
        );

    \I__12442\ : InMux
    port map (
            O => \N__50247\,
            I => \N__50059\
        );

    \I__12441\ : InMux
    port map (
            O => \N__50246\,
            I => \N__50059\
        );

    \I__12440\ : InMux
    port map (
            O => \N__50245\,
            I => \N__50059\
        );

    \I__12439\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50048\
        );

    \I__12438\ : InMux
    port map (
            O => \N__50243\,
            I => \N__50048\
        );

    \I__12437\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50048\
        );

    \I__12436\ : InMux
    port map (
            O => \N__50241\,
            I => \N__50048\
        );

    \I__12435\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50048\
        );

    \I__12434\ : Span4Mux_s3_v
    port map (
            O => \N__50237\,
            I => \N__50033\
        );

    \I__12433\ : Span4Mux_h
    port map (
            O => \N__50234\,
            I => \N__50033\
        );

    \I__12432\ : Span4Mux_v
    port map (
            O => \N__50229\,
            I => \N__50033\
        );

    \I__12431\ : Span4Mux_s3_v
    port map (
            O => \N__50226\,
            I => \N__50033\
        );

    \I__12430\ : Span4Mux_h
    port map (
            O => \N__50219\,
            I => \N__50033\
        );

    \I__12429\ : Span4Mux_h
    port map (
            O => \N__50216\,
            I => \N__50033\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__50201\,
            I => \N__50033\
        );

    \I__12427\ : Span4Mux_s2_v
    port map (
            O => \N__50198\,
            I => \N__50018\
        );

    \I__12426\ : LocalMux
    port map (
            O => \N__50195\,
            I => \N__50018\
        );

    \I__12425\ : Span4Mux_h
    port map (
            O => \N__50188\,
            I => \N__50018\
        );

    \I__12424\ : Span4Mux_v
    port map (
            O => \N__50179\,
            I => \N__50018\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__50170\,
            I => \N__50018\
        );

    \I__12422\ : Span4Mux_s2_v
    port map (
            O => \N__50165\,
            I => \N__50018\
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50018\
        );

    \I__12420\ : InMux
    port map (
            O => \N__50151\,
            I => \N__50001\
        );

    \I__12419\ : InMux
    port map (
            O => \N__50150\,
            I => \N__50001\
        );

    \I__12418\ : InMux
    port map (
            O => \N__50149\,
            I => \N__50001\
        );

    \I__12417\ : InMux
    port map (
            O => \N__50148\,
            I => \N__50001\
        );

    \I__12416\ : InMux
    port map (
            O => \N__50147\,
            I => \N__50001\
        );

    \I__12415\ : InMux
    port map (
            O => \N__50146\,
            I => \N__50001\
        );

    \I__12414\ : InMux
    port map (
            O => \N__50145\,
            I => \N__50001\
        );

    \I__12413\ : InMux
    port map (
            O => \N__50144\,
            I => \N__50001\
        );

    \I__12412\ : InMux
    port map (
            O => \N__50143\,
            I => \N__49988\
        );

    \I__12411\ : InMux
    port map (
            O => \N__50142\,
            I => \N__49988\
        );

    \I__12410\ : InMux
    port map (
            O => \N__50141\,
            I => \N__49988\
        );

    \I__12409\ : InMux
    port map (
            O => \N__50140\,
            I => \N__49988\
        );

    \I__12408\ : InMux
    port map (
            O => \N__50139\,
            I => \N__49988\
        );

    \I__12407\ : InMux
    port map (
            O => \N__50138\,
            I => \N__49988\
        );

    \I__12406\ : InMux
    port map (
            O => \N__50137\,
            I => \N__49973\
        );

    \I__12405\ : InMux
    port map (
            O => \N__50136\,
            I => \N__49973\
        );

    \I__12404\ : InMux
    port map (
            O => \N__50135\,
            I => \N__49973\
        );

    \I__12403\ : InMux
    port map (
            O => \N__50134\,
            I => \N__49973\
        );

    \I__12402\ : InMux
    port map (
            O => \N__50133\,
            I => \N__49973\
        );

    \I__12401\ : InMux
    port map (
            O => \N__50132\,
            I => \N__49973\
        );

    \I__12400\ : InMux
    port map (
            O => \N__50131\,
            I => \N__49973\
        );

    \I__12399\ : InMux
    port map (
            O => \N__50130\,
            I => \N__49958\
        );

    \I__12398\ : InMux
    port map (
            O => \N__50129\,
            I => \N__49958\
        );

    \I__12397\ : InMux
    port map (
            O => \N__50128\,
            I => \N__49958\
        );

    \I__12396\ : InMux
    port map (
            O => \N__50127\,
            I => \N__49958\
        );

    \I__12395\ : InMux
    port map (
            O => \N__50126\,
            I => \N__49958\
        );

    \I__12394\ : InMux
    port map (
            O => \N__50125\,
            I => \N__49958\
        );

    \I__12393\ : InMux
    port map (
            O => \N__50124\,
            I => \N__49958\
        );

    \I__12392\ : InMux
    port map (
            O => \N__50123\,
            I => \N__49945\
        );

    \I__12391\ : InMux
    port map (
            O => \N__50122\,
            I => \N__49945\
        );

    \I__12390\ : InMux
    port map (
            O => \N__50121\,
            I => \N__49945\
        );

    \I__12389\ : InMux
    port map (
            O => \N__50120\,
            I => \N__49945\
        );

    \I__12388\ : InMux
    port map (
            O => \N__50119\,
            I => \N__49945\
        );

    \I__12387\ : InMux
    port map (
            O => \N__50118\,
            I => \N__49945\
        );

    \I__12386\ : Odrv4
    port map (
            O => \N__50115\,
            I => n11114
        );

    \I__12385\ : Odrv4
    port map (
            O => \N__50112\,
            I => n11114
        );

    \I__12384\ : Odrv4
    port map (
            O => \N__50109\,
            I => n11114
        );

    \I__12383\ : Odrv4
    port map (
            O => \N__50100\,
            I => n11114
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__50091\,
            I => n11114
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__50076\,
            I => n11114
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__50059\,
            I => n11114
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__50048\,
            I => n11114
        );

    \I__12378\ : Odrv4
    port map (
            O => \N__50033\,
            I => n11114
        );

    \I__12377\ : Odrv4
    port map (
            O => \N__50018\,
            I => n11114
        );

    \I__12376\ : LocalMux
    port map (
            O => \N__50001\,
            I => n11114
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__49988\,
            I => n11114
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__49973\,
            I => n11114
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__49958\,
            I => n11114
        );

    \I__12372\ : LocalMux
    port map (
            O => \N__49945\,
            I => n11114
        );

    \I__12371\ : CascadeMux
    port map (
            O => \N__49914\,
            I => \N__49911\
        );

    \I__12370\ : InMux
    port map (
            O => \N__49911\,
            I => \N__49908\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__49908\,
            I => \N__49904\
        );

    \I__12368\ : InMux
    port map (
            O => \N__49907\,
            I => \N__49901\
        );

    \I__12367\ : Span4Mux_v
    port map (
            O => \N__49904\,
            I => \N__49898\
        );

    \I__12366\ : LocalMux
    port map (
            O => \N__49901\,
            I => data_out_frame2_17_4
        );

    \I__12365\ : Odrv4
    port map (
            O => \N__49898\,
            I => data_out_frame2_17_4
        );

    \I__12364\ : ClkMux
    port map (
            O => \N__49893\,
            I => \N__49206\
        );

    \I__12363\ : ClkMux
    port map (
            O => \N__49892\,
            I => \N__49206\
        );

    \I__12362\ : ClkMux
    port map (
            O => \N__49891\,
            I => \N__49206\
        );

    \I__12361\ : ClkMux
    port map (
            O => \N__49890\,
            I => \N__49206\
        );

    \I__12360\ : ClkMux
    port map (
            O => \N__49889\,
            I => \N__49206\
        );

    \I__12359\ : ClkMux
    port map (
            O => \N__49888\,
            I => \N__49206\
        );

    \I__12358\ : ClkMux
    port map (
            O => \N__49887\,
            I => \N__49206\
        );

    \I__12357\ : ClkMux
    port map (
            O => \N__49886\,
            I => \N__49206\
        );

    \I__12356\ : ClkMux
    port map (
            O => \N__49885\,
            I => \N__49206\
        );

    \I__12355\ : ClkMux
    port map (
            O => \N__49884\,
            I => \N__49206\
        );

    \I__12354\ : ClkMux
    port map (
            O => \N__49883\,
            I => \N__49206\
        );

    \I__12353\ : ClkMux
    port map (
            O => \N__49882\,
            I => \N__49206\
        );

    \I__12352\ : ClkMux
    port map (
            O => \N__49881\,
            I => \N__49206\
        );

    \I__12351\ : ClkMux
    port map (
            O => \N__49880\,
            I => \N__49206\
        );

    \I__12350\ : ClkMux
    port map (
            O => \N__49879\,
            I => \N__49206\
        );

    \I__12349\ : ClkMux
    port map (
            O => \N__49878\,
            I => \N__49206\
        );

    \I__12348\ : ClkMux
    port map (
            O => \N__49877\,
            I => \N__49206\
        );

    \I__12347\ : ClkMux
    port map (
            O => \N__49876\,
            I => \N__49206\
        );

    \I__12346\ : ClkMux
    port map (
            O => \N__49875\,
            I => \N__49206\
        );

    \I__12345\ : ClkMux
    port map (
            O => \N__49874\,
            I => \N__49206\
        );

    \I__12344\ : ClkMux
    port map (
            O => \N__49873\,
            I => \N__49206\
        );

    \I__12343\ : ClkMux
    port map (
            O => \N__49872\,
            I => \N__49206\
        );

    \I__12342\ : ClkMux
    port map (
            O => \N__49871\,
            I => \N__49206\
        );

    \I__12341\ : ClkMux
    port map (
            O => \N__49870\,
            I => \N__49206\
        );

    \I__12340\ : ClkMux
    port map (
            O => \N__49869\,
            I => \N__49206\
        );

    \I__12339\ : ClkMux
    port map (
            O => \N__49868\,
            I => \N__49206\
        );

    \I__12338\ : ClkMux
    port map (
            O => \N__49867\,
            I => \N__49206\
        );

    \I__12337\ : ClkMux
    port map (
            O => \N__49866\,
            I => \N__49206\
        );

    \I__12336\ : ClkMux
    port map (
            O => \N__49865\,
            I => \N__49206\
        );

    \I__12335\ : ClkMux
    port map (
            O => \N__49864\,
            I => \N__49206\
        );

    \I__12334\ : ClkMux
    port map (
            O => \N__49863\,
            I => \N__49206\
        );

    \I__12333\ : ClkMux
    port map (
            O => \N__49862\,
            I => \N__49206\
        );

    \I__12332\ : ClkMux
    port map (
            O => \N__49861\,
            I => \N__49206\
        );

    \I__12331\ : ClkMux
    port map (
            O => \N__49860\,
            I => \N__49206\
        );

    \I__12330\ : ClkMux
    port map (
            O => \N__49859\,
            I => \N__49206\
        );

    \I__12329\ : ClkMux
    port map (
            O => \N__49858\,
            I => \N__49206\
        );

    \I__12328\ : ClkMux
    port map (
            O => \N__49857\,
            I => \N__49206\
        );

    \I__12327\ : ClkMux
    port map (
            O => \N__49856\,
            I => \N__49206\
        );

    \I__12326\ : ClkMux
    port map (
            O => \N__49855\,
            I => \N__49206\
        );

    \I__12325\ : ClkMux
    port map (
            O => \N__49854\,
            I => \N__49206\
        );

    \I__12324\ : ClkMux
    port map (
            O => \N__49853\,
            I => \N__49206\
        );

    \I__12323\ : ClkMux
    port map (
            O => \N__49852\,
            I => \N__49206\
        );

    \I__12322\ : ClkMux
    port map (
            O => \N__49851\,
            I => \N__49206\
        );

    \I__12321\ : ClkMux
    port map (
            O => \N__49850\,
            I => \N__49206\
        );

    \I__12320\ : ClkMux
    port map (
            O => \N__49849\,
            I => \N__49206\
        );

    \I__12319\ : ClkMux
    port map (
            O => \N__49848\,
            I => \N__49206\
        );

    \I__12318\ : ClkMux
    port map (
            O => \N__49847\,
            I => \N__49206\
        );

    \I__12317\ : ClkMux
    port map (
            O => \N__49846\,
            I => \N__49206\
        );

    \I__12316\ : ClkMux
    port map (
            O => \N__49845\,
            I => \N__49206\
        );

    \I__12315\ : ClkMux
    port map (
            O => \N__49844\,
            I => \N__49206\
        );

    \I__12314\ : ClkMux
    port map (
            O => \N__49843\,
            I => \N__49206\
        );

    \I__12313\ : ClkMux
    port map (
            O => \N__49842\,
            I => \N__49206\
        );

    \I__12312\ : ClkMux
    port map (
            O => \N__49841\,
            I => \N__49206\
        );

    \I__12311\ : ClkMux
    port map (
            O => \N__49840\,
            I => \N__49206\
        );

    \I__12310\ : ClkMux
    port map (
            O => \N__49839\,
            I => \N__49206\
        );

    \I__12309\ : ClkMux
    port map (
            O => \N__49838\,
            I => \N__49206\
        );

    \I__12308\ : ClkMux
    port map (
            O => \N__49837\,
            I => \N__49206\
        );

    \I__12307\ : ClkMux
    port map (
            O => \N__49836\,
            I => \N__49206\
        );

    \I__12306\ : ClkMux
    port map (
            O => \N__49835\,
            I => \N__49206\
        );

    \I__12305\ : ClkMux
    port map (
            O => \N__49834\,
            I => \N__49206\
        );

    \I__12304\ : ClkMux
    port map (
            O => \N__49833\,
            I => \N__49206\
        );

    \I__12303\ : ClkMux
    port map (
            O => \N__49832\,
            I => \N__49206\
        );

    \I__12302\ : ClkMux
    port map (
            O => \N__49831\,
            I => \N__49206\
        );

    \I__12301\ : ClkMux
    port map (
            O => \N__49830\,
            I => \N__49206\
        );

    \I__12300\ : ClkMux
    port map (
            O => \N__49829\,
            I => \N__49206\
        );

    \I__12299\ : ClkMux
    port map (
            O => \N__49828\,
            I => \N__49206\
        );

    \I__12298\ : ClkMux
    port map (
            O => \N__49827\,
            I => \N__49206\
        );

    \I__12297\ : ClkMux
    port map (
            O => \N__49826\,
            I => \N__49206\
        );

    \I__12296\ : ClkMux
    port map (
            O => \N__49825\,
            I => \N__49206\
        );

    \I__12295\ : ClkMux
    port map (
            O => \N__49824\,
            I => \N__49206\
        );

    \I__12294\ : ClkMux
    port map (
            O => \N__49823\,
            I => \N__49206\
        );

    \I__12293\ : ClkMux
    port map (
            O => \N__49822\,
            I => \N__49206\
        );

    \I__12292\ : ClkMux
    port map (
            O => \N__49821\,
            I => \N__49206\
        );

    \I__12291\ : ClkMux
    port map (
            O => \N__49820\,
            I => \N__49206\
        );

    \I__12290\ : ClkMux
    port map (
            O => \N__49819\,
            I => \N__49206\
        );

    \I__12289\ : ClkMux
    port map (
            O => \N__49818\,
            I => \N__49206\
        );

    \I__12288\ : ClkMux
    port map (
            O => \N__49817\,
            I => \N__49206\
        );

    \I__12287\ : ClkMux
    port map (
            O => \N__49816\,
            I => \N__49206\
        );

    \I__12286\ : ClkMux
    port map (
            O => \N__49815\,
            I => \N__49206\
        );

    \I__12285\ : ClkMux
    port map (
            O => \N__49814\,
            I => \N__49206\
        );

    \I__12284\ : ClkMux
    port map (
            O => \N__49813\,
            I => \N__49206\
        );

    \I__12283\ : ClkMux
    port map (
            O => \N__49812\,
            I => \N__49206\
        );

    \I__12282\ : ClkMux
    port map (
            O => \N__49811\,
            I => \N__49206\
        );

    \I__12281\ : ClkMux
    port map (
            O => \N__49810\,
            I => \N__49206\
        );

    \I__12280\ : ClkMux
    port map (
            O => \N__49809\,
            I => \N__49206\
        );

    \I__12279\ : ClkMux
    port map (
            O => \N__49808\,
            I => \N__49206\
        );

    \I__12278\ : ClkMux
    port map (
            O => \N__49807\,
            I => \N__49206\
        );

    \I__12277\ : ClkMux
    port map (
            O => \N__49806\,
            I => \N__49206\
        );

    \I__12276\ : ClkMux
    port map (
            O => \N__49805\,
            I => \N__49206\
        );

    \I__12275\ : ClkMux
    port map (
            O => \N__49804\,
            I => \N__49206\
        );

    \I__12274\ : ClkMux
    port map (
            O => \N__49803\,
            I => \N__49206\
        );

    \I__12273\ : ClkMux
    port map (
            O => \N__49802\,
            I => \N__49206\
        );

    \I__12272\ : ClkMux
    port map (
            O => \N__49801\,
            I => \N__49206\
        );

    \I__12271\ : ClkMux
    port map (
            O => \N__49800\,
            I => \N__49206\
        );

    \I__12270\ : ClkMux
    port map (
            O => \N__49799\,
            I => \N__49206\
        );

    \I__12269\ : ClkMux
    port map (
            O => \N__49798\,
            I => \N__49206\
        );

    \I__12268\ : ClkMux
    port map (
            O => \N__49797\,
            I => \N__49206\
        );

    \I__12267\ : ClkMux
    port map (
            O => \N__49796\,
            I => \N__49206\
        );

    \I__12266\ : ClkMux
    port map (
            O => \N__49795\,
            I => \N__49206\
        );

    \I__12265\ : ClkMux
    port map (
            O => \N__49794\,
            I => \N__49206\
        );

    \I__12264\ : ClkMux
    port map (
            O => \N__49793\,
            I => \N__49206\
        );

    \I__12263\ : ClkMux
    port map (
            O => \N__49792\,
            I => \N__49206\
        );

    \I__12262\ : ClkMux
    port map (
            O => \N__49791\,
            I => \N__49206\
        );

    \I__12261\ : ClkMux
    port map (
            O => \N__49790\,
            I => \N__49206\
        );

    \I__12260\ : ClkMux
    port map (
            O => \N__49789\,
            I => \N__49206\
        );

    \I__12259\ : ClkMux
    port map (
            O => \N__49788\,
            I => \N__49206\
        );

    \I__12258\ : ClkMux
    port map (
            O => \N__49787\,
            I => \N__49206\
        );

    \I__12257\ : ClkMux
    port map (
            O => \N__49786\,
            I => \N__49206\
        );

    \I__12256\ : ClkMux
    port map (
            O => \N__49785\,
            I => \N__49206\
        );

    \I__12255\ : ClkMux
    port map (
            O => \N__49784\,
            I => \N__49206\
        );

    \I__12254\ : ClkMux
    port map (
            O => \N__49783\,
            I => \N__49206\
        );

    \I__12253\ : ClkMux
    port map (
            O => \N__49782\,
            I => \N__49206\
        );

    \I__12252\ : ClkMux
    port map (
            O => \N__49781\,
            I => \N__49206\
        );

    \I__12251\ : ClkMux
    port map (
            O => \N__49780\,
            I => \N__49206\
        );

    \I__12250\ : ClkMux
    port map (
            O => \N__49779\,
            I => \N__49206\
        );

    \I__12249\ : ClkMux
    port map (
            O => \N__49778\,
            I => \N__49206\
        );

    \I__12248\ : ClkMux
    port map (
            O => \N__49777\,
            I => \N__49206\
        );

    \I__12247\ : ClkMux
    port map (
            O => \N__49776\,
            I => \N__49206\
        );

    \I__12246\ : ClkMux
    port map (
            O => \N__49775\,
            I => \N__49206\
        );

    \I__12245\ : ClkMux
    port map (
            O => \N__49774\,
            I => \N__49206\
        );

    \I__12244\ : ClkMux
    port map (
            O => \N__49773\,
            I => \N__49206\
        );

    \I__12243\ : ClkMux
    port map (
            O => \N__49772\,
            I => \N__49206\
        );

    \I__12242\ : ClkMux
    port map (
            O => \N__49771\,
            I => \N__49206\
        );

    \I__12241\ : ClkMux
    port map (
            O => \N__49770\,
            I => \N__49206\
        );

    \I__12240\ : ClkMux
    port map (
            O => \N__49769\,
            I => \N__49206\
        );

    \I__12239\ : ClkMux
    port map (
            O => \N__49768\,
            I => \N__49206\
        );

    \I__12238\ : ClkMux
    port map (
            O => \N__49767\,
            I => \N__49206\
        );

    \I__12237\ : ClkMux
    port map (
            O => \N__49766\,
            I => \N__49206\
        );

    \I__12236\ : ClkMux
    port map (
            O => \N__49765\,
            I => \N__49206\
        );

    \I__12235\ : ClkMux
    port map (
            O => \N__49764\,
            I => \N__49206\
        );

    \I__12234\ : ClkMux
    port map (
            O => \N__49763\,
            I => \N__49206\
        );

    \I__12233\ : ClkMux
    port map (
            O => \N__49762\,
            I => \N__49206\
        );

    \I__12232\ : ClkMux
    port map (
            O => \N__49761\,
            I => \N__49206\
        );

    \I__12231\ : ClkMux
    port map (
            O => \N__49760\,
            I => \N__49206\
        );

    \I__12230\ : ClkMux
    port map (
            O => \N__49759\,
            I => \N__49206\
        );

    \I__12229\ : ClkMux
    port map (
            O => \N__49758\,
            I => \N__49206\
        );

    \I__12228\ : ClkMux
    port map (
            O => \N__49757\,
            I => \N__49206\
        );

    \I__12227\ : ClkMux
    port map (
            O => \N__49756\,
            I => \N__49206\
        );

    \I__12226\ : ClkMux
    port map (
            O => \N__49755\,
            I => \N__49206\
        );

    \I__12225\ : ClkMux
    port map (
            O => \N__49754\,
            I => \N__49206\
        );

    \I__12224\ : ClkMux
    port map (
            O => \N__49753\,
            I => \N__49206\
        );

    \I__12223\ : ClkMux
    port map (
            O => \N__49752\,
            I => \N__49206\
        );

    \I__12222\ : ClkMux
    port map (
            O => \N__49751\,
            I => \N__49206\
        );

    \I__12221\ : ClkMux
    port map (
            O => \N__49750\,
            I => \N__49206\
        );

    \I__12220\ : ClkMux
    port map (
            O => \N__49749\,
            I => \N__49206\
        );

    \I__12219\ : ClkMux
    port map (
            O => \N__49748\,
            I => \N__49206\
        );

    \I__12218\ : ClkMux
    port map (
            O => \N__49747\,
            I => \N__49206\
        );

    \I__12217\ : ClkMux
    port map (
            O => \N__49746\,
            I => \N__49206\
        );

    \I__12216\ : ClkMux
    port map (
            O => \N__49745\,
            I => \N__49206\
        );

    \I__12215\ : ClkMux
    port map (
            O => \N__49744\,
            I => \N__49206\
        );

    \I__12214\ : ClkMux
    port map (
            O => \N__49743\,
            I => \N__49206\
        );

    \I__12213\ : ClkMux
    port map (
            O => \N__49742\,
            I => \N__49206\
        );

    \I__12212\ : ClkMux
    port map (
            O => \N__49741\,
            I => \N__49206\
        );

    \I__12211\ : ClkMux
    port map (
            O => \N__49740\,
            I => \N__49206\
        );

    \I__12210\ : ClkMux
    port map (
            O => \N__49739\,
            I => \N__49206\
        );

    \I__12209\ : ClkMux
    port map (
            O => \N__49738\,
            I => \N__49206\
        );

    \I__12208\ : ClkMux
    port map (
            O => \N__49737\,
            I => \N__49206\
        );

    \I__12207\ : ClkMux
    port map (
            O => \N__49736\,
            I => \N__49206\
        );

    \I__12206\ : ClkMux
    port map (
            O => \N__49735\,
            I => \N__49206\
        );

    \I__12205\ : ClkMux
    port map (
            O => \N__49734\,
            I => \N__49206\
        );

    \I__12204\ : ClkMux
    port map (
            O => \N__49733\,
            I => \N__49206\
        );

    \I__12203\ : ClkMux
    port map (
            O => \N__49732\,
            I => \N__49206\
        );

    \I__12202\ : ClkMux
    port map (
            O => \N__49731\,
            I => \N__49206\
        );

    \I__12201\ : ClkMux
    port map (
            O => \N__49730\,
            I => \N__49206\
        );

    \I__12200\ : ClkMux
    port map (
            O => \N__49729\,
            I => \N__49206\
        );

    \I__12199\ : ClkMux
    port map (
            O => \N__49728\,
            I => \N__49206\
        );

    \I__12198\ : ClkMux
    port map (
            O => \N__49727\,
            I => \N__49206\
        );

    \I__12197\ : ClkMux
    port map (
            O => \N__49726\,
            I => \N__49206\
        );

    \I__12196\ : ClkMux
    port map (
            O => \N__49725\,
            I => \N__49206\
        );

    \I__12195\ : ClkMux
    port map (
            O => \N__49724\,
            I => \N__49206\
        );

    \I__12194\ : ClkMux
    port map (
            O => \N__49723\,
            I => \N__49206\
        );

    \I__12193\ : ClkMux
    port map (
            O => \N__49722\,
            I => \N__49206\
        );

    \I__12192\ : ClkMux
    port map (
            O => \N__49721\,
            I => \N__49206\
        );

    \I__12191\ : ClkMux
    port map (
            O => \N__49720\,
            I => \N__49206\
        );

    \I__12190\ : ClkMux
    port map (
            O => \N__49719\,
            I => \N__49206\
        );

    \I__12189\ : ClkMux
    port map (
            O => \N__49718\,
            I => \N__49206\
        );

    \I__12188\ : ClkMux
    port map (
            O => \N__49717\,
            I => \N__49206\
        );

    \I__12187\ : ClkMux
    port map (
            O => \N__49716\,
            I => \N__49206\
        );

    \I__12186\ : ClkMux
    port map (
            O => \N__49715\,
            I => \N__49206\
        );

    \I__12185\ : ClkMux
    port map (
            O => \N__49714\,
            I => \N__49206\
        );

    \I__12184\ : ClkMux
    port map (
            O => \N__49713\,
            I => \N__49206\
        );

    \I__12183\ : ClkMux
    port map (
            O => \N__49712\,
            I => \N__49206\
        );

    \I__12182\ : ClkMux
    port map (
            O => \N__49711\,
            I => \N__49206\
        );

    \I__12181\ : ClkMux
    port map (
            O => \N__49710\,
            I => \N__49206\
        );

    \I__12180\ : ClkMux
    port map (
            O => \N__49709\,
            I => \N__49206\
        );

    \I__12179\ : ClkMux
    port map (
            O => \N__49708\,
            I => \N__49206\
        );

    \I__12178\ : ClkMux
    port map (
            O => \N__49707\,
            I => \N__49206\
        );

    \I__12177\ : ClkMux
    port map (
            O => \N__49706\,
            I => \N__49206\
        );

    \I__12176\ : ClkMux
    port map (
            O => \N__49705\,
            I => \N__49206\
        );

    \I__12175\ : ClkMux
    port map (
            O => \N__49704\,
            I => \N__49206\
        );

    \I__12174\ : ClkMux
    port map (
            O => \N__49703\,
            I => \N__49206\
        );

    \I__12173\ : ClkMux
    port map (
            O => \N__49702\,
            I => \N__49206\
        );

    \I__12172\ : ClkMux
    port map (
            O => \N__49701\,
            I => \N__49206\
        );

    \I__12171\ : ClkMux
    port map (
            O => \N__49700\,
            I => \N__49206\
        );

    \I__12170\ : ClkMux
    port map (
            O => \N__49699\,
            I => \N__49206\
        );

    \I__12169\ : ClkMux
    port map (
            O => \N__49698\,
            I => \N__49206\
        );

    \I__12168\ : ClkMux
    port map (
            O => \N__49697\,
            I => \N__49206\
        );

    \I__12167\ : ClkMux
    port map (
            O => \N__49696\,
            I => \N__49206\
        );

    \I__12166\ : ClkMux
    port map (
            O => \N__49695\,
            I => \N__49206\
        );

    \I__12165\ : ClkMux
    port map (
            O => \N__49694\,
            I => \N__49206\
        );

    \I__12164\ : ClkMux
    port map (
            O => \N__49693\,
            I => \N__49206\
        );

    \I__12163\ : ClkMux
    port map (
            O => \N__49692\,
            I => \N__49206\
        );

    \I__12162\ : ClkMux
    port map (
            O => \N__49691\,
            I => \N__49206\
        );

    \I__12161\ : ClkMux
    port map (
            O => \N__49690\,
            I => \N__49206\
        );

    \I__12160\ : ClkMux
    port map (
            O => \N__49689\,
            I => \N__49206\
        );

    \I__12159\ : ClkMux
    port map (
            O => \N__49688\,
            I => \N__49206\
        );

    \I__12158\ : ClkMux
    port map (
            O => \N__49687\,
            I => \N__49206\
        );

    \I__12157\ : ClkMux
    port map (
            O => \N__49686\,
            I => \N__49206\
        );

    \I__12156\ : ClkMux
    port map (
            O => \N__49685\,
            I => \N__49206\
        );

    \I__12155\ : ClkMux
    port map (
            O => \N__49684\,
            I => \N__49206\
        );

    \I__12154\ : ClkMux
    port map (
            O => \N__49683\,
            I => \N__49206\
        );

    \I__12153\ : ClkMux
    port map (
            O => \N__49682\,
            I => \N__49206\
        );

    \I__12152\ : ClkMux
    port map (
            O => \N__49681\,
            I => \N__49206\
        );

    \I__12151\ : ClkMux
    port map (
            O => \N__49680\,
            I => \N__49206\
        );

    \I__12150\ : ClkMux
    port map (
            O => \N__49679\,
            I => \N__49206\
        );

    \I__12149\ : ClkMux
    port map (
            O => \N__49678\,
            I => \N__49206\
        );

    \I__12148\ : ClkMux
    port map (
            O => \N__49677\,
            I => \N__49206\
        );

    \I__12147\ : ClkMux
    port map (
            O => \N__49676\,
            I => \N__49206\
        );

    \I__12146\ : ClkMux
    port map (
            O => \N__49675\,
            I => \N__49206\
        );

    \I__12145\ : ClkMux
    port map (
            O => \N__49674\,
            I => \N__49206\
        );

    \I__12144\ : ClkMux
    port map (
            O => \N__49673\,
            I => \N__49206\
        );

    \I__12143\ : ClkMux
    port map (
            O => \N__49672\,
            I => \N__49206\
        );

    \I__12142\ : ClkMux
    port map (
            O => \N__49671\,
            I => \N__49206\
        );

    \I__12141\ : ClkMux
    port map (
            O => \N__49670\,
            I => \N__49206\
        );

    \I__12140\ : ClkMux
    port map (
            O => \N__49669\,
            I => \N__49206\
        );

    \I__12139\ : ClkMux
    port map (
            O => \N__49668\,
            I => \N__49206\
        );

    \I__12138\ : ClkMux
    port map (
            O => \N__49667\,
            I => \N__49206\
        );

    \I__12137\ : ClkMux
    port map (
            O => \N__49666\,
            I => \N__49206\
        );

    \I__12136\ : ClkMux
    port map (
            O => \N__49665\,
            I => \N__49206\
        );

    \I__12135\ : GlobalMux
    port map (
            O => \N__49206\,
            I => \N__49203\
        );

    \I__12134\ : gio2CtrlBuf
    port map (
            O => \N__49203\,
            I => \CLK_c\
        );

    \I__12133\ : InMux
    port map (
            O => \N__49200\,
            I => \N__49197\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__49197\,
            I => \N__49194\
        );

    \I__12131\ : Span4Mux_v
    port map (
            O => \N__49194\,
            I => \N__49191\
        );

    \I__12130\ : Span4Mux_s2_v
    port map (
            O => \N__49191\,
            I => \N__49188\
        );

    \I__12129\ : Span4Mux_h
    port map (
            O => \N__49188\,
            I => \N__49185\
        );

    \I__12128\ : Odrv4
    port map (
            O => \N__49185\,
            I => \c0.n22_adj_2373\
        );

    \I__12127\ : CascadeMux
    port map (
            O => \N__49182\,
            I => \c0.n18726_cascade_\
        );

    \I__12126\ : InMux
    port map (
            O => \N__49179\,
            I => \N__49176\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__49176\,
            I => \N__49173\
        );

    \I__12124\ : Odrv12
    port map (
            O => \N__49173\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__12123\ : InMux
    port map (
            O => \N__49170\,
            I => \N__49167\
        );

    \I__12122\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49164\
        );

    \I__12121\ : Span4Mux_h
    port map (
            O => \N__49164\,
            I => \N__49161\
        );

    \I__12120\ : Odrv4
    port map (
            O => \N__49161\,
            I => \c0.n18160\
        );

    \I__12119\ : CascadeMux
    port map (
            O => \N__49158\,
            I => \N__49155\
        );

    \I__12118\ : InMux
    port map (
            O => \N__49155\,
            I => \N__49152\
        );

    \I__12117\ : LocalMux
    port map (
            O => \N__49152\,
            I => \c0.n18161\
        );

    \I__12116\ : InMux
    port map (
            O => \N__49149\,
            I => \N__49146\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__49146\,
            I => \N__49143\
        );

    \I__12114\ : Span4Mux_v
    port map (
            O => \N__49143\,
            I => \N__49140\
        );

    \I__12113\ : Span4Mux_h
    port map (
            O => \N__49140\,
            I => \N__49137\
        );

    \I__12112\ : Span4Mux_v
    port map (
            O => \N__49137\,
            I => \N__49134\
        );

    \I__12111\ : Odrv4
    port map (
            O => \N__49134\,
            I => \c0.n18067\
        );

    \I__12110\ : CascadeMux
    port map (
            O => \N__49131\,
            I => \c0.n18771_cascade_\
        );

    \I__12109\ : InMux
    port map (
            O => \N__49128\,
            I => \N__49125\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__49125\,
            I => \N__49122\
        );

    \I__12107\ : Span4Mux_h
    port map (
            O => \N__49122\,
            I => \N__49119\
        );

    \I__12106\ : Odrv4
    port map (
            O => \N__49119\,
            I => \c0.n18068\
        );

    \I__12105\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49100\
        );

    \I__12104\ : InMux
    port map (
            O => \N__49115\,
            I => \N__49100\
        );

    \I__12103\ : InMux
    port map (
            O => \N__49114\,
            I => \N__49100\
        );

    \I__12102\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49087\
        );

    \I__12101\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49087\
        );

    \I__12100\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49087\
        );

    \I__12099\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49080\
        );

    \I__12098\ : InMux
    port map (
            O => \N__49109\,
            I => \N__49080\
        );

    \I__12097\ : InMux
    port map (
            O => \N__49108\,
            I => \N__49080\
        );

    \I__12096\ : InMux
    port map (
            O => \N__49107\,
            I => \N__49077\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__49100\,
            I => \N__49071\
        );

    \I__12094\ : InMux
    port map (
            O => \N__49099\,
            I => \N__49064\
        );

    \I__12093\ : InMux
    port map (
            O => \N__49098\,
            I => \N__49064\
        );

    \I__12092\ : InMux
    port map (
            O => \N__49097\,
            I => \N__49064\
        );

    \I__12091\ : InMux
    port map (
            O => \N__49096\,
            I => \N__49057\
        );

    \I__12090\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49057\
        );

    \I__12089\ : InMux
    port map (
            O => \N__49094\,
            I => \N__49057\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__49087\,
            I => \N__49054\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__49080\,
            I => \N__49051\
        );

    \I__12086\ : LocalMux
    port map (
            O => \N__49077\,
            I => \N__49042\
        );

    \I__12085\ : InMux
    port map (
            O => \N__49076\,
            I => \N__49035\
        );

    \I__12084\ : InMux
    port map (
            O => \N__49075\,
            I => \N__49035\
        );

    \I__12083\ : InMux
    port map (
            O => \N__49074\,
            I => \N__49035\
        );

    \I__12082\ : Span4Mux_h
    port map (
            O => \N__49071\,
            I => \N__49028\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__49064\,
            I => \N__49028\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__49057\,
            I => \N__49028\
        );

    \I__12079\ : Span4Mux_v
    port map (
            O => \N__49054\,
            I => \N__49022\
        );

    \I__12078\ : Span4Mux_s2_v
    port map (
            O => \N__49051\,
            I => \N__49022\
        );

    \I__12077\ : InMux
    port map (
            O => \N__49050\,
            I => \N__49015\
        );

    \I__12076\ : InMux
    port map (
            O => \N__49049\,
            I => \N__49015\
        );

    \I__12075\ : InMux
    port map (
            O => \N__49048\,
            I => \N__49015\
        );

    \I__12074\ : InMux
    port map (
            O => \N__49047\,
            I => \N__49008\
        );

    \I__12073\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49008\
        );

    \I__12072\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49008\
        );

    \I__12071\ : Span4Mux_v
    port map (
            O => \N__49042\,
            I => \N__49005\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__49035\,
            I => \N__49002\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__49028\,
            I => \N__48999\
        );

    \I__12068\ : InMux
    port map (
            O => \N__49027\,
            I => \N__48995\
        );

    \I__12067\ : Span4Mux_h
    port map (
            O => \N__49022\,
            I => \N__48992\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__49015\,
            I => \N__48987\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__48987\
        );

    \I__12064\ : Span4Mux_h
    port map (
            O => \N__49005\,
            I => \N__48979\
        );

    \I__12063\ : Span4Mux_s3_v
    port map (
            O => \N__49002\,
            I => \N__48979\
        );

    \I__12062\ : Span4Mux_h
    port map (
            O => \N__48999\,
            I => \N__48979\
        );

    \I__12061\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48976\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__48995\,
            I => \N__48969\
        );

    \I__12059\ : Span4Mux_h
    port map (
            O => \N__48992\,
            I => \N__48969\
        );

    \I__12058\ : Span4Mux_s2_v
    port map (
            O => \N__48987\,
            I => \N__48969\
        );

    \I__12057\ : InMux
    port map (
            O => \N__48986\,
            I => \N__48966\
        );

    \I__12056\ : Span4Mux_h
    port map (
            O => \N__48979\,
            I => \N__48961\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__48976\,
            I => \N__48961\
        );

    \I__12054\ : Odrv4
    port map (
            O => \N__48969\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__48966\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12052\ : Odrv4
    port map (
            O => \N__48961\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__12051\ : CascadeMux
    port map (
            O => \N__48954\,
            I => \c0.n18774_cascade_\
        );

    \I__12050\ : InMux
    port map (
            O => \N__48951\,
            I => \N__48944\
        );

    \I__12049\ : InMux
    port map (
            O => \N__48950\,
            I => \N__48941\
        );

    \I__12048\ : InMux
    port map (
            O => \N__48949\,
            I => \N__48938\
        );

    \I__12047\ : InMux
    port map (
            O => \N__48948\,
            I => \N__48935\
        );

    \I__12046\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48932\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__48944\,
            I => \N__48929\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__48941\,
            I => \N__48918\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__48938\,
            I => \N__48918\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__48935\,
            I => \N__48913\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__48932\,
            I => \N__48913\
        );

    \I__12040\ : Span4Mux_s1_v
    port map (
            O => \N__48929\,
            I => \N__48910\
        );

    \I__12039\ : InMux
    port map (
            O => \N__48928\,
            I => \N__48907\
        );

    \I__12038\ : InMux
    port map (
            O => \N__48927\,
            I => \N__48904\
        );

    \I__12037\ : InMux
    port map (
            O => \N__48926\,
            I => \N__48901\
        );

    \I__12036\ : InMux
    port map (
            O => \N__48925\,
            I => \N__48898\
        );

    \I__12035\ : InMux
    port map (
            O => \N__48924\,
            I => \N__48895\
        );

    \I__12034\ : InMux
    port map (
            O => \N__48923\,
            I => \N__48892\
        );

    \I__12033\ : Span4Mux_v
    port map (
            O => \N__48918\,
            I => \N__48888\
        );

    \I__12032\ : Span4Mux_v
    port map (
            O => \N__48913\,
            I => \N__48883\
        );

    \I__12031\ : Span4Mux_v
    port map (
            O => \N__48910\,
            I => \N__48883\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__48907\,
            I => \N__48880\
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__48904\,
            I => \N__48875\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__48901\,
            I => \N__48875\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__48898\,
            I => \N__48872\
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__48895\,
            I => \N__48867\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__48892\,
            I => \N__48867\
        );

    \I__12024\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48864\
        );

    \I__12023\ : Sp12to4
    port map (
            O => \N__48888\,
            I => \N__48857\
        );

    \I__12022\ : Sp12to4
    port map (
            O => \N__48883\,
            I => \N__48857\
        );

    \I__12021\ : Span12Mux_s5_h
    port map (
            O => \N__48880\,
            I => \N__48857\
        );

    \I__12020\ : Span4Mux_s2_v
    port map (
            O => \N__48875\,
            I => \N__48852\
        );

    \I__12019\ : Span4Mux_h
    port map (
            O => \N__48872\,
            I => \N__48852\
        );

    \I__12018\ : Span4Mux_h
    port map (
            O => \N__48867\,
            I => \N__48849\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__48864\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12016\ : Odrv12
    port map (
            O => \N__48857\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12015\ : Odrv4
    port map (
            O => \N__48852\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12014\ : Odrv4
    port map (
            O => \N__48849\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__12013\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48837\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__48837\,
            I => \N__48834\
        );

    \I__12011\ : Span12Mux_s6_h
    port map (
            O => \N__48834\,
            I => \N__48831\
        );

    \I__12010\ : Odrv12
    port map (
            O => \N__48831\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__12009\ : CEMux
    port map (
            O => \N__48828\,
            I => \N__48825\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__48825\,
            I => \N__48820\
        );

    \I__12007\ : CEMux
    port map (
            O => \N__48824\,
            I => \N__48817\
        );

    \I__12006\ : CEMux
    port map (
            O => \N__48823\,
            I => \N__48813\
        );

    \I__12005\ : Span4Mux_v
    port map (
            O => \N__48820\,
            I => \N__48806\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__48817\,
            I => \N__48806\
        );

    \I__12003\ : CEMux
    port map (
            O => \N__48816\,
            I => \N__48803\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__48813\,
            I => \N__48800\
        );

    \I__12001\ : CEMux
    port map (
            O => \N__48812\,
            I => \N__48797\
        );

    \I__12000\ : CEMux
    port map (
            O => \N__48811\,
            I => \N__48793\
        );

    \I__11999\ : Span4Mux_v
    port map (
            O => \N__48806\,
            I => \N__48790\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__48803\,
            I => \N__48787\
        );

    \I__11997\ : Span4Mux_v
    port map (
            O => \N__48800\,
            I => \N__48783\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__48797\,
            I => \N__48780\
        );

    \I__11995\ : CEMux
    port map (
            O => \N__48796\,
            I => \N__48777\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__48793\,
            I => \N__48774\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__48790\,
            I => \N__48771\
        );

    \I__11992\ : Span4Mux_v
    port map (
            O => \N__48787\,
            I => \N__48768\
        );

    \I__11991\ : CEMux
    port map (
            O => \N__48786\,
            I => \N__48765\
        );

    \I__11990\ : Span4Mux_h
    port map (
            O => \N__48783\,
            I => \N__48762\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__48780\,
            I => \N__48757\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__48777\,
            I => \N__48757\
        );

    \I__11987\ : Span4Mux_h
    port map (
            O => \N__48774\,
            I => \N__48754\
        );

    \I__11986\ : Span4Mux_h
    port map (
            O => \N__48771\,
            I => \N__48751\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__48768\,
            I => \N__48748\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__48765\,
            I => \N__48745\
        );

    \I__11983\ : Span4Mux_h
    port map (
            O => \N__48762\,
            I => \N__48742\
        );

    \I__11982\ : Span4Mux_h
    port map (
            O => \N__48757\,
            I => \N__48737\
        );

    \I__11981\ : Span4Mux_h
    port map (
            O => \N__48754\,
            I => \N__48737\
        );

    \I__11980\ : Span4Mux_v
    port map (
            O => \N__48751\,
            I => \N__48734\
        );

    \I__11979\ : Span4Mux_h
    port map (
            O => \N__48748\,
            I => \N__48731\
        );

    \I__11978\ : Span4Mux_h
    port map (
            O => \N__48745\,
            I => \N__48726\
        );

    \I__11977\ : Span4Mux_v
    port map (
            O => \N__48742\,
            I => \N__48726\
        );

    \I__11976\ : Odrv4
    port map (
            O => \N__48737\,
            I => \c0.tx2.n9639\
        );

    \I__11975\ : Odrv4
    port map (
            O => \N__48734\,
            I => \c0.tx2.n9639\
        );

    \I__11974\ : Odrv4
    port map (
            O => \N__48731\,
            I => \c0.tx2.n9639\
        );

    \I__11973\ : Odrv4
    port map (
            O => \N__48726\,
            I => \c0.tx2.n9639\
        );

    \I__11972\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48714\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__48714\,
            I => \N__48711\
        );

    \I__11970\ : Span4Mux_v
    port map (
            O => \N__48711\,
            I => \N__48708\
        );

    \I__11969\ : Odrv4
    port map (
            O => \N__48708\,
            I => \c0.n18669\
        );

    \I__11968\ : InMux
    port map (
            O => \N__48705\,
            I => \N__48697\
        );

    \I__11967\ : CascadeMux
    port map (
            O => \N__48704\,
            I => \N__48675\
        );

    \I__11966\ : CascadeMux
    port map (
            O => \N__48703\,
            I => \N__48672\
        );

    \I__11965\ : CascadeMux
    port map (
            O => \N__48702\,
            I => \N__48669\
        );

    \I__11964\ : CascadeMux
    port map (
            O => \N__48701\,
            I => \N__48666\
        );

    \I__11963\ : CascadeMux
    port map (
            O => \N__48700\,
            I => \N__48663\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__48697\,
            I => \N__48660\
        );

    \I__11961\ : InMux
    port map (
            O => \N__48696\,
            I => \N__48653\
        );

    \I__11960\ : InMux
    port map (
            O => \N__48695\,
            I => \N__48653\
        );

    \I__11959\ : InMux
    port map (
            O => \N__48694\,
            I => \N__48653\
        );

    \I__11958\ : CascadeMux
    port map (
            O => \N__48693\,
            I => \N__48650\
        );

    \I__11957\ : InMux
    port map (
            O => \N__48692\,
            I => \N__48645\
        );

    \I__11956\ : CascadeMux
    port map (
            O => \N__48691\,
            I => \N__48642\
        );

    \I__11955\ : InMux
    port map (
            O => \N__48690\,
            I => \N__48639\
        );

    \I__11954\ : CascadeMux
    port map (
            O => \N__48689\,
            I => \N__48632\
        );

    \I__11953\ : CascadeMux
    port map (
            O => \N__48688\,
            I => \N__48628\
        );

    \I__11952\ : CascadeMux
    port map (
            O => \N__48687\,
            I => \N__48625\
        );

    \I__11951\ : InMux
    port map (
            O => \N__48686\,
            I => \N__48613\
        );

    \I__11950\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48613\
        );

    \I__11949\ : CascadeMux
    port map (
            O => \N__48684\,
            I => \N__48610\
        );

    \I__11948\ : CascadeMux
    port map (
            O => \N__48683\,
            I => \N__48599\
        );

    \I__11947\ : CascadeMux
    port map (
            O => \N__48682\,
            I => \N__48596\
        );

    \I__11946\ : CascadeMux
    port map (
            O => \N__48681\,
            I => \N__48592\
        );

    \I__11945\ : InMux
    port map (
            O => \N__48680\,
            I => \N__48586\
        );

    \I__11944\ : InMux
    port map (
            O => \N__48679\,
            I => \N__48586\
        );

    \I__11943\ : InMux
    port map (
            O => \N__48678\,
            I => \N__48579\
        );

    \I__11942\ : InMux
    port map (
            O => \N__48675\,
            I => \N__48579\
        );

    \I__11941\ : InMux
    port map (
            O => \N__48672\,
            I => \N__48579\
        );

    \I__11940\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48574\
        );

    \I__11939\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48574\
        );

    \I__11938\ : InMux
    port map (
            O => \N__48663\,
            I => \N__48571\
        );

    \I__11937\ : Span4Mux_v
    port map (
            O => \N__48660\,
            I => \N__48565\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__48653\,
            I => \N__48565\
        );

    \I__11935\ : InMux
    port map (
            O => \N__48650\,
            I => \N__48562\
        );

    \I__11934\ : CascadeMux
    port map (
            O => \N__48649\,
            I => \N__48559\
        );

    \I__11933\ : CascadeMux
    port map (
            O => \N__48648\,
            I => \N__48553\
        );

    \I__11932\ : LocalMux
    port map (
            O => \N__48645\,
            I => \N__48550\
        );

    \I__11931\ : InMux
    port map (
            O => \N__48642\,
            I => \N__48547\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__48639\,
            I => \N__48544\
        );

    \I__11929\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48539\
        );

    \I__11928\ : InMux
    port map (
            O => \N__48637\,
            I => \N__48539\
        );

    \I__11927\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48532\
        );

    \I__11926\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48532\
        );

    \I__11925\ : InMux
    port map (
            O => \N__48632\,
            I => \N__48532\
        );

    \I__11924\ : InMux
    port map (
            O => \N__48631\,
            I => \N__48525\
        );

    \I__11923\ : InMux
    port map (
            O => \N__48628\,
            I => \N__48525\
        );

    \I__11922\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48525\
        );

    \I__11921\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48521\
        );

    \I__11920\ : InMux
    port map (
            O => \N__48623\,
            I => \N__48518\
        );

    \I__11919\ : InMux
    port map (
            O => \N__48622\,
            I => \N__48515\
        );

    \I__11918\ : InMux
    port map (
            O => \N__48621\,
            I => \N__48510\
        );

    \I__11917\ : InMux
    port map (
            O => \N__48620\,
            I => \N__48510\
        );

    \I__11916\ : InMux
    port map (
            O => \N__48619\,
            I => \N__48505\
        );

    \I__11915\ : InMux
    port map (
            O => \N__48618\,
            I => \N__48505\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__48613\,
            I => \N__48502\
        );

    \I__11913\ : InMux
    port map (
            O => \N__48610\,
            I => \N__48497\
        );

    \I__11912\ : InMux
    port map (
            O => \N__48609\,
            I => \N__48497\
        );

    \I__11911\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48492\
        );

    \I__11910\ : InMux
    port map (
            O => \N__48607\,
            I => \N__48492\
        );

    \I__11909\ : CascadeMux
    port map (
            O => \N__48606\,
            I => \N__48484\
        );

    \I__11908\ : InMux
    port map (
            O => \N__48605\,
            I => \N__48475\
        );

    \I__11907\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48475\
        );

    \I__11906\ : InMux
    port map (
            O => \N__48603\,
            I => \N__48470\
        );

    \I__11905\ : InMux
    port map (
            O => \N__48602\,
            I => \N__48470\
        );

    \I__11904\ : InMux
    port map (
            O => \N__48599\,
            I => \N__48459\
        );

    \I__11903\ : InMux
    port map (
            O => \N__48596\,
            I => \N__48459\
        );

    \I__11902\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48459\
        );

    \I__11901\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48459\
        );

    \I__11900\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48459\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__48586\,
            I => \N__48454\
        );

    \I__11898\ : LocalMux
    port map (
            O => \N__48579\,
            I => \N__48454\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__48574\,
            I => \N__48449\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__48571\,
            I => \N__48449\
        );

    \I__11895\ : CascadeMux
    port map (
            O => \N__48570\,
            I => \N__48446\
        );

    \I__11894\ : Span4Mux_v
    port map (
            O => \N__48565\,
            I => \N__48441\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__48562\,
            I => \N__48441\
        );

    \I__11892\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48438\
        );

    \I__11891\ : InMux
    port map (
            O => \N__48558\,
            I => \N__48429\
        );

    \I__11890\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48429\
        );

    \I__11889\ : InMux
    port map (
            O => \N__48556\,
            I => \N__48429\
        );

    \I__11888\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48429\
        );

    \I__11887\ : Span4Mux_v
    port map (
            O => \N__48550\,
            I => \N__48424\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__48547\,
            I => \N__48424\
        );

    \I__11885\ : Span4Mux_v
    port map (
            O => \N__48544\,
            I => \N__48415\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__48539\,
            I => \N__48415\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__48532\,
            I => \N__48415\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__48525\,
            I => \N__48415\
        );

    \I__11881\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48412\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__48521\,
            I => \N__48407\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__48518\,
            I => \N__48407\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__48515\,
            I => \N__48404\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48399\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__48505\,
            I => \N__48390\
        );

    \I__11875\ : Span4Mux_s3_v
    port map (
            O => \N__48502\,
            I => \N__48390\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48390\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__48492\,
            I => \N__48390\
        );

    \I__11872\ : CascadeMux
    port map (
            O => \N__48491\,
            I => \N__48386\
        );

    \I__11871\ : CascadeMux
    port map (
            O => \N__48490\,
            I => \N__48383\
        );

    \I__11870\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48378\
        );

    \I__11869\ : InMux
    port map (
            O => \N__48488\,
            I => \N__48378\
        );

    \I__11868\ : InMux
    port map (
            O => \N__48487\,
            I => \N__48373\
        );

    \I__11867\ : InMux
    port map (
            O => \N__48484\,
            I => \N__48373\
        );

    \I__11866\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48367\
        );

    \I__11865\ : InMux
    port map (
            O => \N__48482\,
            I => \N__48367\
        );

    \I__11864\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48362\
        );

    \I__11863\ : InMux
    port map (
            O => \N__48480\,
            I => \N__48362\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__48475\,
            I => \N__48355\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__48470\,
            I => \N__48355\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__48459\,
            I => \N__48355\
        );

    \I__11859\ : Span4Mux_h
    port map (
            O => \N__48454\,
            I => \N__48352\
        );

    \I__11858\ : Span4Mux_h
    port map (
            O => \N__48449\,
            I => \N__48349\
        );

    \I__11857\ : InMux
    port map (
            O => \N__48446\,
            I => \N__48346\
        );

    \I__11856\ : Span4Mux_h
    port map (
            O => \N__48441\,
            I => \N__48343\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__48438\,
            I => \N__48332\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__48429\,
            I => \N__48332\
        );

    \I__11853\ : Span4Mux_h
    port map (
            O => \N__48424\,
            I => \N__48332\
        );

    \I__11852\ : Span4Mux_v
    port map (
            O => \N__48415\,
            I => \N__48332\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__48412\,
            I => \N__48332\
        );

    \I__11850\ : Span4Mux_s3_v
    port map (
            O => \N__48407\,
            I => \N__48329\
        );

    \I__11849\ : Span4Mux_s3_v
    port map (
            O => \N__48404\,
            I => \N__48326\
        );

    \I__11848\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48321\
        );

    \I__11847\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48321\
        );

    \I__11846\ : Span4Mux_v
    port map (
            O => \N__48399\,
            I => \N__48316\
        );

    \I__11845\ : Span4Mux_v
    port map (
            O => \N__48390\,
            I => \N__48316\
        );

    \I__11844\ : InMux
    port map (
            O => \N__48389\,
            I => \N__48311\
        );

    \I__11843\ : InMux
    port map (
            O => \N__48386\,
            I => \N__48311\
        );

    \I__11842\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48308\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48303\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48303\
        );

    \I__11839\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48300\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48295\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__48362\,
            I => \N__48295\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__48355\,
            I => \N__48292\
        );

    \I__11835\ : Span4Mux_v
    port map (
            O => \N__48352\,
            I => \N__48287\
        );

    \I__11834\ : Span4Mux_v
    port map (
            O => \N__48349\,
            I => \N__48287\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__48346\,
            I => \N__48283\
        );

    \I__11832\ : Span4Mux_h
    port map (
            O => \N__48343\,
            I => \N__48278\
        );

    \I__11831\ : Span4Mux_h
    port map (
            O => \N__48332\,
            I => \N__48278\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__48329\,
            I => \N__48273\
        );

    \I__11829\ : Span4Mux_v
    port map (
            O => \N__48326\,
            I => \N__48273\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__48321\,
            I => \N__48266\
        );

    \I__11827\ : Sp12to4
    port map (
            O => \N__48316\,
            I => \N__48266\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__48311\,
            I => \N__48266\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__48308\,
            I => \N__48259\
        );

    \I__11824\ : Sp12to4
    port map (
            O => \N__48303\,
            I => \N__48259\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__48300\,
            I => \N__48259\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__48295\,
            I => \N__48252\
        );

    \I__11821\ : Span4Mux_v
    port map (
            O => \N__48292\,
            I => \N__48252\
        );

    \I__11820\ : Span4Mux_h
    port map (
            O => \N__48287\,
            I => \N__48252\
        );

    \I__11819\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48249\
        );

    \I__11818\ : Span4Mux_h
    port map (
            O => \N__48283\,
            I => \N__48246\
        );

    \I__11817\ : Span4Mux_h
    port map (
            O => \N__48278\,
            I => \N__48243\
        );

    \I__11816\ : Sp12to4
    port map (
            O => \N__48273\,
            I => \N__48236\
        );

    \I__11815\ : Span12Mux_h
    port map (
            O => \N__48266\,
            I => \N__48236\
        );

    \I__11814\ : Span12Mux_s7_v
    port map (
            O => \N__48259\,
            I => \N__48236\
        );

    \I__11813\ : Span4Mux_h
    port map (
            O => \N__48252\,
            I => \N__48233\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__48249\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11811\ : Odrv4
    port map (
            O => \N__48246\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11810\ : Odrv4
    port map (
            O => \N__48243\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11809\ : Odrv12
    port map (
            O => \N__48236\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11808\ : Odrv4
    port map (
            O => \N__48233\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__11807\ : InMux
    port map (
            O => \N__48222\,
            I => \N__48216\
        );

    \I__11806\ : InMux
    port map (
            O => \N__48221\,
            I => \N__48213\
        );

    \I__11805\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48210\
        );

    \I__11804\ : InMux
    port map (
            O => \N__48219\,
            I => \N__48207\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__48216\,
            I => \N__48204\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__48213\,
            I => \N__48201\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__48210\,
            I => \N__48198\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__48207\,
            I => \N__48193\
        );

    \I__11799\ : Span4Mux_v
    port map (
            O => \N__48204\,
            I => \N__48193\
        );

    \I__11798\ : Span4Mux_h
    port map (
            O => \N__48201\,
            I => \N__48190\
        );

    \I__11797\ : Span4Mux_s1_v
    port map (
            O => \N__48198\,
            I => \N__48187\
        );

    \I__11796\ : Odrv4
    port map (
            O => \N__48193\,
            I => data_out_frame2_16_4
        );

    \I__11795\ : Odrv4
    port map (
            O => \N__48190\,
            I => data_out_frame2_16_4
        );

    \I__11794\ : Odrv4
    port map (
            O => \N__48187\,
            I => data_out_frame2_16_4
        );

    \I__11793\ : InMux
    port map (
            O => \N__48180\,
            I => \N__48177\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__48177\,
            I => \N__48174\
        );

    \I__11791\ : Odrv12
    port map (
            O => \N__48174\,
            I => \c0.data_out_frame2_20_4\
        );

    \I__11790\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48165\
        );

    \I__11789\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48162\
        );

    \I__11788\ : InMux
    port map (
            O => \N__48169\,
            I => \N__48158\
        );

    \I__11787\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48154\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__48165\,
            I => \N__48149\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__48162\,
            I => \N__48149\
        );

    \I__11784\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48146\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__48158\,
            I => \N__48143\
        );

    \I__11782\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48140\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48135\
        );

    \I__11780\ : Span4Mux_h
    port map (
            O => \N__48149\,
            I => \N__48130\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__48146\,
            I => \N__48130\
        );

    \I__11778\ : Span4Mux_s2_v
    port map (
            O => \N__48143\,
            I => \N__48127\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48124\
        );

    \I__11776\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48121\
        );

    \I__11775\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48118\
        );

    \I__11774\ : Span4Mux_s3_v
    port map (
            O => \N__48135\,
            I => \N__48115\
        );

    \I__11773\ : Sp12to4
    port map (
            O => \N__48130\,
            I => \N__48112\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__48127\,
            I => \N__48105\
        );

    \I__11771\ : Span4Mux_v
    port map (
            O => \N__48124\,
            I => \N__48105\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__48121\,
            I => \N__48105\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48102\
        );

    \I__11768\ : Span4Mux_h
    port map (
            O => \N__48115\,
            I => \N__48099\
        );

    \I__11767\ : Span12Mux_s7_v
    port map (
            O => \N__48112\,
            I => \N__48096\
        );

    \I__11766\ : Span4Mux_h
    port map (
            O => \N__48105\,
            I => \N__48093\
        );

    \I__11765\ : Odrv4
    port map (
            O => \N__48102\,
            I => \c0.n7263\
        );

    \I__11764\ : Odrv4
    port map (
            O => \N__48099\,
            I => \c0.n7263\
        );

    \I__11763\ : Odrv12
    port map (
            O => \N__48096\,
            I => \c0.n7263\
        );

    \I__11762\ : Odrv4
    port map (
            O => \N__48093\,
            I => \c0.n7263\
        );

    \I__11761\ : CascadeMux
    port map (
            O => \N__48084\,
            I => \c0.n18672_cascade_\
        );

    \I__11760\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48072\
        );

    \I__11759\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48065\
        );

    \I__11758\ : InMux
    port map (
            O => \N__48079\,
            I => \N__48065\
        );

    \I__11757\ : InMux
    port map (
            O => \N__48078\,
            I => \N__48062\
        );

    \I__11756\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48057\
        );

    \I__11755\ : InMux
    port map (
            O => \N__48076\,
            I => \N__48057\
        );

    \I__11754\ : InMux
    port map (
            O => \N__48075\,
            I => \N__48054\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__48072\,
            I => \N__48051\
        );

    \I__11752\ : InMux
    port map (
            O => \N__48071\,
            I => \N__48046\
        );

    \I__11751\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48046\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__48065\,
            I => \N__48043\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__48062\,
            I => \N__48036\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__48057\,
            I => \N__48036\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__48054\,
            I => \N__48036\
        );

    \I__11746\ : Span4Mux_v
    port map (
            O => \N__48051\,
            I => \N__48026\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__48046\,
            I => \N__48023\
        );

    \I__11744\ : Span4Mux_v
    port map (
            O => \N__48043\,
            I => \N__48018\
        );

    \I__11743\ : Span4Mux_v
    port map (
            O => \N__48036\,
            I => \N__48018\
        );

    \I__11742\ : InMux
    port map (
            O => \N__48035\,
            I => \N__48012\
        );

    \I__11741\ : InMux
    port map (
            O => \N__48034\,
            I => \N__48012\
        );

    \I__11740\ : CascadeMux
    port map (
            O => \N__48033\,
            I => \N__48009\
        );

    \I__11739\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48004\
        );

    \I__11738\ : InMux
    port map (
            O => \N__48031\,
            I => \N__48004\
        );

    \I__11737\ : InMux
    port map (
            O => \N__48030\,
            I => \N__47999\
        );

    \I__11736\ : InMux
    port map (
            O => \N__48029\,
            I => \N__47999\
        );

    \I__11735\ : Span4Mux_v
    port map (
            O => \N__48026\,
            I => \N__47994\
        );

    \I__11734\ : Span4Mux_s1_v
    port map (
            O => \N__48023\,
            I => \N__47994\
        );

    \I__11733\ : Span4Mux_h
    port map (
            O => \N__48018\,
            I => \N__47991\
        );

    \I__11732\ : InMux
    port map (
            O => \N__48017\,
            I => \N__47988\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__48012\,
            I => \N__47985\
        );

    \I__11730\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47982\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__48004\,
            I => \N__47978\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__47999\,
            I => \N__47972\
        );

    \I__11727\ : Span4Mux_h
    port map (
            O => \N__47994\,
            I => \N__47972\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__47991\,
            I => \N__47969\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__47988\,
            I => \N__47966\
        );

    \I__11724\ : Span4Mux_s2_v
    port map (
            O => \N__47985\,
            I => \N__47961\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__47982\,
            I => \N__47961\
        );

    \I__11722\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47957\
        );

    \I__11721\ : Span4Mux_s1_v
    port map (
            O => \N__47978\,
            I => \N__47954\
        );

    \I__11720\ : InMux
    port map (
            O => \N__47977\,
            I => \N__47951\
        );

    \I__11719\ : Span4Mux_h
    port map (
            O => \N__47972\,
            I => \N__47944\
        );

    \I__11718\ : Span4Mux_v
    port map (
            O => \N__47969\,
            I => \N__47944\
        );

    \I__11717\ : Span4Mux_v
    port map (
            O => \N__47966\,
            I => \N__47944\
        );

    \I__11716\ : Span4Mux_h
    port map (
            O => \N__47961\,
            I => \N__47941\
        );

    \I__11715\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47938\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__47957\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11713\ : Odrv4
    port map (
            O => \N__47954\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__47951\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11711\ : Odrv4
    port map (
            O => \N__47944\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11710\ : Odrv4
    port map (
            O => \N__47941\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__47938\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__11708\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47922\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__47922\,
            I => \c0.n22_adj_2243\
        );

    \I__11706\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47916\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__47916\,
            I => \N__47912\
        );

    \I__11704\ : CascadeMux
    port map (
            O => \N__47915\,
            I => \N__47909\
        );

    \I__11703\ : Span4Mux_h
    port map (
            O => \N__47912\,
            I => \N__47906\
        );

    \I__11702\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47903\
        );

    \I__11701\ : Odrv4
    port map (
            O => \N__47906\,
            I => rand_setpoint_14
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__47903\,
            I => rand_setpoint_14
        );

    \I__11699\ : CEMux
    port map (
            O => \N__47898\,
            I => \N__47895\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__47895\,
            I => \N__47890\
        );

    \I__11697\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47887\
        );

    \I__11696\ : CEMux
    port map (
            O => \N__47893\,
            I => \N__47880\
        );

    \I__11695\ : Span4Mux_v
    port map (
            O => \N__47890\,
            I => \N__47875\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__47887\,
            I => \N__47875\
        );

    \I__11693\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47872\
        );

    \I__11692\ : CEMux
    port map (
            O => \N__47885\,
            I => \N__47868\
        );

    \I__11691\ : CEMux
    port map (
            O => \N__47884\,
            I => \N__47865\
        );

    \I__11690\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47862\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47859\
        );

    \I__11688\ : Span4Mux_h
    port map (
            O => \N__47875\,
            I => \N__47854\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__47872\,
            I => \N__47854\
        );

    \I__11686\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47851\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__47868\,
            I => \N__47848\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__47865\,
            I => \N__47845\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__47862\,
            I => \N__47842\
        );

    \I__11682\ : Span4Mux_h
    port map (
            O => \N__47859\,
            I => \N__47839\
        );

    \I__11681\ : Span4Mux_v
    port map (
            O => \N__47854\,
            I => \N__47834\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__47851\,
            I => \N__47834\
        );

    \I__11679\ : Span4Mux_v
    port map (
            O => \N__47848\,
            I => \N__47831\
        );

    \I__11678\ : Span4Mux_h
    port map (
            O => \N__47845\,
            I => \N__47826\
        );

    \I__11677\ : Span4Mux_v
    port map (
            O => \N__47842\,
            I => \N__47826\
        );

    \I__11676\ : Span4Mux_h
    port map (
            O => \N__47839\,
            I => \N__47821\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__47834\,
            I => \N__47821\
        );

    \I__11674\ : Odrv4
    port map (
            O => \N__47831\,
            I => \c0.n11016\
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__47826\,
            I => \c0.n11016\
        );

    \I__11672\ : Odrv4
    port map (
            O => \N__47821\,
            I => \c0.n11016\
        );

    \I__11671\ : CascadeMux
    port map (
            O => \N__47814\,
            I => \N__47811\
        );

    \I__11670\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47806\
        );

    \I__11669\ : CascadeMux
    port map (
            O => \N__47810\,
            I => \N__47803\
        );

    \I__11668\ : CascadeMux
    port map (
            O => \N__47809\,
            I => \N__47800\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47795\
        );

    \I__11666\ : InMux
    port map (
            O => \N__47803\,
            I => \N__47792\
        );

    \I__11665\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47788\
        );

    \I__11664\ : CascadeMux
    port map (
            O => \N__47799\,
            I => \N__47785\
        );

    \I__11663\ : CascadeMux
    port map (
            O => \N__47798\,
            I => \N__47782\
        );

    \I__11662\ : Span4Mux_v
    port map (
            O => \N__47795\,
            I => \N__47777\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47777\
        );

    \I__11660\ : CascadeMux
    port map (
            O => \N__47791\,
            I => \N__47774\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47771\
        );

    \I__11658\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47768\
        );

    \I__11657\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47765\
        );

    \I__11656\ : Span4Mux_h
    port map (
            O => \N__47777\,
            I => \N__47762\
        );

    \I__11655\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47759\
        );

    \I__11654\ : Span4Mux_h
    port map (
            O => \N__47771\,
            I => \N__47754\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__47768\,
            I => \N__47754\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__47765\,
            I => \N__47751\
        );

    \I__11651\ : Span4Mux_v
    port map (
            O => \N__47762\,
            I => \N__47746\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47746\
        );

    \I__11649\ : Span4Mux_v
    port map (
            O => \N__47754\,
            I => \N__47741\
        );

    \I__11648\ : Span4Mux_h
    port map (
            O => \N__47751\,
            I => \N__47741\
        );

    \I__11647\ : Odrv4
    port map (
            O => \N__47746\,
            I => n2732
        );

    \I__11646\ : Odrv4
    port map (
            O => \N__47741\,
            I => n2732
        );

    \I__11645\ : InMux
    port map (
            O => \N__47736\,
            I => \N__47730\
        );

    \I__11644\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47727\
        );

    \I__11643\ : InMux
    port map (
            O => \N__47734\,
            I => \N__47724\
        );

    \I__11642\ : InMux
    port map (
            O => \N__47733\,
            I => \N__47720\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__47730\,
            I => \N__47715\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__47727\,
            I => \N__47715\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47712\
        );

    \I__11638\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47709\
        );

    \I__11637\ : LocalMux
    port map (
            O => \N__47720\,
            I => \N__47706\
        );

    \I__11636\ : Span4Mux_v
    port map (
            O => \N__47715\,
            I => \N__47703\
        );

    \I__11635\ : Span4Mux_h
    port map (
            O => \N__47712\,
            I => \N__47700\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__47709\,
            I => \c0.data_out_7_6\
        );

    \I__11633\ : Odrv12
    port map (
            O => \N__47706\,
            I => \c0.data_out_7_6\
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__47703\,
            I => \c0.data_out_7_6\
        );

    \I__11631\ : Odrv4
    port map (
            O => \N__47700\,
            I => \c0.data_out_7_6\
        );

    \I__11630\ : CascadeMux
    port map (
            O => \N__47691\,
            I => \N__47682\
        );

    \I__11629\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47673\
        );

    \I__11628\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47665\
        );

    \I__11627\ : InMux
    port map (
            O => \N__47688\,
            I => \N__47662\
        );

    \I__11626\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47655\
        );

    \I__11625\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47655\
        );

    \I__11624\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47652\
        );

    \I__11623\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47647\
        );

    \I__11622\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47647\
        );

    \I__11621\ : InMux
    port map (
            O => \N__47680\,
            I => \N__47641\
        );

    \I__11620\ : InMux
    port map (
            O => \N__47679\,
            I => \N__47641\
        );

    \I__11619\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47638\
        );

    \I__11618\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47635\
        );

    \I__11617\ : InMux
    port map (
            O => \N__47676\,
            I => \N__47629\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__47673\,
            I => \N__47626\
        );

    \I__11615\ : CascadeMux
    port map (
            O => \N__47672\,
            I => \N__47622\
        );

    \I__11614\ : InMux
    port map (
            O => \N__47671\,
            I => \N__47619\
        );

    \I__11613\ : CascadeMux
    port map (
            O => \N__47670\,
            I => \N__47616\
        );

    \I__11612\ : CascadeMux
    port map (
            O => \N__47669\,
            I => \N__47611\
        );

    \I__11611\ : InMux
    port map (
            O => \N__47668\,
            I => \N__47607\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__47665\,
            I => \N__47604\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__47662\,
            I => \N__47599\
        );

    \I__11608\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47596\
        );

    \I__11607\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47593\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__47655\,
            I => \N__47590\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__47652\,
            I => \N__47587\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__47647\,
            I => \N__47584\
        );

    \I__11603\ : InMux
    port map (
            O => \N__47646\,
            I => \N__47581\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__47641\,
            I => \N__47578\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__47638\,
            I => \N__47573\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__47635\,
            I => \N__47573\
        );

    \I__11599\ : InMux
    port map (
            O => \N__47634\,
            I => \N__47570\
        );

    \I__11598\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47567\
        );

    \I__11597\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47564\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__47629\,
            I => \N__47561\
        );

    \I__11595\ : Span4Mux_h
    port map (
            O => \N__47626\,
            I => \N__47558\
        );

    \I__11594\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47555\
        );

    \I__11593\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47551\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__47619\,
            I => \N__47546\
        );

    \I__11591\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47543\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__47615\,
            I => \N__47540\
        );

    \I__11589\ : CascadeMux
    port map (
            O => \N__47614\,
            I => \N__47537\
        );

    \I__11588\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47533\
        );

    \I__11587\ : InMux
    port map (
            O => \N__47610\,
            I => \N__47530\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__47607\,
            I => \N__47527\
        );

    \I__11585\ : Span4Mux_v
    port map (
            O => \N__47604\,
            I => \N__47524\
        );

    \I__11584\ : InMux
    port map (
            O => \N__47603\,
            I => \N__47519\
        );

    \I__11583\ : InMux
    port map (
            O => \N__47602\,
            I => \N__47519\
        );

    \I__11582\ : Span4Mux_v
    port map (
            O => \N__47599\,
            I => \N__47512\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__47596\,
            I => \N__47512\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__47593\,
            I => \N__47512\
        );

    \I__11579\ : Span4Mux_v
    port map (
            O => \N__47590\,
            I => \N__47509\
        );

    \I__11578\ : Span4Mux_v
    port map (
            O => \N__47587\,
            I => \N__47506\
        );

    \I__11577\ : Span4Mux_v
    port map (
            O => \N__47584\,
            I => \N__47495\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__47581\,
            I => \N__47495\
        );

    \I__11575\ : Span4Mux_v
    port map (
            O => \N__47578\,
            I => \N__47495\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__47573\,
            I => \N__47495\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__47570\,
            I => \N__47495\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__47567\,
            I => \N__47492\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47483\
        );

    \I__11570\ : Span12Mux_h
    port map (
            O => \N__47561\,
            I => \N__47483\
        );

    \I__11569\ : Sp12to4
    port map (
            O => \N__47558\,
            I => \N__47483\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__47555\,
            I => \N__47483\
        );

    \I__11567\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47480\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__47551\,
            I => \N__47477\
        );

    \I__11565\ : InMux
    port map (
            O => \N__47550\,
            I => \N__47474\
        );

    \I__11564\ : InMux
    port map (
            O => \N__47549\,
            I => \N__47471\
        );

    \I__11563\ : Span4Mux_h
    port map (
            O => \N__47546\,
            I => \N__47466\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__47543\,
            I => \N__47466\
        );

    \I__11561\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47463\
        );

    \I__11560\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47458\
        );

    \I__11559\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47458\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__47533\,
            I => \N__47439\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__47530\,
            I => \N__47439\
        );

    \I__11556\ : Span4Mux_v
    port map (
            O => \N__47527\,
            I => \N__47439\
        );

    \I__11555\ : Span4Mux_h
    port map (
            O => \N__47524\,
            I => \N__47439\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__47519\,
            I => \N__47439\
        );

    \I__11553\ : Span4Mux_v
    port map (
            O => \N__47512\,
            I => \N__47439\
        );

    \I__11552\ : Span4Mux_h
    port map (
            O => \N__47509\,
            I => \N__47439\
        );

    \I__11551\ : Span4Mux_h
    port map (
            O => \N__47506\,
            I => \N__47439\
        );

    \I__11550\ : Span4Mux_v
    port map (
            O => \N__47495\,
            I => \N__47439\
        );

    \I__11549\ : Span12Mux_v
    port map (
            O => \N__47492\,
            I => \N__47436\
        );

    \I__11548\ : Span12Mux_v
    port map (
            O => \N__47483\,
            I => \N__47433\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__47480\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11546\ : Odrv4
    port map (
            O => \N__47477\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__47474\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__47471\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11543\ : Odrv4
    port map (
            O => \N__47466\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__47463\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__47458\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11540\ : Odrv4
    port map (
            O => \N__47439\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11539\ : Odrv12
    port map (
            O => \N__47436\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11538\ : Odrv12
    port map (
            O => \N__47433\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11537\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47395\
        );

    \I__11536\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47391\
        );

    \I__11535\ : InMux
    port map (
            O => \N__47410\,
            I => \N__47388\
        );

    \I__11534\ : InMux
    port map (
            O => \N__47409\,
            I => \N__47381\
        );

    \I__11533\ : InMux
    port map (
            O => \N__47408\,
            I => \N__47381\
        );

    \I__11532\ : InMux
    port map (
            O => \N__47407\,
            I => \N__47381\
        );

    \I__11531\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47375\
        );

    \I__11530\ : InMux
    port map (
            O => \N__47405\,
            I => \N__47375\
        );

    \I__11529\ : InMux
    port map (
            O => \N__47404\,
            I => \N__47372\
        );

    \I__11528\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47369\
        );

    \I__11527\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47366\
        );

    \I__11526\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47362\
        );

    \I__11525\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47359\
        );

    \I__11524\ : InMux
    port map (
            O => \N__47399\,
            I => \N__47350\
        );

    \I__11523\ : InMux
    port map (
            O => \N__47398\,
            I => \N__47347\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__47395\,
            I => \N__47342\
        );

    \I__11521\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47339\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__47391\,
            I => \N__47332\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__47388\,
            I => \N__47332\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__47381\,
            I => \N__47332\
        );

    \I__11517\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47329\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__47375\,
            I => \N__47324\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__47372\,
            I => \N__47324\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__47369\,
            I => \N__47321\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__47366\,
            I => \N__47317\
        );

    \I__11512\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47314\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__47362\,
            I => \N__47308\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__47359\,
            I => \N__47308\
        );

    \I__11509\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47299\
        );

    \I__11508\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47299\
        );

    \I__11507\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47299\
        );

    \I__11506\ : InMux
    port map (
            O => \N__47355\,
            I => \N__47299\
        );

    \I__11505\ : InMux
    port map (
            O => \N__47354\,
            I => \N__47294\
        );

    \I__11504\ : InMux
    port map (
            O => \N__47353\,
            I => \N__47294\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__47350\,
            I => \N__47288\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__47347\,
            I => \N__47285\
        );

    \I__11501\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47282\
        );

    \I__11500\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47279\
        );

    \I__11499\ : Span4Mux_v
    port map (
            O => \N__47342\,
            I => \N__47276\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__47339\,
            I => \N__47273\
        );

    \I__11497\ : Span4Mux_v
    port map (
            O => \N__47332\,
            I => \N__47264\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__47329\,
            I => \N__47264\
        );

    \I__11495\ : Span4Mux_v
    port map (
            O => \N__47324\,
            I => \N__47264\
        );

    \I__11494\ : Span4Mux_h
    port map (
            O => \N__47321\,
            I => \N__47264\
        );

    \I__11493\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47261\
        );

    \I__11492\ : Span4Mux_v
    port map (
            O => \N__47317\,
            I => \N__47249\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__47314\,
            I => \N__47249\
        );

    \I__11490\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47246\
        );

    \I__11489\ : Span4Mux_v
    port map (
            O => \N__47308\,
            I => \N__47243\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__47299\,
            I => \N__47238\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__47294\,
            I => \N__47238\
        );

    \I__11486\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47229\
        );

    \I__11485\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47229\
        );

    \I__11484\ : InMux
    port map (
            O => \N__47291\,
            I => \N__47229\
        );

    \I__11483\ : Span4Mux_h
    port map (
            O => \N__47288\,
            I => \N__47225\
        );

    \I__11482\ : Span4Mux_h
    port map (
            O => \N__47285\,
            I => \N__47210\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__47282\,
            I => \N__47210\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__47279\,
            I => \N__47210\
        );

    \I__11479\ : Span4Mux_h
    port map (
            O => \N__47276\,
            I => \N__47210\
        );

    \I__11478\ : Span4Mux_h
    port map (
            O => \N__47273\,
            I => \N__47210\
        );

    \I__11477\ : Span4Mux_h
    port map (
            O => \N__47264\,
            I => \N__47210\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__47261\,
            I => \N__47210\
        );

    \I__11475\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47205\
        );

    \I__11474\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47205\
        );

    \I__11473\ : InMux
    port map (
            O => \N__47258\,
            I => \N__47202\
        );

    \I__11472\ : InMux
    port map (
            O => \N__47257\,
            I => \N__47197\
        );

    \I__11471\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47197\
        );

    \I__11470\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47192\
        );

    \I__11469\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47192\
        );

    \I__11468\ : Span4Mux_v
    port map (
            O => \N__47249\,
            I => \N__47183\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__47246\,
            I => \N__47183\
        );

    \I__11466\ : Span4Mux_v
    port map (
            O => \N__47243\,
            I => \N__47183\
        );

    \I__11465\ : Span4Mux_v
    port map (
            O => \N__47238\,
            I => \N__47183\
        );

    \I__11464\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47178\
        );

    \I__11463\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47178\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47175\
        );

    \I__11461\ : InMux
    port map (
            O => \N__47228\,
            I => \N__47172\
        );

    \I__11460\ : Span4Mux_h
    port map (
            O => \N__47225\,
            I => \N__47167\
        );

    \I__11459\ : Span4Mux_v
    port map (
            O => \N__47210\,
            I => \N__47167\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__47205\,
            I => \N__47162\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__47202\,
            I => \N__47162\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__47197\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__47192\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11454\ : Odrv4
    port map (
            O => \N__47183\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__47178\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11452\ : Odrv12
    port map (
            O => \N__47175\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__47172\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11450\ : Odrv4
    port map (
            O => \N__47167\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11449\ : Odrv4
    port map (
            O => \N__47162\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11448\ : InMux
    port map (
            O => \N__47145\,
            I => \N__47134\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47131\
        );

    \I__11446\ : InMux
    port map (
            O => \N__47143\,
            I => \N__47124\
        );

    \I__11445\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47112\
        );

    \I__11444\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47108\
        );

    \I__11443\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47105\
        );

    \I__11442\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47102\
        );

    \I__11441\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47097\
        );

    \I__11440\ : InMux
    port map (
            O => \N__47137\,
            I => \N__47097\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__47134\,
            I => \N__47092\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__47131\,
            I => \N__47092\
        );

    \I__11437\ : InMux
    port map (
            O => \N__47130\,
            I => \N__47089\
        );

    \I__11436\ : InMux
    port map (
            O => \N__47129\,
            I => \N__47086\
        );

    \I__11435\ : CascadeMux
    port map (
            O => \N__47128\,
            I => \N__47082\
        );

    \I__11434\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47077\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__47124\,
            I => \N__47074\
        );

    \I__11432\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47067\
        );

    \I__11431\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47060\
        );

    \I__11430\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47055\
        );

    \I__11429\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47050\
        );

    \I__11428\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47050\
        );

    \I__11427\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47047\
        );

    \I__11426\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47040\
        );

    \I__11425\ : InMux
    port map (
            O => \N__47116\,
            I => \N__47040\
        );

    \I__11424\ : InMux
    port map (
            O => \N__47115\,
            I => \N__47040\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47037\
        );

    \I__11422\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47034\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__47108\,
            I => \N__47027\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__47105\,
            I => \N__47027\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__47027\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__47097\,
            I => \N__47024\
        );

    \I__11417\ : Span4Mux_v
    port map (
            O => \N__47092\,
            I => \N__47019\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47019\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__47086\,
            I => \N__47016\
        );

    \I__11414\ : InMux
    port map (
            O => \N__47085\,
            I => \N__47011\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47082\,
            I => \N__47011\
        );

    \I__11412\ : InMux
    port map (
            O => \N__47081\,
            I => \N__47006\
        );

    \I__11411\ : InMux
    port map (
            O => \N__47080\,
            I => \N__47006\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__47077\,
            I => \N__47003\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__47074\,
            I => \N__47000\
        );

    \I__11408\ : InMux
    port map (
            O => \N__47073\,
            I => \N__46995\
        );

    \I__11407\ : InMux
    port map (
            O => \N__47072\,
            I => \N__46995\
        );

    \I__11406\ : InMux
    port map (
            O => \N__47071\,
            I => \N__46990\
        );

    \I__11405\ : InMux
    port map (
            O => \N__47070\,
            I => \N__46990\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__47067\,
            I => \N__46987\
        );

    \I__11403\ : InMux
    port map (
            O => \N__47066\,
            I => \N__46978\
        );

    \I__11402\ : InMux
    port map (
            O => \N__47065\,
            I => \N__46978\
        );

    \I__11401\ : InMux
    port map (
            O => \N__47064\,
            I => \N__46978\
        );

    \I__11400\ : InMux
    port map (
            O => \N__47063\,
            I => \N__46978\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__47060\,
            I => \N__46975\
        );

    \I__11398\ : InMux
    port map (
            O => \N__47059\,
            I => \N__46963\
        );

    \I__11397\ : InMux
    port map (
            O => \N__47058\,
            I => \N__46963\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__46945\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__47050\,
            I => \N__46945\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__47047\,
            I => \N__46945\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__47040\,
            I => \N__46945\
        );

    \I__11392\ : Span4Mux_h
    port map (
            O => \N__47037\,
            I => \N__46945\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__46945\
        );

    \I__11390\ : Span4Mux_v
    port map (
            O => \N__47027\,
            I => \N__46940\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__47024\,
            I => \N__46940\
        );

    \I__11388\ : Span4Mux_v
    port map (
            O => \N__47019\,
            I => \N__46933\
        );

    \I__11387\ : Span4Mux_h
    port map (
            O => \N__47016\,
            I => \N__46933\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__47011\,
            I => \N__46933\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__47006\,
            I => \N__46922\
        );

    \I__11384\ : Span4Mux_h
    port map (
            O => \N__47003\,
            I => \N__46922\
        );

    \I__11383\ : Span4Mux_h
    port map (
            O => \N__47000\,
            I => \N__46922\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__46995\,
            I => \N__46922\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__46990\,
            I => \N__46922\
        );

    \I__11380\ : Span12Mux_h
    port map (
            O => \N__46987\,
            I => \N__46919\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__46978\,
            I => \N__46914\
        );

    \I__11378\ : Span12Mux_v
    port map (
            O => \N__46975\,
            I => \N__46914\
        );

    \I__11377\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46899\
        );

    \I__11376\ : InMux
    port map (
            O => \N__46973\,
            I => \N__46899\
        );

    \I__11375\ : InMux
    port map (
            O => \N__46972\,
            I => \N__46899\
        );

    \I__11374\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46899\
        );

    \I__11373\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46899\
        );

    \I__11372\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46899\
        );

    \I__11371\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46899\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__46963\,
            I => \N__46896\
        );

    \I__11369\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46891\
        );

    \I__11368\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46891\
        );

    \I__11367\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46884\
        );

    \I__11366\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46884\
        );

    \I__11365\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46884\
        );

    \I__11364\ : Span4Mux_v
    port map (
            O => \N__46945\,
            I => \N__46879\
        );

    \I__11363\ : Span4Mux_h
    port map (
            O => \N__46940\,
            I => \N__46879\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__46933\,
            I => \N__46874\
        );

    \I__11361\ : Span4Mux_v
    port map (
            O => \N__46922\,
            I => \N__46874\
        );

    \I__11360\ : Odrv12
    port map (
            O => \N__46919\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11359\ : Odrv12
    port map (
            O => \N__46914\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__46899\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__46896\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__46891\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__46884\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11354\ : Odrv4
    port map (
            O => \N__46879\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11353\ : Odrv4
    port map (
            O => \N__46874\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11352\ : CEMux
    port map (
            O => \N__46857\,
            I => \N__46848\
        );

    \I__11351\ : CEMux
    port map (
            O => \N__46856\,
            I => \N__46840\
        );

    \I__11350\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46837\
        );

    \I__11349\ : CEMux
    port map (
            O => \N__46854\,
            I => \N__46834\
        );

    \I__11348\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46831\
        );

    \I__11347\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46828\
        );

    \I__11346\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46825\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46822\
        );

    \I__11344\ : InMux
    port map (
            O => \N__46847\,
            I => \N__46818\
        );

    \I__11343\ : InMux
    port map (
            O => \N__46846\,
            I => \N__46815\
        );

    \I__11342\ : CEMux
    port map (
            O => \N__46845\,
            I => \N__46811\
        );

    \I__11341\ : CEMux
    port map (
            O => \N__46844\,
            I => \N__46808\
        );

    \I__11340\ : CEMux
    port map (
            O => \N__46843\,
            I => \N__46805\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__46840\,
            I => \N__46802\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__46837\,
            I => \N__46799\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__46834\,
            I => \N__46792\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__46831\,
            I => \N__46792\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__46828\,
            I => \N__46792\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46789\
        );

    \I__11333\ : Span4Mux_v
    port map (
            O => \N__46822\,
            I => \N__46786\
        );

    \I__11332\ : CEMux
    port map (
            O => \N__46821\,
            I => \N__46783\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__46818\,
            I => \N__46778\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__46815\,
            I => \N__46778\
        );

    \I__11329\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46775\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__46811\,
            I => \N__46772\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46769\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__46805\,
            I => \N__46762\
        );

    \I__11325\ : Span4Mux_v
    port map (
            O => \N__46802\,
            I => \N__46762\
        );

    \I__11324\ : Span4Mux_h
    port map (
            O => \N__46799\,
            I => \N__46762\
        );

    \I__11323\ : Span4Mux_v
    port map (
            O => \N__46792\,
            I => \N__46757\
        );

    \I__11322\ : Span4Mux_v
    port map (
            O => \N__46789\,
            I => \N__46757\
        );

    \I__11321\ : Span4Mux_h
    port map (
            O => \N__46786\,
            I => \N__46752\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46752\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__46778\,
            I => \N__46747\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__46775\,
            I => \N__46747\
        );

    \I__11317\ : Span12Mux_h
    port map (
            O => \N__46772\,
            I => \N__46744\
        );

    \I__11316\ : Span4Mux_h
    port map (
            O => \N__46769\,
            I => \N__46741\
        );

    \I__11315\ : Span4Mux_h
    port map (
            O => \N__46762\,
            I => \N__46738\
        );

    \I__11314\ : Span4Mux_h
    port map (
            O => \N__46757\,
            I => \N__46735\
        );

    \I__11313\ : Span4Mux_h
    port map (
            O => \N__46752\,
            I => \N__46730\
        );

    \I__11312\ : Span4Mux_h
    port map (
            O => \N__46747\,
            I => \N__46730\
        );

    \I__11311\ : Odrv12
    port map (
            O => \N__46744\,
            I => \data_out_10__7__N_110\
        );

    \I__11310\ : Odrv4
    port map (
            O => \N__46741\,
            I => \data_out_10__7__N_110\
        );

    \I__11309\ : Odrv4
    port map (
            O => \N__46738\,
            I => \data_out_10__7__N_110\
        );

    \I__11308\ : Odrv4
    port map (
            O => \N__46735\,
            I => \data_out_10__7__N_110\
        );

    \I__11307\ : Odrv4
    port map (
            O => \N__46730\,
            I => \data_out_10__7__N_110\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__46719\,
            I => \N__46716\
        );

    \I__11305\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46712\
        );

    \I__11304\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46709\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__46712\,
            I => \N__46704\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__46709\,
            I => \N__46701\
        );

    \I__11301\ : CascadeMux
    port map (
            O => \N__46708\,
            I => \N__46698\
        );

    \I__11300\ : InMux
    port map (
            O => \N__46707\,
            I => \N__46694\
        );

    \I__11299\ : Span4Mux_h
    port map (
            O => \N__46704\,
            I => \N__46691\
        );

    \I__11298\ : Span4Mux_v
    port map (
            O => \N__46701\,
            I => \N__46688\
        );

    \I__11297\ : InMux
    port map (
            O => \N__46698\,
            I => \N__46685\
        );

    \I__11296\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46682\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__46694\,
            I => \N__46679\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__46691\,
            I => \N__46676\
        );

    \I__11293\ : Span4Mux_h
    port map (
            O => \N__46688\,
            I => \N__46671\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__46685\,
            I => \N__46671\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__46682\,
            I => data_out_frame2_5_4
        );

    \I__11290\ : Odrv12
    port map (
            O => \N__46679\,
            I => data_out_frame2_5_4
        );

    \I__11289\ : Odrv4
    port map (
            O => \N__46676\,
            I => data_out_frame2_5_4
        );

    \I__11288\ : Odrv4
    port map (
            O => \N__46671\,
            I => data_out_frame2_5_4
        );

    \I__11287\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__46659\,
            I => \c0.n17856\
        );

    \I__11285\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46649\
        );

    \I__11284\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46649\
        );

    \I__11283\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46646\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__46649\,
            I => \N__46642\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__46646\,
            I => \N__46639\
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__46645\,
            I => \N__46634\
        );

    \I__11279\ : Span4Mux_v
    port map (
            O => \N__46642\,
            I => \N__46629\
        );

    \I__11278\ : Span4Mux_s3_v
    port map (
            O => \N__46639\,
            I => \N__46629\
        );

    \I__11277\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46626\
        );

    \I__11276\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46623\
        );

    \I__11275\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46620\
        );

    \I__11274\ : Span4Mux_h
    port map (
            O => \N__46629\,
            I => \N__46615\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__46626\,
            I => \N__46615\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__46623\,
            I => data_out_frame2_16_2
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__46620\,
            I => data_out_frame2_16_2
        );

    \I__11270\ : Odrv4
    port map (
            O => \N__46615\,
            I => data_out_frame2_16_2
        );

    \I__11269\ : CascadeMux
    port map (
            O => \N__46608\,
            I => \N__46605\
        );

    \I__11268\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46599\
        );

    \I__11267\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46599\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__46599\,
            I => \N__46596\
        );

    \I__11265\ : Span4Mux_h
    port map (
            O => \N__46596\,
            I => \N__46591\
        );

    \I__11264\ : CascadeMux
    port map (
            O => \N__46595\,
            I => \N__46586\
        );

    \I__11263\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46583\
        );

    \I__11262\ : Sp12to4
    port map (
            O => \N__46591\,
            I => \N__46580\
        );

    \I__11261\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46575\
        );

    \I__11260\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46575\
        );

    \I__11259\ : InMux
    port map (
            O => \N__46586\,
            I => \N__46572\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__46583\,
            I => data_out_frame2_9_2
        );

    \I__11257\ : Odrv12
    port map (
            O => \N__46580\,
            I => data_out_frame2_9_2
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__46575\,
            I => data_out_frame2_9_2
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__46572\,
            I => data_out_frame2_9_2
        );

    \I__11254\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46559\
        );

    \I__11253\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46556\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__46559\,
            I => \N__46553\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__46556\,
            I => \N__46550\
        );

    \I__11250\ : Odrv12
    port map (
            O => \N__46553\,
            I => \c0.n10887\
        );

    \I__11249\ : Odrv4
    port map (
            O => \N__46550\,
            I => \c0.n10887\
        );

    \I__11248\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46542\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46539\
        );

    \I__11246\ : Odrv12
    port map (
            O => \N__46539\,
            I => \c0.n16_adj_2399\
        );

    \I__11245\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46530\
        );

    \I__11244\ : InMux
    port map (
            O => \N__46535\,
            I => \N__46527\
        );

    \I__11243\ : InMux
    port map (
            O => \N__46534\,
            I => \N__46524\
        );

    \I__11242\ : InMux
    port map (
            O => \N__46533\,
            I => \N__46521\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__46530\,
            I => \N__46517\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__46527\,
            I => \N__46512\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__46524\,
            I => \N__46512\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__46521\,
            I => \N__46509\
        );

    \I__11237\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46506\
        );

    \I__11236\ : Span4Mux_v
    port map (
            O => \N__46517\,
            I => \N__46503\
        );

    \I__11235\ : Span4Mux_s3_v
    port map (
            O => \N__46512\,
            I => \N__46500\
        );

    \I__11234\ : Span4Mux_h
    port map (
            O => \N__46509\,
            I => \N__46497\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__46506\,
            I => data_out_frame2_10_0
        );

    \I__11232\ : Odrv4
    port map (
            O => \N__46503\,
            I => data_out_frame2_10_0
        );

    \I__11231\ : Odrv4
    port map (
            O => \N__46500\,
            I => data_out_frame2_10_0
        );

    \I__11230\ : Odrv4
    port map (
            O => \N__46497\,
            I => data_out_frame2_10_0
        );

    \I__11229\ : CascadeMux
    port map (
            O => \N__46488\,
            I => \N__46482\
        );

    \I__11228\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46479\
        );

    \I__11227\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46476\
        );

    \I__11226\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46471\
        );

    \I__11225\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46468\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__46479\,
            I => \N__46464\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__46476\,
            I => \N__46461\
        );

    \I__11222\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46458\
        );

    \I__11221\ : CascadeMux
    port map (
            O => \N__46474\,
            I => \N__46455\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__46471\,
            I => \N__46452\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__46468\,
            I => \N__46449\
        );

    \I__11218\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46446\
        );

    \I__11217\ : Span4Mux_v
    port map (
            O => \N__46464\,
            I => \N__46443\
        );

    \I__11216\ : Span4Mux_v
    port map (
            O => \N__46461\,
            I => \N__46440\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__46458\,
            I => \N__46437\
        );

    \I__11214\ : InMux
    port map (
            O => \N__46455\,
            I => \N__46434\
        );

    \I__11213\ : Span4Mux_h
    port map (
            O => \N__46452\,
            I => \N__46429\
        );

    \I__11212\ : Span4Mux_h
    port map (
            O => \N__46449\,
            I => \N__46429\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__46446\,
            I => data_out_frame2_11_0
        );

    \I__11210\ : Odrv4
    port map (
            O => \N__46443\,
            I => data_out_frame2_11_0
        );

    \I__11209\ : Odrv4
    port map (
            O => \N__46440\,
            I => data_out_frame2_11_0
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__46437\,
            I => data_out_frame2_11_0
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__46434\,
            I => data_out_frame2_11_0
        );

    \I__11206\ : Odrv4
    port map (
            O => \N__46429\,
            I => data_out_frame2_11_0
        );

    \I__11205\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46412\
        );

    \I__11204\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46407\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__46412\,
            I => \N__46404\
        );

    \I__11202\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46401\
        );

    \I__11201\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46398\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__46407\,
            I => \N__46394\
        );

    \I__11199\ : Span4Mux_h
    port map (
            O => \N__46404\,
            I => \N__46389\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__46401\,
            I => \N__46389\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__46398\,
            I => \N__46386\
        );

    \I__11196\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46383\
        );

    \I__11195\ : Span4Mux_s1_v
    port map (
            O => \N__46394\,
            I => \N__46379\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__46389\,
            I => \N__46372\
        );

    \I__11193\ : Span4Mux_v
    port map (
            O => \N__46386\,
            I => \N__46372\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__46383\,
            I => \N__46372\
        );

    \I__11191\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46369\
        );

    \I__11190\ : Span4Mux_v
    port map (
            O => \N__46379\,
            I => \N__46366\
        );

    \I__11189\ : Span4Mux_h
    port map (
            O => \N__46372\,
            I => \N__46363\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__46369\,
            I => data_out_frame2_9_0
        );

    \I__11187\ : Odrv4
    port map (
            O => \N__46366\,
            I => data_out_frame2_9_0
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__46363\,
            I => data_out_frame2_9_0
        );

    \I__11185\ : CascadeMux
    port map (
            O => \N__46356\,
            I => \c0.n18891_cascade_\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46349\
        );

    \I__11183\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46346\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__46349\,
            I => \N__46342\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__46346\,
            I => \N__46338\
        );

    \I__11180\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46335\
        );

    \I__11179\ : Span4Mux_h
    port map (
            O => \N__46342\,
            I => \N__46332\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46328\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__46338\,
            I => \N__46325\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46320\
        );

    \I__11175\ : Span4Mux_v
    port map (
            O => \N__46332\,
            I => \N__46320\
        );

    \I__11174\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46317\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__46328\,
            I => data_out_frame2_8_0
        );

    \I__11172\ : Odrv4
    port map (
            O => \N__46325\,
            I => data_out_frame2_8_0
        );

    \I__11171\ : Odrv4
    port map (
            O => \N__46320\,
            I => data_out_frame2_8_0
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__46317\,
            I => data_out_frame2_8_0
        );

    \I__11169\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46305\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46305\,
            I => \N__46300\
        );

    \I__11167\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46297\
        );

    \I__11166\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46294\
        );

    \I__11165\ : Span4Mux_s2_v
    port map (
            O => \N__46300\,
            I => \N__46291\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__46297\,
            I => \N__46288\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46284\
        );

    \I__11162\ : Span4Mux_v
    port map (
            O => \N__46291\,
            I => \N__46279\
        );

    \I__11161\ : Span4Mux_h
    port map (
            O => \N__46288\,
            I => \N__46279\
        );

    \I__11160\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46276\
        );

    \I__11159\ : Span12Mux_s9_v
    port map (
            O => \N__46284\,
            I => \N__46273\
        );

    \I__11158\ : Span4Mux_h
    port map (
            O => \N__46279\,
            I => \N__46270\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__46276\,
            I => data_out_frame2_14_0
        );

    \I__11156\ : Odrv12
    port map (
            O => \N__46273\,
            I => data_out_frame2_14_0
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__46270\,
            I => data_out_frame2_14_0
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__46263\,
            I => \N__46258\
        );

    \I__11153\ : InMux
    port map (
            O => \N__46262\,
            I => \N__46255\
        );

    \I__11152\ : InMux
    port map (
            O => \N__46261\,
            I => \N__46252\
        );

    \I__11151\ : InMux
    port map (
            O => \N__46258\,
            I => \N__46249\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__46255\,
            I => \N__46246\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__46252\,
            I => \N__46243\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__46249\,
            I => \N__46240\
        );

    \I__11147\ : IoSpan4Mux
    port map (
            O => \N__46246\,
            I => \N__46235\
        );

    \I__11146\ : Span4Mux_v
    port map (
            O => \N__46243\,
            I => \N__46235\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__46240\,
            I => \N__46230\
        );

    \I__11144\ : Span4Mux_s0_v
    port map (
            O => \N__46235\,
            I => \N__46227\
        );

    \I__11143\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46222\
        );

    \I__11142\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46222\
        );

    \I__11141\ : Span4Mux_v
    port map (
            O => \N__46230\,
            I => \N__46219\
        );

    \I__11140\ : Odrv4
    port map (
            O => \N__46227\,
            I => data_out_frame2_15_0
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__46222\,
            I => data_out_frame2_15_0
        );

    \I__11138\ : Odrv4
    port map (
            O => \N__46219\,
            I => data_out_frame2_15_0
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__46212\,
            I => \N__46207\
        );

    \I__11136\ : CascadeMux
    port map (
            O => \N__46211\,
            I => \N__46202\
        );

    \I__11135\ : CascadeMux
    port map (
            O => \N__46210\,
            I => \N__46198\
        );

    \I__11134\ : InMux
    port map (
            O => \N__46207\,
            I => \N__46181\
        );

    \I__11133\ : InMux
    port map (
            O => \N__46206\,
            I => \N__46170\
        );

    \I__11132\ : InMux
    port map (
            O => \N__46205\,
            I => \N__46170\
        );

    \I__11131\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46170\
        );

    \I__11130\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46170\
        );

    \I__11129\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46170\
        );

    \I__11128\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46167\
        );

    \I__11127\ : InMux
    port map (
            O => \N__46196\,
            I => \N__46152\
        );

    \I__11126\ : InMux
    port map (
            O => \N__46195\,
            I => \N__46152\
        );

    \I__11125\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46145\
        );

    \I__11124\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46145\
        );

    \I__11123\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46140\
        );

    \I__11122\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46140\
        );

    \I__11121\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46136\
        );

    \I__11120\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46127\
        );

    \I__11119\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46127\
        );

    \I__11118\ : InMux
    port map (
            O => \N__46187\,
            I => \N__46127\
        );

    \I__11117\ : InMux
    port map (
            O => \N__46186\,
            I => \N__46127\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46185\,
            I => \N__46124\
        );

    \I__11115\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46113\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__46181\,
            I => \N__46106\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__46170\,
            I => \N__46106\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__46167\,
            I => \N__46106\
        );

    \I__11111\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46101\
        );

    \I__11110\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46101\
        );

    \I__11109\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46096\
        );

    \I__11108\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46096\
        );

    \I__11107\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46093\
        );

    \I__11106\ : InMux
    port map (
            O => \N__46161\,
            I => \N__46085\
        );

    \I__11105\ : InMux
    port map (
            O => \N__46160\,
            I => \N__46082\
        );

    \I__11104\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46077\
        );

    \I__11103\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46072\
        );

    \I__11102\ : InMux
    port map (
            O => \N__46157\,
            I => \N__46072\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__46152\,
            I => \N__46069\
        );

    \I__11100\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46066\
        );

    \I__11099\ : InMux
    port map (
            O => \N__46150\,
            I => \N__46061\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__46145\,
            I => \N__46056\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__46056\
        );

    \I__11096\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46053\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__46136\,
            I => \N__46046\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__46127\,
            I => \N__46046\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__46124\,
            I => \N__46046\
        );

    \I__11092\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46039\
        );

    \I__11091\ : InMux
    port map (
            O => \N__46122\,
            I => \N__46039\
        );

    \I__11090\ : InMux
    port map (
            O => \N__46121\,
            I => \N__46039\
        );

    \I__11089\ : InMux
    port map (
            O => \N__46120\,
            I => \N__46034\
        );

    \I__11088\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46034\
        );

    \I__11087\ : InMux
    port map (
            O => \N__46118\,
            I => \N__46027\
        );

    \I__11086\ : InMux
    port map (
            O => \N__46117\,
            I => \N__46027\
        );

    \I__11085\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46027\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__46113\,
            I => \N__46018\
        );

    \I__11083\ : Span4Mux_h
    port map (
            O => \N__46106\,
            I => \N__46018\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46101\,
            I => \N__46018\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__46096\,
            I => \N__46018\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__46093\,
            I => \N__46014\
        );

    \I__11079\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46007\
        );

    \I__11078\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46007\
        );

    \I__11077\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46007\
        );

    \I__11076\ : InMux
    port map (
            O => \N__46089\,
            I => \N__46002\
        );

    \I__11075\ : InMux
    port map (
            O => \N__46088\,
            I => \N__46002\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__46085\,
            I => \N__45999\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__46082\,
            I => \N__45996\
        );

    \I__11072\ : InMux
    port map (
            O => \N__46081\,
            I => \N__45993\
        );

    \I__11071\ : InMux
    port map (
            O => \N__46080\,
            I => \N__45990\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__46077\,
            I => \N__45987\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__46072\,
            I => \N__45982\
        );

    \I__11068\ : Span4Mux_v
    port map (
            O => \N__46069\,
            I => \N__45982\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__46066\,
            I => \N__45979\
        );

    \I__11066\ : InMux
    port map (
            O => \N__46065\,
            I => \N__45976\
        );

    \I__11065\ : InMux
    port map (
            O => \N__46064\,
            I => \N__45973\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__46061\,
            I => \N__45968\
        );

    \I__11063\ : Span4Mux_v
    port map (
            O => \N__46056\,
            I => \N__45968\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__46053\,
            I => \N__45963\
        );

    \I__11061\ : Span4Mux_v
    port map (
            O => \N__46046\,
            I => \N__45963\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__46039\,
            I => \N__45956\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__46034\,
            I => \N__45956\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__45956\
        );

    \I__11057\ : Span4Mux_h
    port map (
            O => \N__46018\,
            I => \N__45953\
        );

    \I__11056\ : InMux
    port map (
            O => \N__46017\,
            I => \N__45949\
        );

    \I__11055\ : Span4Mux_s1_v
    port map (
            O => \N__46014\,
            I => \N__45944\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__46007\,
            I => \N__45944\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45939\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__45999\,
            I => \N__45939\
        );

    \I__11051\ : Span4Mux_v
    port map (
            O => \N__45996\,
            I => \N__45936\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__45993\,
            I => \N__45933\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__45990\,
            I => \N__45926\
        );

    \I__11048\ : Span4Mux_v
    port map (
            O => \N__45987\,
            I => \N__45926\
        );

    \I__11047\ : Span4Mux_v
    port map (
            O => \N__45982\,
            I => \N__45926\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__45979\,
            I => \N__45921\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__45976\,
            I => \N__45921\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__45973\,
            I => \N__45916\
        );

    \I__11043\ : Span4Mux_v
    port map (
            O => \N__45968\,
            I => \N__45916\
        );

    \I__11042\ : Span4Mux_v
    port map (
            O => \N__45963\,
            I => \N__45913\
        );

    \I__11041\ : Span4Mux_v
    port map (
            O => \N__45956\,
            I => \N__45908\
        );

    \I__11040\ : Span4Mux_v
    port map (
            O => \N__45953\,
            I => \N__45908\
        );

    \I__11039\ : InMux
    port map (
            O => \N__45952\,
            I => \N__45905\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__45949\,
            I => \N__45902\
        );

    \I__11037\ : Span4Mux_v
    port map (
            O => \N__45944\,
            I => \N__45899\
        );

    \I__11036\ : Span4Mux_h
    port map (
            O => \N__45939\,
            I => \N__45896\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__45936\,
            I => \N__45889\
        );

    \I__11034\ : Span4Mux_v
    port map (
            O => \N__45933\,
            I => \N__45889\
        );

    \I__11033\ : Span4Mux_h
    port map (
            O => \N__45926\,
            I => \N__45889\
        );

    \I__11032\ : Span4Mux_h
    port map (
            O => \N__45921\,
            I => \N__45886\
        );

    \I__11031\ : Span4Mux_h
    port map (
            O => \N__45916\,
            I => \N__45881\
        );

    \I__11030\ : Span4Mux_h
    port map (
            O => \N__45913\,
            I => \N__45881\
        );

    \I__11029\ : Span4Mux_h
    port map (
            O => \N__45908\,
            I => \N__45878\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__45905\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11027\ : Odrv12
    port map (
            O => \N__45902\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11026\ : Odrv4
    port map (
            O => \N__45899\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11025\ : Odrv4
    port map (
            O => \N__45896\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11024\ : Odrv4
    port map (
            O => \N__45889\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__45886\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11022\ : Odrv4
    port map (
            O => \N__45881\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11021\ : Odrv4
    port map (
            O => \N__45878\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__45861\,
            I => \N__45858\
        );

    \I__11019\ : InMux
    port map (
            O => \N__45858\,
            I => \N__45853\
        );

    \I__11018\ : InMux
    port map (
            O => \N__45857\,
            I => \N__45850\
        );

    \I__11017\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45846\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45843\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45840\
        );

    \I__11014\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45837\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__45846\,
            I => \N__45834\
        );

    \I__11012\ : Span4Mux_h
    port map (
            O => \N__45843\,
            I => \N__45831\
        );

    \I__11011\ : Span4Mux_v
    port map (
            O => \N__45840\,
            I => \N__45828\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__45837\,
            I => data_out_frame2_13_0
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__45834\,
            I => data_out_frame2_13_0
        );

    \I__11008\ : Odrv4
    port map (
            O => \N__45831\,
            I => data_out_frame2_13_0
        );

    \I__11007\ : Odrv4
    port map (
            O => \N__45828\,
            I => data_out_frame2_13_0
        );

    \I__11006\ : CascadeMux
    port map (
            O => \N__45819\,
            I => \c0.n18897_cascade_\
        );

    \I__11005\ : InMux
    port map (
            O => \N__45816\,
            I => \N__45811\
        );

    \I__11004\ : InMux
    port map (
            O => \N__45815\,
            I => \N__45808\
        );

    \I__11003\ : InMux
    port map (
            O => \N__45814\,
            I => \N__45805\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45802\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__45808\,
            I => \N__45798\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__45805\,
            I => \N__45795\
        );

    \I__10999\ : Span4Mux_v
    port map (
            O => \N__45802\,
            I => \N__45792\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__45801\,
            I => \N__45786\
        );

    \I__10997\ : Span4Mux_s3_v
    port map (
            O => \N__45798\,
            I => \N__45781\
        );

    \I__10996\ : Span4Mux_s3_v
    port map (
            O => \N__45795\,
            I => \N__45781\
        );

    \I__10995\ : Span4Mux_v
    port map (
            O => \N__45792\,
            I => \N__45778\
        );

    \I__10994\ : InMux
    port map (
            O => \N__45791\,
            I => \N__45773\
        );

    \I__10993\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45773\
        );

    \I__10992\ : InMux
    port map (
            O => \N__45789\,
            I => \N__45770\
        );

    \I__10991\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45767\
        );

    \I__10990\ : Span4Mux_h
    port map (
            O => \N__45781\,
            I => \N__45763\
        );

    \I__10989\ : Span4Mux_s1_v
    port map (
            O => \N__45778\,
            I => \N__45758\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__45773\,
            I => \N__45758\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__45770\,
            I => \N__45755\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__45767\,
            I => \N__45752\
        );

    \I__10985\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45749\
        );

    \I__10984\ : Sp12to4
    port map (
            O => \N__45763\,
            I => \N__45746\
        );

    \I__10983\ : Span4Mux_h
    port map (
            O => \N__45758\,
            I => \N__45739\
        );

    \I__10982\ : Span4Mux_h
    port map (
            O => \N__45755\,
            I => \N__45739\
        );

    \I__10981\ : Span4Mux_h
    port map (
            O => \N__45752\,
            I => \N__45739\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__45749\,
            I => data_out_frame2_12_0
        );

    \I__10979\ : Odrv12
    port map (
            O => \N__45746\,
            I => data_out_frame2_12_0
        );

    \I__10978\ : Odrv4
    port map (
            O => \N__45739\,
            I => data_out_frame2_12_0
        );

    \I__10977\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__45729\,
            I => \c0.n18060\
        );

    \I__10975\ : CascadeMux
    port map (
            O => \N__45726\,
            I => \c0.n18057_cascade_\
        );

    \I__10974\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45720\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__45720\,
            I => \N__45717\
        );

    \I__10972\ : Odrv12
    port map (
            O => \N__45717\,
            I => \c0.n18374\
        );

    \I__10971\ : CascadeMux
    port map (
            O => \N__45714\,
            I => \c0.n18723_cascade_\
        );

    \I__10970\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__45708\,
            I => \N__45705\
        );

    \I__10968\ : Span4Mux_v
    port map (
            O => \N__45705\,
            I => \N__45702\
        );

    \I__10967\ : Span4Mux_h
    port map (
            O => \N__45702\,
            I => \N__45699\
        );

    \I__10966\ : Odrv4
    port map (
            O => \N__45699\,
            I => \c0.n6_adj_2275\
        );

    \I__10965\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45692\
        );

    \I__10964\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45689\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__45692\,
            I => \N__45684\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__45689\,
            I => \N__45684\
        );

    \I__10961\ : Span4Mux_s3_v
    port map (
            O => \N__45684\,
            I => \N__45679\
        );

    \I__10960\ : InMux
    port map (
            O => \N__45683\,
            I => \N__45674\
        );

    \I__10959\ : InMux
    port map (
            O => \N__45682\,
            I => \N__45674\
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__45679\,
            I => \c0.n17810\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__45674\,
            I => \c0.n17810\
        );

    \I__10956\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45664\
        );

    \I__10955\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45659\
        );

    \I__10954\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45659\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__45664\,
            I => \N__45656\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__45659\,
            I => \N__45651\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__45656\,
            I => \N__45647\
        );

    \I__10950\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45642\
        );

    \I__10949\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45642\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__45651\,
            I => \N__45639\
        );

    \I__10947\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45636\
        );

    \I__10946\ : Odrv4
    port map (
            O => \N__45647\,
            I => data_out_frame2_11_2
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__45642\,
            I => data_out_frame2_11_2
        );

    \I__10944\ : Odrv4
    port map (
            O => \N__45639\,
            I => data_out_frame2_11_2
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__45636\,
            I => data_out_frame2_11_2
        );

    \I__10942\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45622\
        );

    \I__10941\ : CascadeMux
    port map (
            O => \N__45626\,
            I => \N__45618\
        );

    \I__10940\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45615\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45610\
        );

    \I__10938\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45605\
        );

    \I__10937\ : InMux
    port map (
            O => \N__45618\,
            I => \N__45605\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__45615\,
            I => \N__45602\
        );

    \I__10935\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45599\
        );

    \I__10934\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45596\
        );

    \I__10933\ : Span4Mux_s1_v
    port map (
            O => \N__45610\,
            I => \N__45593\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__45605\,
            I => \N__45590\
        );

    \I__10931\ : Span4Mux_h
    port map (
            O => \N__45602\,
            I => \N__45587\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__45599\,
            I => data_out_frame2_11_3
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__45596\,
            I => data_out_frame2_11_3
        );

    \I__10928\ : Odrv4
    port map (
            O => \N__45593\,
            I => data_out_frame2_11_3
        );

    \I__10927\ : Odrv12
    port map (
            O => \N__45590\,
            I => data_out_frame2_11_3
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__45587\,
            I => data_out_frame2_11_3
        );

    \I__10925\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45571\
        );

    \I__10924\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45567\
        );

    \I__10923\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45564\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__45571\,
            I => \N__45561\
        );

    \I__10921\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45558\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__45567\,
            I => \N__45555\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__45564\,
            I => data_out_frame2_11_1
        );

    \I__10918\ : Odrv12
    port map (
            O => \N__45561\,
            I => data_out_frame2_11_1
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__45558\,
            I => data_out_frame2_11_1
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__45555\,
            I => data_out_frame2_11_1
        );

    \I__10915\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45543\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__45543\,
            I => \c0.n17798\
        );

    \I__10913\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45537\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__45537\,
            I => \N__45533\
        );

    \I__10911\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45530\
        );

    \I__10910\ : Span4Mux_v
    port map (
            O => \N__45533\,
            I => \N__45527\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__45530\,
            I => \N__45524\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__45527\,
            I => \N__45520\
        );

    \I__10907\ : Span4Mux_s1_v
    port map (
            O => \N__45524\,
            I => \N__45517\
        );

    \I__10906\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45514\
        );

    \I__10905\ : Odrv4
    port map (
            O => \N__45520\,
            I => \c0.n17751\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__45517\,
            I => \c0.n17751\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__45514\,
            I => \c0.n17751\
        );

    \I__10902\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45503\
        );

    \I__10901\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45500\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__45503\,
            I => \N__45497\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__45500\,
            I => \N__45494\
        );

    \I__10898\ : Odrv4
    port map (
            O => \N__45497\,
            I => \c0.n17868\
        );

    \I__10897\ : Odrv12
    port map (
            O => \N__45494\,
            I => \c0.n17868\
        );

    \I__10896\ : CascadeMux
    port map (
            O => \N__45489\,
            I => \c0.n17798_cascade_\
        );

    \I__10895\ : InMux
    port map (
            O => \N__45486\,
            I => \N__45483\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__45483\,
            I => \N__45479\
        );

    \I__10893\ : InMux
    port map (
            O => \N__45482\,
            I => \N__45476\
        );

    \I__10892\ : Span4Mux_h
    port map (
            O => \N__45479\,
            I => \N__45473\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__45476\,
            I => \c0.n17902\
        );

    \I__10890\ : Odrv4
    port map (
            O => \N__45473\,
            I => \c0.n17902\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45468\,
            I => \N__45465\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__45465\,
            I => \c0.n18_adj_2393\
        );

    \I__10887\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45459\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__45459\,
            I => \N__45456\
        );

    \I__10885\ : Span4Mux_v
    port map (
            O => \N__45456\,
            I => \N__45451\
        );

    \I__10884\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45448\
        );

    \I__10883\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45445\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__45451\,
            I => \N__45439\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__45448\,
            I => \N__45439\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__45445\,
            I => \N__45436\
        );

    \I__10879\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45432\
        );

    \I__10878\ : Span4Mux_s1_v
    port map (
            O => \N__45439\,
            I => \N__45427\
        );

    \I__10877\ : Span4Mux_h
    port map (
            O => \N__45436\,
            I => \N__45427\
        );

    \I__10876\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45424\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__45432\,
            I => data_out_frame2_16_5
        );

    \I__10874\ : Odrv4
    port map (
            O => \N__45427\,
            I => data_out_frame2_16_5
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__45424\,
            I => data_out_frame2_16_5
        );

    \I__10872\ : CascadeMux
    port map (
            O => \N__45417\,
            I => \c0.n24_adj_2394_cascade_\
        );

    \I__10871\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__45411\,
            I => \N__45407\
        );

    \I__10869\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45404\
        );

    \I__10868\ : Span4Mux_v
    port map (
            O => \N__45407\,
            I => \N__45398\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__45404\,
            I => \N__45398\
        );

    \I__10866\ : CascadeMux
    port map (
            O => \N__45403\,
            I => \N__45395\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__45398\,
            I => \N__45391\
        );

    \I__10864\ : InMux
    port map (
            O => \N__45395\,
            I => \N__45386\
        );

    \I__10863\ : InMux
    port map (
            O => \N__45394\,
            I => \N__45386\
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__45391\,
            I => data_out_frame2_15_5
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__45386\,
            I => data_out_frame2_15_5
        );

    \I__10860\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45375\
        );

    \I__10859\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45375\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__45375\,
            I => \N__45372\
        );

    \I__10857\ : Odrv4
    port map (
            O => \N__45372\,
            I => \c0.n17920\
        );

    \I__10856\ : InMux
    port map (
            O => \N__45369\,
            I => \N__45366\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__45366\,
            I => \N__45363\
        );

    \I__10854\ : Odrv12
    port map (
            O => \N__45363\,
            I => \c0.n22_adj_2395\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__45360\,
            I => \c0.n26_adj_2396_cascade_\
        );

    \I__10852\ : InMux
    port map (
            O => \N__45357\,
            I => \N__45354\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45350\
        );

    \I__10850\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45347\
        );

    \I__10849\ : Span4Mux_h
    port map (
            O => \N__45350\,
            I => \N__45344\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__45347\,
            I => \N__45339\
        );

    \I__10847\ : Span4Mux_h
    port map (
            O => \N__45344\,
            I => \N__45339\
        );

    \I__10846\ : Odrv4
    port map (
            O => \N__45339\,
            I => \c0.n17917\
        );

    \I__10845\ : CascadeMux
    port map (
            O => \N__45336\,
            I => \N__45333\
        );

    \I__10844\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45330\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45327\
        );

    \I__10842\ : Span4Mux_h
    port map (
            O => \N__45327\,
            I => \N__45324\
        );

    \I__10841\ : Span4Mux_h
    port map (
            O => \N__45324\,
            I => \N__45321\
        );

    \I__10840\ : Sp12to4
    port map (
            O => \N__45321\,
            I => \N__45318\
        );

    \I__10839\ : Odrv12
    port map (
            O => \N__45318\,
            I => \c0.data_out_frame2_20_7\
        );

    \I__10838\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45312\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__45312\,
            I => \N__45309\
        );

    \I__10836\ : Span4Mux_v
    port map (
            O => \N__45309\,
            I => \N__45306\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__45306\,
            I => \N__45302\
        );

    \I__10834\ : InMux
    port map (
            O => \N__45305\,
            I => \N__45299\
        );

    \I__10833\ : Sp12to4
    port map (
            O => \N__45302\,
            I => \N__45296\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45293\
        );

    \I__10831\ : Odrv12
    port map (
            O => \N__45296\,
            I => \c0.n10778\
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__45293\,
            I => \c0.n10778\
        );

    \I__10829\ : InMux
    port map (
            O => \N__45288\,
            I => \N__45284\
        );

    \I__10828\ : InMux
    port map (
            O => \N__45287\,
            I => \N__45281\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__45284\,
            I => \N__45278\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__45281\,
            I => \N__45275\
        );

    \I__10825\ : Odrv4
    port map (
            O => \N__45278\,
            I => \c0.n17871\
        );

    \I__10824\ : Odrv4
    port map (
            O => \N__45275\,
            I => \c0.n17871\
        );

    \I__10823\ : CascadeMux
    port map (
            O => \N__45270\,
            I => \c0.n14_adj_2406_cascade_\
        );

    \I__10822\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45260\
        );

    \I__10820\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45257\
        );

    \I__10819\ : Span4Mux_s1_v
    port map (
            O => \N__45260\,
            I => \N__45254\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__45257\,
            I => \c0.n10583\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__45254\,
            I => \c0.n10583\
        );

    \I__10816\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45245\
        );

    \I__10815\ : InMux
    port map (
            O => \N__45248\,
            I => \N__45241\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__45245\,
            I => \N__45238\
        );

    \I__10813\ : InMux
    port map (
            O => \N__45244\,
            I => \N__45235\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__45241\,
            I => \N__45230\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__45238\,
            I => \N__45225\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45225\
        );

    \I__10809\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45222\
        );

    \I__10808\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45219\
        );

    \I__10807\ : Span4Mux_h
    port map (
            O => \N__45230\,
            I => \N__45214\
        );

    \I__10806\ : Span4Mux_h
    port map (
            O => \N__45225\,
            I => \N__45214\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__45222\,
            I => data_out_frame2_11_5
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__45219\,
            I => data_out_frame2_11_5
        );

    \I__10803\ : Odrv4
    port map (
            O => \N__45214\,
            I => data_out_frame2_11_5
        );

    \I__10802\ : CascadeMux
    port map (
            O => \N__45207\,
            I => \N__45203\
        );

    \I__10801\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45198\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45195\
        );

    \I__10799\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45192\
        );

    \I__10798\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45189\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__45198\,
            I => \N__45186\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__45195\,
            I => \N__45182\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__45192\,
            I => \N__45179\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__45189\,
            I => \N__45176\
        );

    \I__10793\ : Span4Mux_h
    port map (
            O => \N__45186\,
            I => \N__45173\
        );

    \I__10792\ : InMux
    port map (
            O => \N__45185\,
            I => \N__45170\
        );

    \I__10791\ : Span4Mux_h
    port map (
            O => \N__45182\,
            I => \N__45167\
        );

    \I__10790\ : Span12Mux_s11_h
    port map (
            O => \N__45179\,
            I => \N__45164\
        );

    \I__10789\ : Span4Mux_h
    port map (
            O => \N__45176\,
            I => \N__45161\
        );

    \I__10788\ : Span4Mux_v
    port map (
            O => \N__45173\,
            I => \N__45158\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__45170\,
            I => data_out_frame2_12_4
        );

    \I__10786\ : Odrv4
    port map (
            O => \N__45167\,
            I => data_out_frame2_12_4
        );

    \I__10785\ : Odrv12
    port map (
            O => \N__45164\,
            I => data_out_frame2_12_4
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__45161\,
            I => data_out_frame2_12_4
        );

    \I__10783\ : Odrv4
    port map (
            O => \N__45158\,
            I => data_out_frame2_12_4
        );

    \I__10782\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45143\
        );

    \I__10781\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45140\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__45143\,
            I => \N__45137\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__45140\,
            I => \N__45134\
        );

    \I__10778\ : Span4Mux_h
    port map (
            O => \N__45137\,
            I => \N__45131\
        );

    \I__10777\ : Span4Mux_s3_v
    port map (
            O => \N__45134\,
            I => \N__45128\
        );

    \I__10776\ : Odrv4
    port map (
            O => \N__45131\,
            I => \c0.n17780\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__45128\,
            I => \c0.n17780\
        );

    \I__10774\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__45120\,
            I => \c0.n15_adj_2407\
        );

    \I__10772\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45108\
        );

    \I__10771\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45108\
        );

    \I__10770\ : InMux
    port map (
            O => \N__45115\,
            I => \N__45108\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__45108\,
            I => \N__45104\
        );

    \I__10768\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45101\
        );

    \I__10767\ : Span4Mux_s3_v
    port map (
            O => \N__45104\,
            I => \N__45098\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__45101\,
            I => data_out_frame2_7_3
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__45098\,
            I => data_out_frame2_7_3
        );

    \I__10764\ : InMux
    port map (
            O => \N__45093\,
            I => \N__45089\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__45092\,
            I => \N__45085\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__45089\,
            I => \N__45082\
        );

    \I__10761\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45079\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45085\,
            I => \N__45074\
        );

    \I__10759\ : Span4Mux_v
    port map (
            O => \N__45082\,
            I => \N__45071\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__45079\,
            I => \N__45068\
        );

    \I__10757\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45065\
        );

    \I__10756\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45062\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__45074\,
            I => \N__45055\
        );

    \I__10754\ : Span4Mux_h
    port map (
            O => \N__45071\,
            I => \N__45055\
        );

    \I__10753\ : Span4Mux_v
    port map (
            O => \N__45068\,
            I => \N__45055\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__45065\,
            I => \N__45052\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__45062\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__10750\ : Odrv4
    port map (
            O => \N__45055\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__10749\ : Odrv12
    port map (
            O => \N__45052\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__10748\ : InMux
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__45042\,
            I => \N__45036\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45041\,
            I => \N__45033\
        );

    \I__10745\ : InMux
    port map (
            O => \N__45040\,
            I => \N__45030\
        );

    \I__10744\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45027\
        );

    \I__10743\ : Span4Mux_h
    port map (
            O => \N__45036\,
            I => \N__45022\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45022\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__45030\,
            I => data_out_frame2_14_3
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__45027\,
            I => data_out_frame2_14_3
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__45022\,
            I => data_out_frame2_14_3
        );

    \I__10738\ : InMux
    port map (
            O => \N__45015\,
            I => \N__45010\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45014\,
            I => \N__45007\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45013\,
            I => \N__45004\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__44998\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__45007\,
            I => \N__44998\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44995\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44991\
        );

    \I__10731\ : Span4Mux_h
    port map (
            O => \N__44998\,
            I => \N__44988\
        );

    \I__10730\ : Span4Mux_h
    port map (
            O => \N__44995\,
            I => \N__44985\
        );

    \I__10729\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44982\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__44991\,
            I => data_out_frame2_15_4
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__44988\,
            I => data_out_frame2_15_4
        );

    \I__10726\ : Odrv4
    port map (
            O => \N__44985\,
            I => data_out_frame2_15_4
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__44982\,
            I => data_out_frame2_15_4
        );

    \I__10724\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44968\
        );

    \I__10723\ : CascadeMux
    port map (
            O => \N__44972\,
            I => \N__44964\
        );

    \I__10722\ : CascadeMux
    port map (
            O => \N__44971\,
            I => \N__44961\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__44968\,
            I => \N__44958\
        );

    \I__10720\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44953\
        );

    \I__10719\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44953\
        );

    \I__10718\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44950\
        );

    \I__10717\ : Span4Mux_s3_v
    port map (
            O => \N__44958\,
            I => \N__44944\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44944\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44941\
        );

    \I__10714\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44938\
        );

    \I__10713\ : Span4Mux_v
    port map (
            O => \N__44944\,
            I => \N__44933\
        );

    \I__10712\ : Span4Mux_h
    port map (
            O => \N__44941\,
            I => \N__44933\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__44938\,
            I => data_out_frame2_7_4
        );

    \I__10710\ : Odrv4
    port map (
            O => \N__44933\,
            I => data_out_frame2_7_4
        );

    \I__10709\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44925\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__44925\,
            I => \c0.n10710\
        );

    \I__10707\ : CascadeMux
    port map (
            O => \N__44922\,
            I => \c0.n10710_cascade_\
        );

    \I__10706\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44916\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__44916\,
            I => \c0.n18_adj_2402\
        );

    \I__10704\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44910\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__44910\,
            I => \N__44907\
        );

    \I__10702\ : Span4Mux_s3_v
    port map (
            O => \N__44907\,
            I => \N__44904\
        );

    \I__10701\ : Odrv4
    port map (
            O => \N__44904\,
            I => \c0.n20_adj_2404\
        );

    \I__10700\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44895\
        );

    \I__10699\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44892\
        );

    \I__10698\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44889\
        );

    \I__10697\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44885\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44880\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44880\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__44889\,
            I => \N__44877\
        );

    \I__10693\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44874\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__44885\,
            I => \N__44871\
        );

    \I__10691\ : Span4Mux_h
    port map (
            O => \N__44880\,
            I => \N__44866\
        );

    \I__10690\ : Span4Mux_s3_v
    port map (
            O => \N__44877\,
            I => \N__44866\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__44874\,
            I => data_out_frame2_6_5
        );

    \I__10688\ : Odrv4
    port map (
            O => \N__44871\,
            I => data_out_frame2_6_5
        );

    \I__10687\ : Odrv4
    port map (
            O => \N__44866\,
            I => data_out_frame2_6_5
        );

    \I__10686\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44854\
        );

    \I__10685\ : InMux
    port map (
            O => \N__44858\,
            I => \N__44847\
        );

    \I__10684\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44847\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__44854\,
            I => \N__44844\
        );

    \I__10682\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44841\
        );

    \I__10681\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44838\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__44847\,
            I => \N__44835\
        );

    \I__10679\ : Span4Mux_h
    port map (
            O => \N__44844\,
            I => \N__44832\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__44841\,
            I => \N__44829\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__44838\,
            I => data_out_frame2_7_5
        );

    \I__10676\ : Odrv12
    port map (
            O => \N__44835\,
            I => data_out_frame2_7_5
        );

    \I__10675\ : Odrv4
    port map (
            O => \N__44832\,
            I => data_out_frame2_7_5
        );

    \I__10674\ : Odrv4
    port map (
            O => \N__44829\,
            I => data_out_frame2_7_5
        );

    \I__10673\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44817\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__44817\,
            I => \N__44814\
        );

    \I__10671\ : Odrv12
    port map (
            O => \N__44814\,
            I => \c0.n5_adj_2386\
        );

    \I__10670\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44807\
        );

    \I__10669\ : InMux
    port map (
            O => \N__44810\,
            I => \N__44802\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__44807\,
            I => \N__44799\
        );

    \I__10667\ : InMux
    port map (
            O => \N__44806\,
            I => \N__44796\
        );

    \I__10666\ : CascadeMux
    port map (
            O => \N__44805\,
            I => \N__44793\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44789\
        );

    \I__10664\ : Span4Mux_v
    port map (
            O => \N__44799\,
            I => \N__44786\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44783\
        );

    \I__10662\ : InMux
    port map (
            O => \N__44793\,
            I => \N__44780\
        );

    \I__10661\ : InMux
    port map (
            O => \N__44792\,
            I => \N__44777\
        );

    \I__10660\ : Span4Mux_h
    port map (
            O => \N__44789\,
            I => \N__44774\
        );

    \I__10659\ : Span4Mux_h
    port map (
            O => \N__44786\,
            I => \N__44771\
        );

    \I__10658\ : Span4Mux_h
    port map (
            O => \N__44783\,
            I => \N__44768\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__44780\,
            I => \N__44765\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__44777\,
            I => data_out_frame2_13_5
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__44774\,
            I => data_out_frame2_13_5
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__44771\,
            I => data_out_frame2_13_5
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__44768\,
            I => data_out_frame2_13_5
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__44765\,
            I => data_out_frame2_13_5
        );

    \I__10651\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44750\
        );

    \I__10650\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44746\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__44750\,
            I => \N__44743\
        );

    \I__10648\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44738\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__44746\,
            I => \N__44735\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__44743\,
            I => \N__44732\
        );

    \I__10645\ : InMux
    port map (
            O => \N__44742\,
            I => \N__44727\
        );

    \I__10644\ : InMux
    port map (
            O => \N__44741\,
            I => \N__44727\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__44738\,
            I => data_out_frame2_10_7
        );

    \I__10642\ : Odrv12
    port map (
            O => \N__44735\,
            I => data_out_frame2_10_7
        );

    \I__10641\ : Odrv4
    port map (
            O => \N__44732\,
            I => data_out_frame2_10_7
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__44727\,
            I => data_out_frame2_10_7
        );

    \I__10639\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__44715\,
            I => \c0.n10877\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__44712\,
            I => \c0.n10593_cascade_\
        );

    \I__10636\ : InMux
    port map (
            O => \N__44709\,
            I => \N__44706\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__44706\,
            I => \N__44703\
        );

    \I__10634\ : Span4Mux_h
    port map (
            O => \N__44703\,
            I => \N__44700\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__44700\,
            I => \c0.n14\
        );

    \I__10632\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44691\
        );

    \I__10631\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44691\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__44691\,
            I => \N__44687\
        );

    \I__10629\ : InMux
    port map (
            O => \N__44690\,
            I => \N__44684\
        );

    \I__10628\ : Span4Mux_v
    port map (
            O => \N__44687\,
            I => \N__44678\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__44684\,
            I => \N__44678\
        );

    \I__10626\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44674\
        );

    \I__10625\ : Span4Mux_h
    port map (
            O => \N__44678\,
            I => \N__44671\
        );

    \I__10624\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44668\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__44674\,
            I => data_out_frame2_7_6
        );

    \I__10622\ : Odrv4
    port map (
            O => \N__44671\,
            I => data_out_frame2_7_6
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__44668\,
            I => data_out_frame2_7_6
        );

    \I__10620\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44656\
        );

    \I__10619\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44653\
        );

    \I__10618\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44650\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__44656\,
            I => \N__44646\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__44653\,
            I => \N__44641\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__44650\,
            I => \N__44641\
        );

    \I__10614\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44638\
        );

    \I__10613\ : Span4Mux_h
    port map (
            O => \N__44646\,
            I => \N__44635\
        );

    \I__10612\ : Span4Mux_s3_v
    port map (
            O => \N__44641\,
            I => \N__44632\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__44638\,
            I => data_out_frame2_5_7
        );

    \I__10610\ : Odrv4
    port map (
            O => \N__44635\,
            I => data_out_frame2_5_7
        );

    \I__10609\ : Odrv4
    port map (
            O => \N__44632\,
            I => data_out_frame2_5_7
        );

    \I__10608\ : CascadeMux
    port map (
            O => \N__44625\,
            I => \N__44621\
        );

    \I__10607\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44618\
        );

    \I__10606\ : InMux
    port map (
            O => \N__44621\,
            I => \N__44615\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__44618\,
            I => \N__44610\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__44615\,
            I => \N__44607\
        );

    \I__10603\ : InMux
    port map (
            O => \N__44614\,
            I => \N__44604\
        );

    \I__10602\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44601\
        );

    \I__10601\ : Span4Mux_h
    port map (
            O => \N__44610\,
            I => \N__44594\
        );

    \I__10600\ : Span4Mux_v
    port map (
            O => \N__44607\,
            I => \N__44594\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__44604\,
            I => \N__44594\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__44601\,
            I => data_out_frame2_9_5
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__44594\,
            I => data_out_frame2_9_5
        );

    \I__10596\ : CascadeMux
    port map (
            O => \N__44589\,
            I => \N__44586\
        );

    \I__10595\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44583\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__44583\,
            I => \N__44578\
        );

    \I__10593\ : InMux
    port map (
            O => \N__44582\,
            I => \N__44575\
        );

    \I__10592\ : CascadeMux
    port map (
            O => \N__44581\,
            I => \N__44572\
        );

    \I__10591\ : Span4Mux_s1_v
    port map (
            O => \N__44578\,
            I => \N__44568\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__44575\,
            I => \N__44565\
        );

    \I__10589\ : InMux
    port map (
            O => \N__44572\,
            I => \N__44561\
        );

    \I__10588\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44558\
        );

    \I__10587\ : Span4Mux_v
    port map (
            O => \N__44568\,
            I => \N__44555\
        );

    \I__10586\ : Span4Mux_s3_v
    port map (
            O => \N__44565\,
            I => \N__44552\
        );

    \I__10585\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44549\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__44561\,
            I => \N__44546\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__44558\,
            I => data_out_frame2_9_3
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__44555\,
            I => data_out_frame2_9_3
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__44552\,
            I => data_out_frame2_9_3
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__44549\,
            I => data_out_frame2_9_3
        );

    \I__10579\ : Odrv12
    port map (
            O => \N__44546\,
            I => data_out_frame2_9_3
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__44535\,
            I => \N__44532\
        );

    \I__10577\ : InMux
    port map (
            O => \N__44532\,
            I => \N__44529\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__44529\,
            I => \c0.n10929\
        );

    \I__10575\ : CascadeMux
    port map (
            O => \N__44526\,
            I => \c0.n10929_cascade_\
        );

    \I__10574\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44520\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__44520\,
            I => \c0.n17823\
        );

    \I__10572\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44514\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44510\
        );

    \I__10570\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44507\
        );

    \I__10569\ : Odrv12
    port map (
            O => \N__44510\,
            I => \c0.n17853\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__44507\,
            I => \c0.n17853\
        );

    \I__10567\ : CascadeMux
    port map (
            O => \N__44502\,
            I => \c0.n17823_cascade_\
        );

    \I__10566\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44496\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__44496\,
            I => \c0.n17895\
        );

    \I__10564\ : CascadeMux
    port map (
            O => \N__44493\,
            I => \c0.n17_adj_2401_cascade_\
        );

    \I__10563\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44486\
        );

    \I__10562\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44483\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__44486\,
            I => \N__44480\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__44483\,
            I => \N__44477\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__44480\,
            I => \N__44474\
        );

    \I__10558\ : Odrv4
    port map (
            O => \N__44477\,
            I => \c0.n17914\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__44474\,
            I => \c0.n17914\
        );

    \I__10556\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44466\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__44466\,
            I => \N__44463\
        );

    \I__10554\ : Span4Mux_v
    port map (
            O => \N__44463\,
            I => \N__44460\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__44460\,
            I => \c0.data_out_frame2_20_6\
        );

    \I__10552\ : InMux
    port map (
            O => \N__44457\,
            I => \N__44454\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__44454\,
            I => \N__44450\
        );

    \I__10550\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44447\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__44450\,
            I => \N__44444\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__44447\,
            I => \c0.n10703\
        );

    \I__10547\ : Odrv4
    port map (
            O => \N__44444\,
            I => \c0.n10703\
        );

    \I__10546\ : CascadeMux
    port map (
            O => \N__44439\,
            I => \N__44434\
        );

    \I__10545\ : CascadeMux
    port map (
            O => \N__44438\,
            I => \N__44430\
        );

    \I__10544\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44427\
        );

    \I__10543\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44424\
        );

    \I__10542\ : InMux
    port map (
            O => \N__44433\,
            I => \N__44419\
        );

    \I__10541\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44419\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44415\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__44424\,
            I => \N__44412\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__44419\,
            I => \N__44409\
        );

    \I__10537\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44406\
        );

    \I__10536\ : Span12Mux_s5_v
    port map (
            O => \N__44415\,
            I => \N__44403\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__44412\,
            I => \N__44400\
        );

    \I__10534\ : Span4Mux_v
    port map (
            O => \N__44409\,
            I => \N__44397\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__44406\,
            I => data_out_frame2_14_4
        );

    \I__10532\ : Odrv12
    port map (
            O => \N__44403\,
            I => data_out_frame2_14_4
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__44400\,
            I => data_out_frame2_14_4
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__44397\,
            I => data_out_frame2_14_4
        );

    \I__10529\ : InMux
    port map (
            O => \N__44388\,
            I => \N__44385\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__44385\,
            I => \N__44382\
        );

    \I__10527\ : Span4Mux_h
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__10526\ : Odrv4
    port map (
            O => \N__44379\,
            I => \c0.n10825\
        );

    \I__10525\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44371\
        );

    \I__10524\ : InMux
    port map (
            O => \N__44375\,
            I => \N__44368\
        );

    \I__10523\ : InMux
    port map (
            O => \N__44374\,
            I => \N__44364\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__44371\,
            I => \N__44361\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44358\
        );

    \I__10520\ : CascadeMux
    port map (
            O => \N__44367\,
            I => \N__44355\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__44364\,
            I => \N__44352\
        );

    \I__10518\ : Span4Mux_h
    port map (
            O => \N__44361\,
            I => \N__44347\
        );

    \I__10517\ : Span4Mux_s2_v
    port map (
            O => \N__44358\,
            I => \N__44347\
        );

    \I__10516\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44344\
        );

    \I__10515\ : Span4Mux_h
    port map (
            O => \N__44352\,
            I => \N__44341\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__44347\,
            I => \N__44338\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__44344\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__44341\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__10511\ : Odrv4
    port map (
            O => \N__44338\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__10510\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44326\
        );

    \I__10509\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44321\
        );

    \I__10508\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44318\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__44326\,
            I => \N__44315\
        );

    \I__10506\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44310\
        );

    \I__10505\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44310\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__44321\,
            I => \N__44304\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__44318\,
            I => \N__44304\
        );

    \I__10502\ : Span4Mux_v
    port map (
            O => \N__44315\,
            I => \N__44299\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__44310\,
            I => \N__44299\
        );

    \I__10500\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44296\
        );

    \I__10499\ : Span4Mux_v
    port map (
            O => \N__44304\,
            I => \N__44291\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__44299\,
            I => \N__44291\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__44296\,
            I => data_out_frame2_8_1
        );

    \I__10496\ : Odrv4
    port map (
            O => \N__44291\,
            I => data_out_frame2_8_1
        );

    \I__10495\ : InMux
    port map (
            O => \N__44286\,
            I => \N__44281\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__44285\,
            I => \N__44278\
        );

    \I__10493\ : InMux
    port map (
            O => \N__44284\,
            I => \N__44275\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__44281\,
            I => \N__44272\
        );

    \I__10491\ : InMux
    port map (
            O => \N__44278\,
            I => \N__44269\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44264\
        );

    \I__10489\ : Span4Mux_s2_v
    port map (
            O => \N__44272\,
            I => \N__44261\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__44269\,
            I => \N__44258\
        );

    \I__10487\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44255\
        );

    \I__10486\ : InMux
    port map (
            O => \N__44267\,
            I => \N__44252\
        );

    \I__10485\ : Span4Mux_s2_v
    port map (
            O => \N__44264\,
            I => \N__44249\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__44261\,
            I => \N__44244\
        );

    \I__10483\ : Span4Mux_h
    port map (
            O => \N__44258\,
            I => \N__44244\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__44255\,
            I => \N__44241\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__44252\,
            I => data_out_frame2_12_7
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__44249\,
            I => data_out_frame2_12_7
        );

    \I__10479\ : Odrv4
    port map (
            O => \N__44244\,
            I => data_out_frame2_12_7
        );

    \I__10478\ : Odrv12
    port map (
            O => \N__44241\,
            I => data_out_frame2_12_7
        );

    \I__10477\ : InMux
    port map (
            O => \N__44232\,
            I => \N__44225\
        );

    \I__10476\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44222\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44219\
        );

    \I__10474\ : InMux
    port map (
            O => \N__44229\,
            I => \N__44216\
        );

    \I__10473\ : CascadeMux
    port map (
            O => \N__44228\,
            I => \N__44213\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__44225\,
            I => \N__44210\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44207\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__44219\,
            I => \N__44204\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__44216\,
            I => \N__44200\
        );

    \I__10468\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44197\
        );

    \I__10467\ : Span4Mux_v
    port map (
            O => \N__44210\,
            I => \N__44194\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__44207\,
            I => \N__44189\
        );

    \I__10465\ : Span4Mux_h
    port map (
            O => \N__44204\,
            I => \N__44189\
        );

    \I__10464\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44186\
        );

    \I__10463\ : Span12Mux_h
    port map (
            O => \N__44200\,
            I => \N__44181\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__44197\,
            I => \N__44181\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__44194\,
            I => rand_data_5
        );

    \I__10460\ : Odrv4
    port map (
            O => \N__44189\,
            I => rand_data_5
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__44186\,
            I => rand_data_5
        );

    \I__10458\ : Odrv12
    port map (
            O => \N__44181\,
            I => rand_data_5
        );

    \I__10457\ : CascadeMux
    port map (
            O => \N__44172\,
            I => \N__44168\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__44171\,
            I => \N__44164\
        );

    \I__10455\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44161\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44157\
        );

    \I__10453\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44154\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44161\,
            I => \N__44151\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44147\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44144\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__44154\,
            I => \N__44141\
        );

    \I__10448\ : Span4Mux_h
    port map (
            O => \N__44151\,
            I => \N__44137\
        );

    \I__10447\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44134\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__44147\,
            I => \N__44131\
        );

    \I__10445\ : Span4Mux_s3_v
    port map (
            O => \N__44144\,
            I => \N__44126\
        );

    \I__10444\ : Span4Mux_s3_v
    port map (
            O => \N__44141\,
            I => \N__44126\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44123\
        );

    \I__10442\ : Span4Mux_h
    port map (
            O => \N__44137\,
            I => \N__44120\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__44134\,
            I => \N__44117\
        );

    \I__10440\ : Span4Mux_s3_v
    port map (
            O => \N__44131\,
            I => \N__44112\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__44126\,
            I => \N__44112\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__44123\,
            I => data_out_frame2_12_5
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__44120\,
            I => data_out_frame2_12_5
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__44117\,
            I => data_out_frame2_12_5
        );

    \I__10435\ : Odrv4
    port map (
            O => \N__44112\,
            I => data_out_frame2_12_5
        );

    \I__10434\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44100\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__44100\,
            I => \N__44096\
        );

    \I__10432\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44093\
        );

    \I__10431\ : Span4Mux_v
    port map (
            O => \N__44096\,
            I => \N__44088\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__44093\,
            I => \N__44088\
        );

    \I__10429\ : Span4Mux_h
    port map (
            O => \N__44088\,
            I => \N__44083\
        );

    \I__10428\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44080\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44077\
        );

    \I__10426\ : Span4Mux_v
    port map (
            O => \N__44083\,
            I => \N__44074\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__44080\,
            I => data_out_frame2_6_3
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__44077\,
            I => data_out_frame2_6_3
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__44074\,
            I => data_out_frame2_6_3
        );

    \I__10422\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44064\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__44064\,
            I => \c0.n5_adj_2381\
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__44061\,
            I => \N__44058\
        );

    \I__10419\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44054\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44050\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__44054\,
            I => \N__44047\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44053\,
            I => \N__44044\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44050\,
            I => \N__44041\
        );

    \I__10414\ : Span4Mux_v
    port map (
            O => \N__44047\,
            I => \N__44037\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__44044\,
            I => \N__44034\
        );

    \I__10412\ : Span4Mux_h
    port map (
            O => \N__44041\,
            I => \N__44031\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44040\,
            I => \N__44028\
        );

    \I__10410\ : Span4Mux_h
    port map (
            O => \N__44037\,
            I => \N__44025\
        );

    \I__10409\ : Span4Mux_v
    port map (
            O => \N__44034\,
            I => \N__44022\
        );

    \I__10408\ : Span4Mux_h
    port map (
            O => \N__44031\,
            I => \N__44019\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__44028\,
            I => data_out_frame2_6_1
        );

    \I__10406\ : Odrv4
    port map (
            O => \N__44025\,
            I => data_out_frame2_6_1
        );

    \I__10405\ : Odrv4
    port map (
            O => \N__44022\,
            I => data_out_frame2_6_1
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__44019\,
            I => data_out_frame2_6_1
        );

    \I__10403\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44007\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44007\,
            I => \N__44004\
        );

    \I__10401\ : Span4Mux_s2_v
    port map (
            O => \N__44004\,
            I => \N__44001\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__44001\,
            I => \c0.n30_adj_2434\
        );

    \I__10399\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__43995\,
            I => \c0.data_out_frame2_20_2\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__43992\,
            I => \c0.n18636_cascade_\
        );

    \I__10396\ : InMux
    port map (
            O => \N__43989\,
            I => \N__43986\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__43986\,
            I => \c0.n22_adj_2268\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__43983\,
            I => \N__43980\
        );

    \I__10393\ : InMux
    port map (
            O => \N__43980\,
            I => \N__43976\
        );

    \I__10392\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43973\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__43976\,
            I => \N__43970\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__43973\,
            I => \N__43967\
        );

    \I__10389\ : Span4Mux_s2_v
    port map (
            O => \N__43970\,
            I => \N__43964\
        );

    \I__10388\ : Odrv12
    port map (
            O => \N__43967\,
            I => \c0.n17892\
        );

    \I__10387\ : Odrv4
    port map (
            O => \N__43964\,
            I => \c0.n17892\
        );

    \I__10386\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43955\
        );

    \I__10385\ : CascadeMux
    port map (
            O => \N__43958\,
            I => \N__43951\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__43955\,
            I => \N__43946\
        );

    \I__10383\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43943\
        );

    \I__10382\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43940\
        );

    \I__10381\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43937\
        );

    \I__10380\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43934\
        );

    \I__10379\ : Span4Mux_s2_v
    port map (
            O => \N__43946\,
            I => \N__43931\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__43943\,
            I => \N__43928\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__43940\,
            I => \N__43925\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__43937\,
            I => \N__43922\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__43934\,
            I => data_out_frame2_9_1
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__43931\,
            I => data_out_frame2_9_1
        );

    \I__10373\ : Odrv12
    port map (
            O => \N__43928\,
            I => data_out_frame2_9_1
        );

    \I__10372\ : Odrv4
    port map (
            O => \N__43925\,
            I => data_out_frame2_9_1
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__43922\,
            I => data_out_frame2_9_1
        );

    \I__10370\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43908\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__43908\,
            I => \N__43905\
        );

    \I__10368\ : Odrv12
    port map (
            O => \N__43905\,
            I => \c0.n10893\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__43902\,
            I => \c0.n20_adj_2438_cascade_\
        );

    \I__10366\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43896\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__43893\,
            I => \N__43889\
        );

    \I__10363\ : InMux
    port map (
            O => \N__43892\,
            I => \N__43886\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__43889\,
            I => \c0.n17755\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__43886\,
            I => \c0.n17755\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__10359\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43875\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__43875\,
            I => \N__43872\
        );

    \I__10357\ : Span4Mux_v
    port map (
            O => \N__43872\,
            I => \N__43869\
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__43869\,
            I => \c0.data_out_frame2_19_6\
        );

    \I__10355\ : InMux
    port map (
            O => \N__43866\,
            I => \N__43862\
        );

    \I__10354\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43859\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43852\
        );

    \I__10351\ : Span4Mux_v
    port map (
            O => \N__43856\,
            I => \N__43849\
        );

    \I__10350\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43846\
        );

    \I__10349\ : Span4Mux_v
    port map (
            O => \N__43852\,
            I => \N__43842\
        );

    \I__10348\ : Sp12to4
    port map (
            O => \N__43849\,
            I => \N__43837\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__43846\,
            I => \N__43837\
        );

    \I__10346\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43834\
        );

    \I__10345\ : Span4Mux_v
    port map (
            O => \N__43842\,
            I => \N__43831\
        );

    \I__10344\ : Span12Mux_h
    port map (
            O => \N__43837\,
            I => \N__43828\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__43834\,
            I => data_out_frame2_5_3
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__43831\,
            I => data_out_frame2_5_3
        );

    \I__10341\ : Odrv12
    port map (
            O => \N__43828\,
            I => data_out_frame2_5_3
        );

    \I__10340\ : CascadeMux
    port map (
            O => \N__43821\,
            I => \N__43815\
        );

    \I__10339\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43812\
        );

    \I__10338\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43807\
        );

    \I__10337\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43807\
        );

    \I__10336\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43804\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__43812\,
            I => \N__43801\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43798\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43794\
        );

    \I__10332\ : Span4Mux_h
    port map (
            O => \N__43801\,
            I => \N__43789\
        );

    \I__10331\ : Span4Mux_h
    port map (
            O => \N__43798\,
            I => \N__43789\
        );

    \I__10330\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43786\
        );

    \I__10329\ : Span4Mux_h
    port map (
            O => \N__43794\,
            I => \N__43781\
        );

    \I__10328\ : Span4Mux_v
    port map (
            O => \N__43789\,
            I => \N__43781\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__43786\,
            I => data_out_frame2_12_3
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__43781\,
            I => data_out_frame2_12_3
        );

    \I__10325\ : InMux
    port map (
            O => \N__43776\,
            I => \N__43773\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__43773\,
            I => \c0.n10905\
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__43770\,
            I => \c0.n10905_cascade_\
        );

    \I__10322\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43764\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__43764\,
            I => \c0.n16_adj_2391\
        );

    \I__10320\ : InMux
    port map (
            O => \N__43761\,
            I => \N__43756\
        );

    \I__10319\ : InMux
    port map (
            O => \N__43760\,
            I => \N__43753\
        );

    \I__10318\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43749\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__43756\,
            I => \N__43746\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__43753\,
            I => \N__43742\
        );

    \I__10315\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43739\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__43749\,
            I => \N__43734\
        );

    \I__10313\ : Span4Mux_v
    port map (
            O => \N__43746\,
            I => \N__43734\
        );

    \I__10312\ : InMux
    port map (
            O => \N__43745\,
            I => \N__43731\
        );

    \I__10311\ : Span4Mux_h
    port map (
            O => \N__43742\,
            I => \N__43726\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__43739\,
            I => \N__43726\
        );

    \I__10309\ : Sp12to4
    port map (
            O => \N__43734\,
            I => \N__43723\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__43731\,
            I => \N__43720\
        );

    \I__10307\ : Span4Mux_v
    port map (
            O => \N__43726\,
            I => \N__43717\
        );

    \I__10306\ : Odrv12
    port map (
            O => \N__43723\,
            I => data_out_frame2_8_2
        );

    \I__10305\ : Odrv4
    port map (
            O => \N__43720\,
            I => data_out_frame2_8_2
        );

    \I__10304\ : Odrv4
    port map (
            O => \N__43717\,
            I => data_out_frame2_8_2
        );

    \I__10303\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43703\
        );

    \I__10302\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43703\
        );

    \I__10301\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43700\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__43703\,
            I => \N__43696\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__43700\,
            I => \N__43693\
        );

    \I__10298\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43690\
        );

    \I__10297\ : Span4Mux_h
    port map (
            O => \N__43696\,
            I => \N__43685\
        );

    \I__10296\ : Span4Mux_s1_v
    port map (
            O => \N__43693\,
            I => \N__43685\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__43690\,
            I => data_out_frame2_14_6
        );

    \I__10294\ : Odrv4
    port map (
            O => \N__43685\,
            I => data_out_frame2_14_6
        );

    \I__10293\ : InMux
    port map (
            O => \N__43680\,
            I => \N__43676\
        );

    \I__10292\ : CascadeMux
    port map (
            O => \N__43679\,
            I => \N__43672\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43669\
        );

    \I__10290\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43666\
        );

    \I__10289\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43663\
        );

    \I__10288\ : Span4Mux_h
    port map (
            O => \N__43669\,
            I => \N__43657\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__43666\,
            I => \N__43650\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__43663\,
            I => \N__43650\
        );

    \I__10285\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43645\
        );

    \I__10284\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43645\
        );

    \I__10283\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43642\
        );

    \I__10282\ : Span4Mux_h
    port map (
            O => \N__43657\,
            I => \N__43639\
        );

    \I__10281\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43636\
        );

    \I__10280\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43633\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__43650\,
            I => \N__43630\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__43645\,
            I => \N__43627\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__43642\,
            I => data_out_frame2_11_7
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__43639\,
            I => data_out_frame2_11_7
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__43636\,
            I => data_out_frame2_11_7
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__43633\,
            I => data_out_frame2_11_7
        );

    \I__10273\ : Odrv4
    port map (
            O => \N__43630\,
            I => data_out_frame2_11_7
        );

    \I__10272\ : Odrv4
    port map (
            O => \N__43627\,
            I => data_out_frame2_11_7
        );

    \I__10271\ : InMux
    port map (
            O => \N__43614\,
            I => \N__43611\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43607\
        );

    \I__10269\ : InMux
    port map (
            O => \N__43610\,
            I => \N__43604\
        );

    \I__10268\ : Span4Mux_h
    port map (
            O => \N__43607\,
            I => \N__43599\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__43604\,
            I => \N__43596\
        );

    \I__10266\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43591\
        );

    \I__10265\ : InMux
    port map (
            O => \N__43602\,
            I => \N__43591\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__43599\,
            I => data_out_frame2_14_5
        );

    \I__10263\ : Odrv4
    port map (
            O => \N__43596\,
            I => data_out_frame2_14_5
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__43591\,
            I => data_out_frame2_14_5
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__43584\,
            I => \N__43580\
        );

    \I__10260\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43576\
        );

    \I__10259\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43571\
        );

    \I__10258\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43568\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__43576\,
            I => \N__43565\
        );

    \I__10256\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43562\
        );

    \I__10255\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43559\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__43571\,
            I => \N__43556\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__43568\,
            I => data_out_frame2_12_6
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__43565\,
            I => data_out_frame2_12_6
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__43562\,
            I => data_out_frame2_12_6
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__43559\,
            I => data_out_frame2_12_6
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__43556\,
            I => data_out_frame2_12_6
        );

    \I__10248\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43541\
        );

    \I__10247\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43538\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__43541\,
            I => rand_setpoint_31
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__43538\,
            I => rand_setpoint_31
        );

    \I__10244\ : CascadeMux
    port map (
            O => \N__43533\,
            I => \N__43530\
        );

    \I__10243\ : InMux
    port map (
            O => \N__43530\,
            I => \N__43524\
        );

    \I__10242\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43521\
        );

    \I__10241\ : InMux
    port map (
            O => \N__43528\,
            I => \N__43518\
        );

    \I__10240\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43515\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__43524\,
            I => \N__43511\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43508\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__43518\,
            I => \N__43505\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__43515\,
            I => \N__43502\
        );

    \I__10235\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43499\
        );

    \I__10234\ : Span4Mux_h
    port map (
            O => \N__43511\,
            I => \N__43494\
        );

    \I__10233\ : Span4Mux_v
    port map (
            O => \N__43508\,
            I => \N__43494\
        );

    \I__10232\ : Span4Mux_h
    port map (
            O => \N__43505\,
            I => \N__43491\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__43502\,
            I => \N__43488\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__43499\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__43494\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10228\ : Odrv4
    port map (
            O => \N__43491\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__43488\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__10226\ : SRMux
    port map (
            O => \N__43479\,
            I => \N__43474\
        );

    \I__10225\ : SRMux
    port map (
            O => \N__43478\,
            I => \N__43471\
        );

    \I__10224\ : SRMux
    port map (
            O => \N__43477\,
            I => \N__43468\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__43474\,
            I => \N__43463\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__43471\,
            I => \N__43463\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__43468\,
            I => \N__43459\
        );

    \I__10220\ : Span4Mux_h
    port map (
            O => \N__43463\,
            I => \N__43456\
        );

    \I__10219\ : SRMux
    port map (
            O => \N__43462\,
            I => \N__43453\
        );

    \I__10218\ : Span4Mux_v
    port map (
            O => \N__43459\,
            I => \N__43450\
        );

    \I__10217\ : Span4Mux_h
    port map (
            O => \N__43456\,
            I => \N__43447\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__43453\,
            I => \N__43444\
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__43450\,
            I => \c0.n11277\
        );

    \I__10214\ : Odrv4
    port map (
            O => \N__43447\,
            I => \c0.n11277\
        );

    \I__10213\ : Odrv12
    port map (
            O => \N__43444\,
            I => \c0.n11277\
        );

    \I__10212\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43434\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__43434\,
            I => \N__43431\
        );

    \I__10210\ : Span4Mux_h
    port map (
            O => \N__43431\,
            I => \N__43428\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__43428\,
            I => \c0.data_out_1_1\
        );

    \I__10208\ : CEMux
    port map (
            O => \N__43425\,
            I => \N__43420\
        );

    \I__10207\ : CEMux
    port map (
            O => \N__43424\,
            I => \N__43414\
        );

    \I__10206\ : CEMux
    port map (
            O => \N__43423\,
            I => \N__43406\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__43420\,
            I => \N__43403\
        );

    \I__10204\ : CEMux
    port map (
            O => \N__43419\,
            I => \N__43400\
        );

    \I__10203\ : CEMux
    port map (
            O => \N__43418\,
            I => \N__43397\
        );

    \I__10202\ : CEMux
    port map (
            O => \N__43417\,
            I => \N__43390\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43387\
        );

    \I__10200\ : CEMux
    port map (
            O => \N__43413\,
            I => \N__43384\
        );

    \I__10199\ : InMux
    port map (
            O => \N__43412\,
            I => \N__43377\
        );

    \I__10198\ : InMux
    port map (
            O => \N__43411\,
            I => \N__43377\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__43410\,
            I => \N__43373\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__43409\,
            I => \N__43369\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43365\
        );

    \I__10194\ : Span4Mux_v
    port map (
            O => \N__43403\,
            I => \N__43362\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__43400\,
            I => \N__43357\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43357\
        );

    \I__10191\ : CEMux
    port map (
            O => \N__43396\,
            I => \N__43354\
        );

    \I__10190\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43351\
        );

    \I__10189\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43348\
        );

    \I__10188\ : CascadeMux
    port map (
            O => \N__43393\,
            I => \N__43343\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__43390\,
            I => \N__43336\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__43387\,
            I => \N__43336\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43336\
        );

    \I__10184\ : CEMux
    port map (
            O => \N__43383\,
            I => \N__43333\
        );

    \I__10183\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43330\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__43377\,
            I => \N__43327\
        );

    \I__10181\ : InMux
    port map (
            O => \N__43376\,
            I => \N__43320\
        );

    \I__10180\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43320\
        );

    \I__10179\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43320\
        );

    \I__10178\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43314\
        );

    \I__10177\ : InMux
    port map (
            O => \N__43368\,
            I => \N__43311\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__43365\,
            I => \N__43308\
        );

    \I__10175\ : Span4Mux_v
    port map (
            O => \N__43362\,
            I => \N__43301\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__43357\,
            I => \N__43301\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__43354\,
            I => \N__43301\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__43351\,
            I => \N__43296\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__43348\,
            I => \N__43296\
        );

    \I__10170\ : InMux
    port map (
            O => \N__43347\,
            I => \N__43293\
        );

    \I__10169\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43290\
        );

    \I__10168\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43287\
        );

    \I__10167\ : Span4Mux_h
    port map (
            O => \N__43336\,
            I => \N__43282\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43282\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43279\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__43327\,
            I => \N__43274\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__43320\,
            I => \N__43274\
        );

    \I__10162\ : InMux
    port map (
            O => \N__43319\,
            I => \N__43271\
        );

    \I__10161\ : CascadeMux
    port map (
            O => \N__43318\,
            I => \N__43266\
        );

    \I__10160\ : CascadeMux
    port map (
            O => \N__43317\,
            I => \N__43261\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__43314\,
            I => \N__43254\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N__43254\
        );

    \I__10157\ : Span4Mux_h
    port map (
            O => \N__43308\,
            I => \N__43249\
        );

    \I__10156\ : Span4Mux_h
    port map (
            O => \N__43301\,
            I => \N__43249\
        );

    \I__10155\ : Span4Mux_h
    port map (
            O => \N__43296\,
            I => \N__43244\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43244\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43239\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__43287\,
            I => \N__43239\
        );

    \I__10151\ : Span4Mux_v
    port map (
            O => \N__43282\,
            I => \N__43230\
        );

    \I__10150\ : Span4Mux_v
    port map (
            O => \N__43279\,
            I => \N__43230\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__43274\,
            I => \N__43230\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43230\
        );

    \I__10147\ : InMux
    port map (
            O => \N__43270\,
            I => \N__43227\
        );

    \I__10146\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43222\
        );

    \I__10145\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43222\
        );

    \I__10144\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43217\
        );

    \I__10143\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43217\
        );

    \I__10142\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43212\
        );

    \I__10141\ : InMux
    port map (
            O => \N__43260\,
            I => \N__43212\
        );

    \I__10140\ : InMux
    port map (
            O => \N__43259\,
            I => \N__43209\
        );

    \I__10139\ : Span4Mux_h
    port map (
            O => \N__43254\,
            I => \N__43206\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__43249\,
            I => n11017
        );

    \I__10137\ : Odrv4
    port map (
            O => \N__43244\,
            I => n11017
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__43239\,
            I => n11017
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__43230\,
            I => n11017
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__43227\,
            I => n11017
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__43222\,
            I => n11017
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__43217\,
            I => n11017
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__43212\,
            I => n11017
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__43209\,
            I => n11017
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__43206\,
            I => n11017
        );

    \I__10128\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43179\
        );

    \I__10126\ : Odrv4
    port map (
            O => \N__43179\,
            I => \c0.n18250\
        );

    \I__10125\ : CascadeMux
    port map (
            O => \N__43176\,
            I => \N__43173\
        );

    \I__10124\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__43170\,
            I => \N__43166\
        );

    \I__10122\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \N__43163\
        );

    \I__10121\ : Span4Mux_v
    port map (
            O => \N__43166\,
            I => \N__43160\
        );

    \I__10120\ : InMux
    port map (
            O => \N__43163\,
            I => \N__43157\
        );

    \I__10119\ : Odrv4
    port map (
            O => \N__43160\,
            I => rand_setpoint_8
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43157\,
            I => rand_setpoint_8
        );

    \I__10117\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43149\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__43149\,
            I => \N__43144\
        );

    \I__10115\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43141\
        );

    \I__10114\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43138\
        );

    \I__10113\ : Span4Mux_v
    port map (
            O => \N__43144\,
            I => \N__43133\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__43141\,
            I => \N__43133\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__43138\,
            I => \N__43130\
        );

    \I__10110\ : Span4Mux_h
    port map (
            O => \N__43133\,
            I => \N__43127\
        );

    \I__10109\ : Odrv12
    port map (
            O => \N__43130\,
            I => \c0.data_out_7_0\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__43127\,
            I => \c0.data_out_7_0\
        );

    \I__10107\ : InMux
    port map (
            O => \N__43122\,
            I => \N__43119\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__10105\ : Odrv4
    port map (
            O => \N__43116\,
            I => \c0.n18648\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__43113\,
            I => \N__43110\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__43107\,
            I => \N__43104\
        );

    \I__10101\ : Odrv12
    port map (
            O => \N__43104\,
            I => \c0.n18642\
        );

    \I__10100\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43098\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43095\
        );

    \I__10098\ : Span4Mux_h
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__43092\,
            I => \c0.n18221\
        );

    \I__10096\ : CascadeMux
    port map (
            O => \N__43089\,
            I => \c0.n18765_cascade_\
        );

    \I__10095\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43083\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__43083\,
            I => \N__43080\
        );

    \I__10093\ : Odrv4
    port map (
            O => \N__43080\,
            I => \c0.n6_adj_2227\
        );

    \I__10092\ : CascadeMux
    port map (
            O => \N__43077\,
            I => \c0.n18768_cascade_\
        );

    \I__10091\ : InMux
    port map (
            O => \N__43074\,
            I => \N__43071\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__43071\,
            I => \N__43068\
        );

    \I__10089\ : Span4Mux_h
    port map (
            O => \N__43068\,
            I => \N__43065\
        );

    \I__10088\ : Span4Mux_h
    port map (
            O => \N__43065\,
            I => \N__43062\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__43062\,
            I => \N__43059\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__43059\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__10085\ : InMux
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__43053\,
            I => \N__43049\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43052\,
            I => \N__43046\
        );

    \I__10082\ : Span4Mux_s2_v
    port map (
            O => \N__43049\,
            I => \N__43043\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__43046\,
            I => data_out_frame2_18_2
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__43043\,
            I => data_out_frame2_18_2
        );

    \I__10079\ : CascadeMux
    port map (
            O => \N__43038\,
            I => \N__43035\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43035\,
            I => \N__43032\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__43032\,
            I => \N__43029\
        );

    \I__10076\ : Odrv12
    port map (
            O => \N__43029\,
            I => \c0.data_out_frame2_19_2\
        );

    \I__10075\ : InMux
    port map (
            O => \N__43026\,
            I => \N__43023\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__10073\ : Sp12to4
    port map (
            O => \N__43020\,
            I => \N__43016\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43013\
        );

    \I__10071\ : Span12Mux_s2_v
    port map (
            O => \N__43016\,
            I => \N__43010\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__43013\,
            I => data_out_frame2_17_2
        );

    \I__10069\ : Odrv12
    port map (
            O => \N__43010\,
            I => data_out_frame2_17_2
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__43005\,
            I => \c0.n18633_cascade_\
        );

    \I__10067\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__42999\,
            I => \c0.n18780\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__42996\,
            I => \c0.n22_adj_2240_cascade_\
        );

    \I__10064\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42990\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42987\
        );

    \I__10062\ : Span12Mux_s5_h
    port map (
            O => \N__42987\,
            I => \N__42984\
        );

    \I__10061\ : Odrv12
    port map (
            O => \N__42984\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__42981\,
            I => \c0.n18783_cascade_\
        );

    \I__10059\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42973\
        );

    \I__10058\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42970\
        );

    \I__10057\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42966\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__42973\,
            I => \N__42963\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__42970\,
            I => \N__42960\
        );

    \I__10054\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42957\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__42966\,
            I => \N__42952\
        );

    \I__10052\ : Span12Mux_h
    port map (
            O => \N__42963\,
            I => \N__42952\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__42960\,
            I => \N__42949\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__42957\,
            I => data_out_frame2_13_4
        );

    \I__10049\ : Odrv12
    port map (
            O => \N__42952\,
            I => data_out_frame2_13_4
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__42949\,
            I => data_out_frame2_13_4
        );

    \I__10047\ : InMux
    port map (
            O => \N__42942\,
            I => \N__42938\
        );

    \I__10046\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42934\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__42938\,
            I => \N__42930\
        );

    \I__10044\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42926\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__42934\,
            I => \N__42923\
        );

    \I__10042\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42920\
        );

    \I__10041\ : Span4Mux_v
    port map (
            O => \N__42930\,
            I => \N__42917\
        );

    \I__10040\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42914\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__42926\,
            I => \N__42911\
        );

    \I__10038\ : Span4Mux_h
    port map (
            O => \N__42923\,
            I => \N__42906\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__42920\,
            I => \N__42906\
        );

    \I__10036\ : Odrv4
    port map (
            O => \N__42917\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__42914\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__42911\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__42906\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__10032\ : InMux
    port map (
            O => \N__42897\,
            I => \N__42894\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__42894\,
            I => \N__42891\
        );

    \I__10030\ : Odrv12
    port map (
            O => \N__42891\,
            I => \c0.n18311\
        );

    \I__10029\ : CascadeMux
    port map (
            O => \N__42888\,
            I => \N__42884\
        );

    \I__10028\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42881\
        );

    \I__10027\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42878\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__42881\,
            I => rand_setpoint_11
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__42878\,
            I => rand_setpoint_11
        );

    \I__10024\ : InMux
    port map (
            O => \N__42873\,
            I => \N__42852\
        );

    \I__10023\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42852\
        );

    \I__10022\ : InMux
    port map (
            O => \N__42871\,
            I => \N__42843\
        );

    \I__10021\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42843\
        );

    \I__10020\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42843\
        );

    \I__10019\ : InMux
    port map (
            O => \N__42868\,
            I => \N__42843\
        );

    \I__10018\ : InMux
    port map (
            O => \N__42867\,
            I => \N__42836\
        );

    \I__10017\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42836\
        );

    \I__10016\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42836\
        );

    \I__10015\ : InMux
    port map (
            O => \N__42864\,
            I => \N__42831\
        );

    \I__10014\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42831\
        );

    \I__10013\ : InMux
    port map (
            O => \N__42862\,
            I => \N__42827\
        );

    \I__10012\ : InMux
    port map (
            O => \N__42861\,
            I => \N__42824\
        );

    \I__10011\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42805\
        );

    \I__10010\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42792\
        );

    \I__10009\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42792\
        );

    \I__10008\ : InMux
    port map (
            O => \N__42857\,
            I => \N__42789\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__42852\,
            I => \N__42782\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__42843\,
            I => \N__42782\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__42836\,
            I => \N__42782\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__42831\,
            I => \N__42776\
        );

    \I__10003\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42773\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42770\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__42824\,
            I => \N__42767\
        );

    \I__10000\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42758\
        );

    \I__9999\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42758\
        );

    \I__9998\ : InMux
    port map (
            O => \N__42821\,
            I => \N__42758\
        );

    \I__9997\ : InMux
    port map (
            O => \N__42820\,
            I => \N__42758\
        );

    \I__9996\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42749\
        );

    \I__9995\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42749\
        );

    \I__9994\ : InMux
    port map (
            O => \N__42817\,
            I => \N__42749\
        );

    \I__9993\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42749\
        );

    \I__9992\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42742\
        );

    \I__9991\ : InMux
    port map (
            O => \N__42814\,
            I => \N__42742\
        );

    \I__9990\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42742\
        );

    \I__9989\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42739\
        );

    \I__9988\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42736\
        );

    \I__9987\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42731\
        );

    \I__9986\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42731\
        );

    \I__9985\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42728\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__42805\,
            I => \N__42725\
        );

    \I__9983\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42718\
        );

    \I__9982\ : InMux
    port map (
            O => \N__42803\,
            I => \N__42718\
        );

    \I__9981\ : InMux
    port map (
            O => \N__42802\,
            I => \N__42718\
        );

    \I__9980\ : InMux
    port map (
            O => \N__42801\,
            I => \N__42713\
        );

    \I__9979\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42713\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__42799\,
            I => \N__42709\
        );

    \I__9977\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42704\
        );

    \I__9976\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42701\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42694\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__42789\,
            I => \N__42694\
        );

    \I__9973\ : Span4Mux_v
    port map (
            O => \N__42782\,
            I => \N__42694\
        );

    \I__9972\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42691\
        );

    \I__9971\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42686\
        );

    \I__9970\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42686\
        );

    \I__9969\ : Span4Mux_v
    port map (
            O => \N__42776\,
            I => \N__42683\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__42773\,
            I => \N__42670\
        );

    \I__9967\ : Span4Mux_h
    port map (
            O => \N__42770\,
            I => \N__42670\
        );

    \I__9966\ : Span4Mux_v
    port map (
            O => \N__42767\,
            I => \N__42670\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42670\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__42749\,
            I => \N__42670\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__42742\,
            I => \N__42670\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__42739\,
            I => \N__42655\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__42736\,
            I => \N__42655\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__42731\,
            I => \N__42655\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__42728\,
            I => \N__42655\
        );

    \I__9958\ : Span4Mux_v
    port map (
            O => \N__42725\,
            I => \N__42655\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__42718\,
            I => \N__42655\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__42713\,
            I => \N__42655\
        );

    \I__9955\ : InMux
    port map (
            O => \N__42712\,
            I => \N__42652\
        );

    \I__9954\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42649\
        );

    \I__9953\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42646\
        );

    \I__9952\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42643\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42636\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__42701\,
            I => \N__42636\
        );

    \I__9949\ : Span4Mux_v
    port map (
            O => \N__42694\,
            I => \N__42636\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__42691\,
            I => \N__42627\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__42686\,
            I => \N__42627\
        );

    \I__9946\ : Span4Mux_h
    port map (
            O => \N__42683\,
            I => \N__42627\
        );

    \I__9945\ : Span4Mux_v
    port map (
            O => \N__42670\,
            I => \N__42627\
        );

    \I__9944\ : Sp12to4
    port map (
            O => \N__42655\,
            I => \N__42622\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__42652\,
            I => \N__42622\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__42649\,
            I => \N__42619\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__42646\,
            I => byte_transmit_counter_0
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__42643\,
            I => byte_transmit_counter_0
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__42636\,
            I => byte_transmit_counter_0
        );

    \I__9938\ : Odrv4
    port map (
            O => \N__42627\,
            I => byte_transmit_counter_0
        );

    \I__9937\ : Odrv12
    port map (
            O => \N__42622\,
            I => byte_transmit_counter_0
        );

    \I__9936\ : Odrv4
    port map (
            O => \N__42619\,
            I => byte_transmit_counter_0
        );

    \I__9935\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42601\
        );

    \I__9934\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42597\
        );

    \I__9933\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42594\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__42601\,
            I => \N__42591\
        );

    \I__9931\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42588\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__42597\,
            I => \N__42585\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__42594\,
            I => \N__42582\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__42591\,
            I => \N__42577\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__42588\,
            I => \N__42577\
        );

    \I__9926\ : Span4Mux_h
    port map (
            O => \N__42585\,
            I => \N__42574\
        );

    \I__9925\ : Span4Mux_h
    port map (
            O => \N__42582\,
            I => \N__42571\
        );

    \I__9924\ : Span4Mux_v
    port map (
            O => \N__42577\,
            I => \N__42568\
        );

    \I__9923\ : Odrv4
    port map (
            O => \N__42574\,
            I => \c0.data_out_6_3\
        );

    \I__9922\ : Odrv4
    port map (
            O => \N__42571\,
            I => \c0.data_out_6_3\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__42568\,
            I => \c0.data_out_6_3\
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__42561\,
            I => \N__42558\
        );

    \I__9919\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9917\ : Odrv12
    port map (
            O => \N__42552\,
            I => \c0.n5_adj_2217\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__42549\,
            I => \N__42546\
        );

    \I__9915\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__42543\,
            I => \c0.n18201\
        );

    \I__9913\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42537\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42533\
        );

    \I__9911\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42530\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__42533\,
            I => \N__42525\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__42530\,
            I => \N__42525\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__42525\,
            I => \N__42521\
        );

    \I__9907\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42518\
        );

    \I__9906\ : Odrv4
    port map (
            O => \N__42521\,
            I => \c0.data_out_7_3\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__42518\,
            I => \c0.data_out_7_3\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__42513\,
            I => \N__42509\
        );

    \I__9903\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42506\
        );

    \I__9902\ : InMux
    port map (
            O => \N__42509\,
            I => \N__42503\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__42506\,
            I => rand_setpoint_24
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__42503\,
            I => rand_setpoint_24
        );

    \I__9899\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42495\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__42495\,
            I => \N__42490\
        );

    \I__9897\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42486\
        );

    \I__9896\ : InMux
    port map (
            O => \N__42493\,
            I => \N__42482\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__42490\,
            I => \N__42479\
        );

    \I__9894\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42476\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__42486\,
            I => \N__42473\
        );

    \I__9892\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42470\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__42482\,
            I => \N__42466\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__42479\,
            I => \N__42461\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__42476\,
            I => \N__42461\
        );

    \I__9888\ : Sp12to4
    port map (
            O => \N__42473\,
            I => \N__42456\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__42470\,
            I => \N__42456\
        );

    \I__9886\ : InMux
    port map (
            O => \N__42469\,
            I => \N__42453\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__42466\,
            I => \N__42448\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__42461\,
            I => \N__42448\
        );

    \I__9883\ : Span12Mux_v
    port map (
            O => \N__42456\,
            I => \N__42443\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42443\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__42448\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__9880\ : Odrv12
    port map (
            O => \N__42443\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__9879\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42435\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42432\
        );

    \I__9877\ : Odrv12
    port map (
            O => \N__42432\,
            I => \c0.n18666\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__42429\,
            I => \N__42426\
        );

    \I__9875\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42423\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__42420\,
            I => \c0.n18660\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42414\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__42414\,
            I => \N__42411\
        );

    \I__9870\ : Odrv12
    port map (
            O => \N__42411\,
            I => \c0.n18371\
        );

    \I__9869\ : CascadeMux
    port map (
            O => \N__42408\,
            I => \c0.n18735_cascade_\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__42402\,
            I => \N__42399\
        );

    \I__9866\ : Odrv4
    port map (
            O => \N__42399\,
            I => \c0.n6_adj_2360\
        );

    \I__9865\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42393\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__42393\,
            I => \c0.n22_adj_2259\
        );

    \I__9863\ : CascadeMux
    port map (
            O => \N__42390\,
            I => \c0.n18738_cascade_\
        );

    \I__9862\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__42384\,
            I => \N__42381\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__42378\,
            I => \N__42375\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__42375\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__9857\ : InMux
    port map (
            O => \N__42372\,
            I => \N__42369\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__42369\,
            I => \N__42365\
        );

    \I__9855\ : InMux
    port map (
            O => \N__42368\,
            I => \N__42362\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__42365\,
            I => \N__42359\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__42362\,
            I => data_out_frame2_18_6
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__42359\,
            I => data_out_frame2_18_6
        );

    \I__9851\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42351\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__42351\,
            I => \N__42348\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__42348\,
            I => \c0.n18708\
        );

    \I__9848\ : CascadeMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9847\ : InMux
    port map (
            O => \N__42342\,
            I => \N__42339\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9845\ : Span4Mux_h
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__9843\ : Odrv4
    port map (
            O => \N__42330\,
            I => \c0.n18762\
        );

    \I__9842\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42324\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__42324\,
            I => \N__42321\
        );

    \I__9840\ : Span4Mux_h
    port map (
            O => \N__42321\,
            I => \N__42318\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__42318\,
            I => \c0.n18308\
        );

    \I__9838\ : CascadeMux
    port map (
            O => \N__42315\,
            I => \c0.n18777_cascade_\
        );

    \I__9837\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42309\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__9835\ : Odrv12
    port map (
            O => \N__42306\,
            I => \c0.n6_adj_2218\
        );

    \I__9834\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__42300\,
            I => \c0.n18699\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9831\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42291\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42287\
        );

    \I__9829\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42284\
        );

    \I__9828\ : Span4Mux_h
    port map (
            O => \N__42287\,
            I => \N__42281\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__42284\,
            I => data_out_frame2_17_6
        );

    \I__9826\ : Odrv4
    port map (
            O => \N__42281\,
            I => data_out_frame2_17_6
        );

    \I__9825\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42272\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__42275\,
            I => \N__42269\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__42272\,
            I => \N__42266\
        );

    \I__9822\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42262\
        );

    \I__9821\ : Span4Mux_v
    port map (
            O => \N__42266\,
            I => \N__42258\
        );

    \I__9820\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42255\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__42262\,
            I => \N__42252\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42249\
        );

    \I__9817\ : Span4Mux_v
    port map (
            O => \N__42258\,
            I => \N__42246\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__42255\,
            I => \N__42241\
        );

    \I__9815\ : Span4Mux_s0_v
    port map (
            O => \N__42252\,
            I => \N__42241\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__42249\,
            I => data_out_frame2_16_6
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__42246\,
            I => data_out_frame2_16_6
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__42241\,
            I => data_out_frame2_16_6
        );

    \I__9811\ : CascadeMux
    port map (
            O => \N__42234\,
            I => \c0.n18702_cascade_\
        );

    \I__9810\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42227\
        );

    \I__9809\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42224\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__42227\,
            I => \N__42220\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__42224\,
            I => \N__42217\
        );

    \I__9806\ : InMux
    port map (
            O => \N__42223\,
            I => \N__42214\
        );

    \I__9805\ : Span4Mux_s2_v
    port map (
            O => \N__42220\,
            I => \N__42211\
        );

    \I__9804\ : Span4Mux_h
    port map (
            O => \N__42217\,
            I => \N__42208\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__42214\,
            I => data_out_frame2_13_7
        );

    \I__9802\ : Odrv4
    port map (
            O => \N__42211\,
            I => data_out_frame2_13_7
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__42208\,
            I => data_out_frame2_13_7
        );

    \I__9800\ : InMux
    port map (
            O => \N__42201\,
            I => \N__42198\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__42198\,
            I => \N__42195\
        );

    \I__9798\ : Odrv12
    port map (
            O => \N__42195\,
            I => \c0.n10_adj_2411\
        );

    \I__9797\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42189\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42186\
        );

    \I__9795\ : Span4Mux_v
    port map (
            O => \N__42186\,
            I => \N__42183\
        );

    \I__9794\ : Odrv4
    port map (
            O => \N__42183\,
            I => \c0.n18705\
        );

    \I__9793\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42177\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__42177\,
            I => \N__42174\
        );

    \I__9791\ : Span4Mux_s1_v
    port map (
            O => \N__42174\,
            I => \N__42170\
        );

    \I__9790\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42167\
        );

    \I__9789\ : Span4Mux_v
    port map (
            O => \N__42170\,
            I => \N__42160\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__42167\,
            I => \N__42160\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42166\,
            I => \N__42155\
        );

    \I__9786\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42155\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__42160\,
            I => data_out_frame2_13_6
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__42155\,
            I => data_out_frame2_13_6
        );

    \I__9783\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42145\
        );

    \I__9782\ : InMux
    port map (
            O => \N__42149\,
            I => \N__42142\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__42148\,
            I => \N__42139\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__42145\,
            I => \N__42135\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42142\,
            I => \N__42132\
        );

    \I__9778\ : InMux
    port map (
            O => \N__42139\,
            I => \N__42129\
        );

    \I__9777\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42125\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__42135\,
            I => \N__42122\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__42132\,
            I => \N__42119\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__42129\,
            I => \N__42116\
        );

    \I__9773\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42113\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__42110\
        );

    \I__9771\ : Odrv4
    port map (
            O => \N__42122\,
            I => rand_data_27
        );

    \I__9770\ : Odrv4
    port map (
            O => \N__42119\,
            I => rand_data_27
        );

    \I__9769\ : Odrv4
    port map (
            O => \N__42116\,
            I => rand_data_27
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__42113\,
            I => rand_data_27
        );

    \I__9767\ : Odrv12
    port map (
            O => \N__42110\,
            I => rand_data_27
        );

    \I__9766\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42092\
        );

    \I__9765\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42092\
        );

    \I__9764\ : CascadeMux
    port map (
            O => \N__42097\,
            I => \N__42088\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__42092\,
            I => \N__42084\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42091\,
            I => \N__42081\
        );

    \I__9761\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42077\
        );

    \I__9760\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42074\
        );

    \I__9759\ : Span12Mux_s4_v
    port map (
            O => \N__42084\,
            I => \N__42069\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__42081\,
            I => \N__42069\
        );

    \I__9757\ : InMux
    port map (
            O => \N__42080\,
            I => \N__42066\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42077\,
            I => \N__42063\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42074\,
            I => rand_data_7
        );

    \I__9754\ : Odrv12
    port map (
            O => \N__42069\,
            I => rand_data_7
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__42066\,
            I => rand_data_7
        );

    \I__9752\ : Odrv12
    port map (
            O => \N__42063\,
            I => rand_data_7
        );

    \I__9751\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42049\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42046\
        );

    \I__9749\ : InMux
    port map (
            O => \N__42052\,
            I => \N__42043\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__42049\,
            I => \N__42040\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__42046\,
            I => \N__42036\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__42043\,
            I => \N__42031\
        );

    \I__9745\ : Span4Mux_h
    port map (
            O => \N__42040\,
            I => \N__42031\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42039\,
            I => \N__42028\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__42036\,
            I => \N__42025\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__42031\,
            I => \N__42022\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42028\,
            I => data_out_frame2_13_3
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__42025\,
            I => data_out_frame2_13_3
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__42022\,
            I => data_out_frame2_13_3
        );

    \I__9738\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__42012\,
            I => \N__42009\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__42009\,
            I => \N__42006\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__42006\,
            I => \c0.n18657\
        );

    \I__9734\ : InMux
    port map (
            O => \N__42003\,
            I => \N__42000\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__42000\,
            I => \N__41996\
        );

    \I__9732\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41993\
        );

    \I__9731\ : Span4Mux_h
    port map (
            O => \N__41996\,
            I => \N__41990\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__41993\,
            I => data_out_frame2_18_3
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__41990\,
            I => data_out_frame2_18_3
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__9727\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41979\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__41976\,
            I => \c0.data_out_frame2_19_3\
        );

    \I__9724\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41969\
        );

    \I__9723\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41966\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__41969\,
            I => data_out_frame2_17_3
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__41966\,
            I => data_out_frame2_17_3
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__41961\,
            I => \c0.n18651_cascade_\
        );

    \I__9719\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41951\
        );

    \I__9717\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41947\
        );

    \I__9716\ : Span4Mux_h
    port map (
            O => \N__41951\,
            I => \N__41943\
        );

    \I__9715\ : InMux
    port map (
            O => \N__41950\,
            I => \N__41940\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__41947\,
            I => \N__41937\
        );

    \I__9713\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41934\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__41943\,
            I => \N__41931\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41928\
        );

    \I__9710\ : Span4Mux_h
    port map (
            O => \N__41937\,
            I => \N__41925\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__41934\,
            I => data_out_frame2_16_3
        );

    \I__9708\ : Odrv4
    port map (
            O => \N__41931\,
            I => data_out_frame2_16_3
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__41928\,
            I => data_out_frame2_16_3
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__41925\,
            I => data_out_frame2_16_3
        );

    \I__9705\ : InMux
    port map (
            O => \N__41916\,
            I => \N__41913\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__41913\,
            I => \N__41910\
        );

    \I__9703\ : Span4Mux_v
    port map (
            O => \N__41910\,
            I => \N__41907\
        );

    \I__9702\ : Odrv4
    port map (
            O => \N__41907\,
            I => \c0.data_out_frame2_20_3\
        );

    \I__9701\ : CascadeMux
    port map (
            O => \N__41904\,
            I => \c0.n18654_cascade_\
        );

    \I__9700\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__41898\,
            I => \N__41894\
        );

    \I__9698\ : InMux
    port map (
            O => \N__41897\,
            I => \N__41891\
        );

    \I__9697\ : Span4Mux_v
    port map (
            O => \N__41894\,
            I => \N__41888\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__41891\,
            I => \c0.n17880\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__41888\,
            I => \c0.n17880\
        );

    \I__9694\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41879\
        );

    \I__9693\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41876\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__41879\,
            I => \N__41873\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__41876\,
            I => \N__41868\
        );

    \I__9690\ : Span4Mux_s1_v
    port map (
            O => \N__41873\,
            I => \N__41868\
        );

    \I__9689\ : Odrv4
    port map (
            O => \N__41868\,
            I => \c0.n17789\
        );

    \I__9688\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41860\
        );

    \I__9687\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41854\
        );

    \I__9686\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41854\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41850\
        );

    \I__9684\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41847\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__41854\,
            I => \N__41844\
        );

    \I__9682\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41841\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__41850\,
            I => \N__41836\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41836\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__41844\,
            I => \N__41833\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__41841\,
            I => data_out_frame2_5_6
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__41836\,
            I => data_out_frame2_5_6
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__41833\,
            I => data_out_frame2_5_6
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__9674\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41820\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__41820\,
            I => \c0.n5_adj_2439\
        );

    \I__9672\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41812\
        );

    \I__9671\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41808\
        );

    \I__9670\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41805\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__41812\,
            I => \N__41802\
        );

    \I__9668\ : CascadeMux
    port map (
            O => \N__41811\,
            I => \N__41799\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__41808\,
            I => \N__41796\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__41805\,
            I => \N__41793\
        );

    \I__9665\ : Span4Mux_h
    port map (
            O => \N__41802\,
            I => \N__41790\
        );

    \I__9664\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41787\
        );

    \I__9663\ : Span4Mux_h
    port map (
            O => \N__41796\,
            I => \N__41782\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__41793\,
            I => \N__41782\
        );

    \I__9661\ : Span4Mux_h
    port map (
            O => \N__41790\,
            I => \N__41779\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__41787\,
            I => \N__41774\
        );

    \I__9659\ : Sp12to4
    port map (
            O => \N__41782\,
            I => \N__41774\
        );

    \I__9658\ : Span4Mux_h
    port map (
            O => \N__41779\,
            I => \N__41771\
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__41774\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__41771\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__9655\ : InMux
    port map (
            O => \N__41766\,
            I => \N__41760\
        );

    \I__9654\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41755\
        );

    \I__9653\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41755\
        );

    \I__9652\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41752\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__41760\,
            I => \N__41748\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__41755\,
            I => \N__41745\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__41752\,
            I => \N__41742\
        );

    \I__9648\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41739\
        );

    \I__9647\ : Span4Mux_h
    port map (
            O => \N__41748\,
            I => \N__41736\
        );

    \I__9646\ : Span4Mux_h
    port map (
            O => \N__41745\,
            I => \N__41731\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__41742\,
            I => \N__41731\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__41739\,
            I => data_out_frame2_15_6
        );

    \I__9643\ : Odrv4
    port map (
            O => \N__41736\,
            I => data_out_frame2_15_6
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__41731\,
            I => data_out_frame2_15_6
        );

    \I__9641\ : InMux
    port map (
            O => \N__41724\,
            I => \N__41719\
        );

    \I__9640\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41716\
        );

    \I__9639\ : CascadeMux
    port map (
            O => \N__41722\,
            I => \N__41713\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41710\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__41716\,
            I => \N__41707\
        );

    \I__9636\ : InMux
    port map (
            O => \N__41713\,
            I => \N__41704\
        );

    \I__9635\ : Span4Mux_s2_v
    port map (
            O => \N__41710\,
            I => \N__41698\
        );

    \I__9634\ : Span4Mux_v
    port map (
            O => \N__41707\,
            I => \N__41698\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__41704\,
            I => \N__41695\
        );

    \I__9632\ : InMux
    port map (
            O => \N__41703\,
            I => \N__41692\
        );

    \I__9631\ : Span4Mux_h
    port map (
            O => \N__41698\,
            I => \N__41689\
        );

    \I__9630\ : Span4Mux_s3_v
    port map (
            O => \N__41695\,
            I => \N__41686\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__41692\,
            I => data_out_frame2_13_1
        );

    \I__9628\ : Odrv4
    port map (
            O => \N__41689\,
            I => data_out_frame2_13_1
        );

    \I__9627\ : Odrv4
    port map (
            O => \N__41686\,
            I => data_out_frame2_13_1
        );

    \I__9626\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41675\
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__41678\,
            I => \N__41671\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__41675\,
            I => \N__41667\
        );

    \I__9623\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41664\
        );

    \I__9622\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41661\
        );

    \I__9621\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41658\
        );

    \I__9620\ : Span4Mux_h
    port map (
            O => \N__41667\,
            I => \N__41654\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41651\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__41661\,
            I => \N__41648\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41645\
        );

    \I__9616\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41642\
        );

    \I__9615\ : Span4Mux_s1_v
    port map (
            O => \N__41654\,
            I => \N__41639\
        );

    \I__9614\ : Span4Mux_v
    port map (
            O => \N__41651\,
            I => \N__41632\
        );

    \I__9613\ : Span4Mux_v
    port map (
            O => \N__41648\,
            I => \N__41632\
        );

    \I__9612\ : Span4Mux_h
    port map (
            O => \N__41645\,
            I => \N__41632\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__41642\,
            I => data_out_frame2_8_7
        );

    \I__9610\ : Odrv4
    port map (
            O => \N__41639\,
            I => data_out_frame2_8_7
        );

    \I__9609\ : Odrv4
    port map (
            O => \N__41632\,
            I => data_out_frame2_8_7
        );

    \I__9608\ : CascadeMux
    port map (
            O => \N__41625\,
            I => \N__41621\
        );

    \I__9607\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41617\
        );

    \I__9606\ : InMux
    port map (
            O => \N__41621\,
            I => \N__41614\
        );

    \I__9605\ : InMux
    port map (
            O => \N__41620\,
            I => \N__41610\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__41617\,
            I => \N__41607\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__41614\,
            I => \N__41604\
        );

    \I__9602\ : CascadeMux
    port map (
            O => \N__41613\,
            I => \N__41601\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__41610\,
            I => \N__41598\
        );

    \I__9600\ : Span4Mux_v
    port map (
            O => \N__41607\,
            I => \N__41593\
        );

    \I__9599\ : Span4Mux_h
    port map (
            O => \N__41604\,
            I => \N__41593\
        );

    \I__9598\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41590\
        );

    \I__9597\ : Span12Mux_h
    port map (
            O => \N__41598\,
            I => \N__41587\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__41593\,
            I => \N__41584\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__41590\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9594\ : Odrv12
    port map (
            O => \N__41587\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__41584\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9592\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41574\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__41574\,
            I => \N__41571\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__41571\,
            I => \c0.n10_adj_2431\
        );

    \I__9589\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41561\
        );

    \I__9588\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41556\
        );

    \I__9587\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41556\
        );

    \I__9586\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41552\
        );

    \I__9585\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41549\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__41561\,
            I => \N__41546\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__41556\,
            I => \N__41543\
        );

    \I__9582\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41540\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__41552\,
            I => \N__41537\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__41549\,
            I => \N__41530\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__41546\,
            I => \N__41530\
        );

    \I__9578\ : Span4Mux_h
    port map (
            O => \N__41543\,
            I => \N__41530\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41540\,
            I => data_out_frame2_5_2
        );

    \I__9576\ : Odrv4
    port map (
            O => \N__41537\,
            I => data_out_frame2_5_2
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__41530\,
            I => data_out_frame2_5_2
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__9573\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41517\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__9571\ : Sp12to4
    port map (
            O => \N__41514\,
            I => \N__41511\
        );

    \I__9570\ : Odrv12
    port map (
            O => \N__41511\,
            I => \c0.n17865\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__41508\,
            I => \N__41504\
        );

    \I__9568\ : InMux
    port map (
            O => \N__41507\,
            I => \N__41501\
        );

    \I__9567\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41496\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__41501\,
            I => \N__41493\
        );

    \I__9565\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41490\
        );

    \I__9564\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41487\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__41496\,
            I => \N__41484\
        );

    \I__9562\ : Span4Mux_v
    port map (
            O => \N__41493\,
            I => \N__41479\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41479\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__41487\,
            I => \N__41475\
        );

    \I__9559\ : Span4Mux_v
    port map (
            O => \N__41484\,
            I => \N__41472\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__41479\,
            I => \N__41469\
        );

    \I__9557\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41466\
        );

    \I__9556\ : Span4Mux_v
    port map (
            O => \N__41475\,
            I => \N__41463\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__41472\,
            I => rand_data_28
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__41469\,
            I => rand_data_28
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__41466\,
            I => rand_data_28
        );

    \I__9552\ : Odrv4
    port map (
            O => \N__41463\,
            I => rand_data_28
        );

    \I__9551\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41448\
        );

    \I__9550\ : InMux
    port map (
            O => \N__41453\,
            I => \N__41443\
        );

    \I__9549\ : InMux
    port map (
            O => \N__41452\,
            I => \N__41438\
        );

    \I__9548\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41438\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41435\
        );

    \I__9546\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41432\
        );

    \I__9545\ : InMux
    port map (
            O => \N__41446\,
            I => \N__41429\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__41443\,
            I => \N__41426\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__41438\,
            I => rand_data_11
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__41435\,
            I => rand_data_11
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__41432\,
            I => rand_data_11
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__41429\,
            I => rand_data_11
        );

    \I__9539\ : Odrv12
    port map (
            O => \N__41426\,
            I => rand_data_11
        );

    \I__9538\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41410\
        );

    \I__9537\ : InMux
    port map (
            O => \N__41414\,
            I => \N__41407\
        );

    \I__9536\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41402\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__41410\,
            I => \N__41399\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41407\,
            I => \N__41396\
        );

    \I__9533\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41393\
        );

    \I__9532\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41390\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__41402\,
            I => \N__41383\
        );

    \I__9530\ : Span4Mux_s3_v
    port map (
            O => \N__41399\,
            I => \N__41383\
        );

    \I__9529\ : Span4Mux_h
    port map (
            O => \N__41396\,
            I => \N__41383\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__41393\,
            I => data_out_frame2_10_3
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__41390\,
            I => data_out_frame2_10_3
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__41383\,
            I => data_out_frame2_10_3
        );

    \I__9525\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41373\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__41373\,
            I => \c0.n18663\
        );

    \I__9523\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41367\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41361\
        );

    \I__9521\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41358\
        );

    \I__9520\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41354\
        );

    \I__9519\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41351\
        );

    \I__9518\ : Span12Mux_s7_v
    port map (
            O => \N__41361\,
            I => \N__41348\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__41358\,
            I => \N__41345\
        );

    \I__9516\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41342\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__41354\,
            I => data_out_frame2_5_0
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__41351\,
            I => data_out_frame2_5_0
        );

    \I__9513\ : Odrv12
    port map (
            O => \N__41348\,
            I => data_out_frame2_5_0
        );

    \I__9512\ : Odrv12
    port map (
            O => \N__41345\,
            I => data_out_frame2_5_0
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__41342\,
            I => data_out_frame2_5_0
        );

    \I__9510\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__41328\,
            I => \c0.n10911\
        );

    \I__9508\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41319\
        );

    \I__9507\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41316\
        );

    \I__9506\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41313\
        );

    \I__9505\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41309\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__41319\,
            I => \N__41306\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__41316\,
            I => \N__41301\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41301\
        );

    \I__9501\ : InMux
    port map (
            O => \N__41312\,
            I => \N__41298\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__41309\,
            I => data_out_frame2_11_6
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__41306\,
            I => data_out_frame2_11_6
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__41301\,
            I => data_out_frame2_11_6
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__41298\,
            I => data_out_frame2_11_6
        );

    \I__9496\ : InMux
    port map (
            O => \N__41289\,
            I => \N__41285\
        );

    \I__9495\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41281\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__41285\,
            I => \N__41277\
        );

    \I__9493\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41274\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41271\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__41280\,
            I => \N__41268\
        );

    \I__9490\ : Span4Mux_h
    port map (
            O => \N__41277\,
            I => \N__41263\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__41274\,
            I => \N__41263\
        );

    \I__9488\ : Span4Mux_h
    port map (
            O => \N__41271\,
            I => \N__41259\
        );

    \I__9487\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41255\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__41263\,
            I => \N__41252\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41249\
        );

    \I__9484\ : Span4Mux_s2_v
    port map (
            O => \N__41259\,
            I => \N__41246\
        );

    \I__9483\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41243\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__41255\,
            I => \N__41240\
        );

    \I__9481\ : Odrv4
    port map (
            O => \N__41252\,
            I => rand_data_6
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__41249\,
            I => rand_data_6
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__41246\,
            I => rand_data_6
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__41243\,
            I => rand_data_6
        );

    \I__9477\ : Odrv12
    port map (
            O => \N__41240\,
            I => rand_data_6
        );

    \I__9476\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41224\
        );

    \I__9475\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41219\
        );

    \I__9474\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41219\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41214\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__41219\,
            I => \N__41211\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41208\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41205\
        );

    \I__9469\ : Span4Mux_s2_v
    port map (
            O => \N__41214\,
            I => \N__41200\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__41211\,
            I => \N__41200\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__41208\,
            I => \N__41197\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__41205\,
            I => data_out_frame2_9_4
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__41200\,
            I => data_out_frame2_9_4
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__41197\,
            I => data_out_frame2_9_4
        );

    \I__9463\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41186\
        );

    \I__9462\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41181\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__41186\,
            I => \N__41178\
        );

    \I__9460\ : InMux
    port map (
            O => \N__41185\,
            I => \N__41175\
        );

    \I__9459\ : InMux
    port map (
            O => \N__41184\,
            I => \N__41172\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__41181\,
            I => \N__41169\
        );

    \I__9457\ : Span4Mux_h
    port map (
            O => \N__41178\,
            I => \N__41166\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__41175\,
            I => \N__41163\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__41172\,
            I => data_out_frame2_7_7
        );

    \I__9454\ : Odrv4
    port map (
            O => \N__41169\,
            I => data_out_frame2_7_7
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__41166\,
            I => data_out_frame2_7_7
        );

    \I__9452\ : Odrv4
    port map (
            O => \N__41163\,
            I => data_out_frame2_7_7
        );

    \I__9451\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41151\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__41151\,
            I => \N__41146\
        );

    \I__9449\ : CascadeMux
    port map (
            O => \N__41150\,
            I => \N__41142\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41139\
        );

    \I__9447\ : Span12Mux_h
    port map (
            O => \N__41146\,
            I => \N__41136\
        );

    \I__9446\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41133\
        );

    \I__9445\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41130\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41139\,
            I => data_out_frame2_9_7
        );

    \I__9443\ : Odrv12
    port map (
            O => \N__41136\,
            I => data_out_frame2_9_7
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__41133\,
            I => data_out_frame2_9_7
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__41130\,
            I => data_out_frame2_9_7
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__41121\,
            I => \N__41118\
        );

    \I__9439\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41112\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__41112\,
            I => \c0.n10617\
        );

    \I__9436\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41106\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41103\
        );

    \I__9434\ : Span4Mux_s2_v
    port map (
            O => \N__41103\,
            I => \N__41100\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__41100\,
            I => \N__41097\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__41097\,
            I => \c0.n14_adj_2362\
        );

    \I__9431\ : CascadeMux
    port map (
            O => \N__41094\,
            I => \N__41091\
        );

    \I__9430\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41086\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41090\,
            I => \N__41083\
        );

    \I__9428\ : InMux
    port map (
            O => \N__41089\,
            I => \N__41079\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__41086\,
            I => \N__41073\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__41083\,
            I => \N__41070\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41082\,
            I => \N__41067\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__41079\,
            I => \N__41064\
        );

    \I__9423\ : InMux
    port map (
            O => \N__41078\,
            I => \N__41059\
        );

    \I__9422\ : InMux
    port map (
            O => \N__41077\,
            I => \N__41059\
        );

    \I__9421\ : InMux
    port map (
            O => \N__41076\,
            I => \N__41056\
        );

    \I__9420\ : Span4Mux_h
    port map (
            O => \N__41073\,
            I => \N__41051\
        );

    \I__9419\ : Span4Mux_v
    port map (
            O => \N__41070\,
            I => \N__41051\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__41067\,
            I => \N__41044\
        );

    \I__9417\ : Span4Mux_h
    port map (
            O => \N__41064\,
            I => \N__41044\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__41059\,
            I => \N__41044\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__41056\,
            I => data_out_frame2_12_2
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__41051\,
            I => data_out_frame2_12_2
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__41044\,
            I => data_out_frame2_12_2
        );

    \I__9412\ : InMux
    port map (
            O => \N__41037\,
            I => \N__41032\
        );

    \I__9411\ : InMux
    port map (
            O => \N__41036\,
            I => \N__41029\
        );

    \I__9410\ : InMux
    port map (
            O => \N__41035\,
            I => \N__41026\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__41032\,
            I => \N__41022\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__41029\,
            I => \N__41019\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__41026\,
            I => \N__41016\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41025\,
            I => \N__41012\
        );

    \I__9405\ : Span4Mux_v
    port map (
            O => \N__41022\,
            I => \N__41009\
        );

    \I__9404\ : Span4Mux_h
    port map (
            O => \N__41019\,
            I => \N__41004\
        );

    \I__9403\ : Span4Mux_s1_v
    port map (
            O => \N__41016\,
            I => \N__41004\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41015\,
            I => \N__41001\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__41012\,
            I => data_out_frame2_10_4
        );

    \I__9400\ : Odrv4
    port map (
            O => \N__41009\,
            I => data_out_frame2_10_4
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__41004\,
            I => data_out_frame2_10_4
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__41001\,
            I => data_out_frame2_10_4
        );

    \I__9397\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40988\
        );

    \I__9396\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40985\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__40988\,
            I => \N__40980\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__40985\,
            I => \N__40977\
        );

    \I__9393\ : InMux
    port map (
            O => \N__40984\,
            I => \N__40973\
        );

    \I__9392\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40970\
        );

    \I__9391\ : Span4Mux_s2_v
    port map (
            O => \N__40980\,
            I => \N__40967\
        );

    \I__9390\ : Span4Mux_s2_v
    port map (
            O => \N__40977\,
            I => \N__40964\
        );

    \I__9389\ : InMux
    port map (
            O => \N__40976\,
            I => \N__40961\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__40973\,
            I => data_out_frame2_16_7
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__40970\,
            I => data_out_frame2_16_7
        );

    \I__9386\ : Odrv4
    port map (
            O => \N__40967\,
            I => data_out_frame2_16_7
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__40964\,
            I => data_out_frame2_16_7
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__40961\,
            I => data_out_frame2_16_7
        );

    \I__9383\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40946\
        );

    \I__9382\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40943\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__40946\,
            I => \N__40937\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__40943\,
            I => \N__40934\
        );

    \I__9379\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40929\
        );

    \I__9378\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40929\
        );

    \I__9377\ : InMux
    port map (
            O => \N__40940\,
            I => \N__40925\
        );

    \I__9376\ : Span4Mux_v
    port map (
            O => \N__40937\,
            I => \N__40918\
        );

    \I__9375\ : Span4Mux_s0_v
    port map (
            O => \N__40934\,
            I => \N__40918\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__40929\,
            I => \N__40918\
        );

    \I__9373\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40915\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__40925\,
            I => \N__40910\
        );

    \I__9371\ : Span4Mux_h
    port map (
            O => \N__40918\,
            I => \N__40910\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__40915\,
            I => data_out_frame2_15_7
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__40910\,
            I => data_out_frame2_15_7
        );

    \I__9368\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__40902\,
            I => \c0.n17889\
        );

    \I__9366\ : InMux
    port map (
            O => \N__40899\,
            I => \N__40896\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__40896\,
            I => \N__40893\
        );

    \I__9364\ : Span4Mux_h
    port map (
            O => \N__40893\,
            I => \N__40888\
        );

    \I__9363\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40885\
        );

    \I__9362\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40882\
        );

    \I__9361\ : Span4Mux_s2_v
    port map (
            O => \N__40888\,
            I => \N__40877\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__40885\,
            I => \N__40877\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__40882\,
            I => \N__40873\
        );

    \I__9358\ : Span4Mux_h
    port map (
            O => \N__40877\,
            I => \N__40870\
        );

    \I__9357\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40866\
        );

    \I__9356\ : Span4Mux_h
    port map (
            O => \N__40873\,
            I => \N__40863\
        );

    \I__9355\ : Span4Mux_v
    port map (
            O => \N__40870\,
            I => \N__40860\
        );

    \I__9354\ : InMux
    port map (
            O => \N__40869\,
            I => \N__40857\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__40866\,
            I => \N__40854\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__40863\,
            I => rand_data_18
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__40860\,
            I => rand_data_18
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__40857\,
            I => rand_data_18
        );

    \I__9349\ : Odrv12
    port map (
            O => \N__40854\,
            I => rand_data_18
        );

    \I__9348\ : CascadeMux
    port map (
            O => \N__40845\,
            I => \N__40841\
        );

    \I__9347\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40836\
        );

    \I__9346\ : InMux
    port map (
            O => \N__40841\,
            I => \N__40831\
        );

    \I__9345\ : InMux
    port map (
            O => \N__40840\,
            I => \N__40831\
        );

    \I__9344\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40828\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40825\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40822\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__40828\,
            I => data_out_frame2_6_2
        );

    \I__9340\ : Odrv12
    port map (
            O => \N__40825\,
            I => data_out_frame2_6_2
        );

    \I__9339\ : Odrv4
    port map (
            O => \N__40822\,
            I => data_out_frame2_6_2
        );

    \I__9338\ : InMux
    port map (
            O => \N__40815\,
            I => \N__40812\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__40812\,
            I => \N__40809\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__40809\,
            I => \N__40806\
        );

    \I__9335\ : Odrv4
    port map (
            O => \N__40806\,
            I => \c0.n18645\
        );

    \I__9334\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40800\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__40800\,
            I => \N__40797\
        );

    \I__9332\ : Span12Mux_h
    port map (
            O => \N__40797\,
            I => \N__40794\
        );

    \I__9331\ : Odrv12
    port map (
            O => \N__40794\,
            I => \c0.n18_adj_2441\
        );

    \I__9330\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40783\
        );

    \I__9328\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40778\
        );

    \I__9327\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40778\
        );

    \I__9326\ : Span4Mux_s2_v
    port map (
            O => \N__40783\,
            I => \N__40772\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__40778\,
            I => \N__40769\
        );

    \I__9324\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40766\
        );

    \I__9323\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40761\
        );

    \I__9322\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40761\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__40772\,
            I => data_out_frame2_8_3
        );

    \I__9320\ : Odrv12
    port map (
            O => \N__40769\,
            I => data_out_frame2_8_3
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__40766\,
            I => data_out_frame2_8_3
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__40761\,
            I => data_out_frame2_8_3
        );

    \I__9317\ : InMux
    port map (
            O => \N__40752\,
            I => \N__40747\
        );

    \I__9316\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40743\
        );

    \I__9315\ : CascadeMux
    port map (
            O => \N__40750\,
            I => \N__40740\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__40747\,
            I => \N__40736\
        );

    \I__9313\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40733\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40730\
        );

    \I__9311\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40725\
        );

    \I__9310\ : InMux
    port map (
            O => \N__40739\,
            I => \N__40725\
        );

    \I__9309\ : Span4Mux_h
    port map (
            O => \N__40736\,
            I => \N__40722\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__40733\,
            I => \N__40719\
        );

    \I__9307\ : Span4Mux_s2_v
    port map (
            O => \N__40730\,
            I => \N__40716\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__40725\,
            I => data_out_frame2_10_1
        );

    \I__9305\ : Odrv4
    port map (
            O => \N__40722\,
            I => data_out_frame2_10_1
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__40719\,
            I => data_out_frame2_10_1
        );

    \I__9303\ : Odrv4
    port map (
            O => \N__40716\,
            I => data_out_frame2_10_1
        );

    \I__9302\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__40704\,
            I => \N__40700\
        );

    \I__9300\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__40700\,
            I => \N__40694\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__40697\,
            I => \c0.n17838\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__40694\,
            I => \c0.n17838\
        );

    \I__9296\ : InMux
    port map (
            O => \N__40689\,
            I => \N__40685\
        );

    \I__9295\ : InMux
    port map (
            O => \N__40688\,
            I => \N__40682\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__40685\,
            I => \N__40679\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__40682\,
            I => \N__40676\
        );

    \I__9292\ : Odrv12
    port map (
            O => \N__40679\,
            I => \c0.n17792\
        );

    \I__9291\ : Odrv4
    port map (
            O => \N__40676\,
            I => \c0.n17792\
        );

    \I__9290\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__40668\,
            I => \c0.n33\
        );

    \I__9288\ : InMux
    port map (
            O => \N__40665\,
            I => \N__40661\
        );

    \I__9287\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40658\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__40661\,
            I => \N__40653\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40650\
        );

    \I__9284\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40647\
        );

    \I__9283\ : InMux
    port map (
            O => \N__40656\,
            I => \N__40644\
        );

    \I__9282\ : Span12Mux_s9_v
    port map (
            O => \N__40653\,
            I => \N__40641\
        );

    \I__9281\ : Span12Mux_s2_v
    port map (
            O => \N__40650\,
            I => \N__40638\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__40647\,
            I => data_out_frame2_6_6
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__40644\,
            I => data_out_frame2_6_6
        );

    \I__9278\ : Odrv12
    port map (
            O => \N__40641\,
            I => data_out_frame2_6_6
        );

    \I__9277\ : Odrv12
    port map (
            O => \N__40638\,
            I => data_out_frame2_6_6
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__40629\,
            I => \N__40626\
        );

    \I__9275\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40623\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__40623\,
            I => \N__40620\
        );

    \I__9273\ : Span4Mux_h
    port map (
            O => \N__40620\,
            I => \N__40617\
        );

    \I__9272\ : Sp12to4
    port map (
            O => \N__40617\,
            I => \N__40614\
        );

    \I__9271\ : Odrv12
    port map (
            O => \N__40614\,
            I => \c0.n17736\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__40611\,
            I => \c0.n17736_cascade_\
        );

    \I__9269\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40605\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__40605\,
            I => \c0.n18813\
        );

    \I__9267\ : CascadeMux
    port map (
            O => \N__40602\,
            I => \N__40599\
        );

    \I__9266\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__40596\,
            I => \N__40593\
        );

    \I__9264\ : Odrv12
    port map (
            O => \N__40593\,
            I => \c0.n18816\
        );

    \I__9263\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40582\
        );

    \I__9262\ : InMux
    port map (
            O => \N__40589\,
            I => \N__40582\
        );

    \I__9261\ : InMux
    port map (
            O => \N__40588\,
            I => \N__40577\
        );

    \I__9260\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40577\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__40582\,
            I => \N__40571\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40577\,
            I => \N__40571\
        );

    \I__9257\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40568\
        );

    \I__9256\ : Span4Mux_s1_v
    port map (
            O => \N__40571\,
            I => \N__40565\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__40568\,
            I => data_out_frame2_9_6
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__40565\,
            I => data_out_frame2_9_6
        );

    \I__9253\ : InMux
    port map (
            O => \N__40560\,
            I => \N__40557\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__40557\,
            I => \N__40554\
        );

    \I__9251\ : Odrv12
    port map (
            O => \N__40554\,
            I => \c0.n10725\
        );

    \I__9250\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40546\
        );

    \I__9249\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40543\
        );

    \I__9248\ : InMux
    port map (
            O => \N__40549\,
            I => \N__40540\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__40546\,
            I => \N__40537\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__40543\,
            I => \N__40530\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40530\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__40537\,
            I => \N__40527\
        );

    \I__9243\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40524\
        );

    \I__9242\ : InMux
    port map (
            O => \N__40535\,
            I => \N__40521\
        );

    \I__9241\ : Span4Mux_h
    port map (
            O => \N__40530\,
            I => \N__40516\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__40527\,
            I => \N__40516\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__40524\,
            I => data_out_frame2_7_0
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__40521\,
            I => data_out_frame2_7_0
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__40516\,
            I => data_out_frame2_7_0
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \N__40506\
        );

    \I__9235\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40503\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__40503\,
            I => \N__40500\
        );

    \I__9233\ : Span4Mux_h
    port map (
            O => \N__40500\,
            I => \N__40497\
        );

    \I__9232\ : IoSpan4Mux
    port map (
            O => \N__40497\,
            I => \N__40494\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__40494\,
            I => \c0.n10700\
        );

    \I__9230\ : InMux
    port map (
            O => \N__40491\,
            I => \N__40488\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__40488\,
            I => \N__40485\
        );

    \I__9228\ : Span12Mux_h
    port map (
            O => \N__40485\,
            I => \N__40482\
        );

    \I__9227\ : Odrv12
    port map (
            O => \N__40482\,
            I => \c0.n16_adj_2412\
        );

    \I__9226\ : CascadeMux
    port map (
            O => \N__40479\,
            I => \c0.n17_adj_2413_cascade_\
        );

    \I__9225\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40472\
        );

    \I__9224\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40469\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__40472\,
            I => \N__40463\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__40469\,
            I => \N__40463\
        );

    \I__9221\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40459\
        );

    \I__9220\ : Span4Mux_v
    port map (
            O => \N__40463\,
            I => \N__40456\
        );

    \I__9219\ : CascadeMux
    port map (
            O => \N__40462\,
            I => \N__40453\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__40459\,
            I => \N__40448\
        );

    \I__9217\ : Sp12to4
    port map (
            O => \N__40456\,
            I => \N__40448\
        );

    \I__9216\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40445\
        );

    \I__9215\ : Span12Mux_h
    port map (
            O => \N__40448\,
            I => \N__40442\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__40445\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__9213\ : Odrv12
    port map (
            O => \N__40442\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__9212\ : InMux
    port map (
            O => \N__40437\,
            I => \N__40433\
        );

    \I__9211\ : CascadeMux
    port map (
            O => \N__40436\,
            I => \N__40430\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__40433\,
            I => \N__40427\
        );

    \I__9209\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40424\
        );

    \I__9208\ : Span4Mux_h
    port map (
            O => \N__40427\,
            I => \N__40421\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__40424\,
            I => \N__40418\
        );

    \I__9206\ : Span4Mux_v
    port map (
            O => \N__40421\,
            I => \N__40415\
        );

    \I__9205\ : Span12Mux_s8_v
    port map (
            O => \N__40418\,
            I => \N__40412\
        );

    \I__9204\ : Odrv4
    port map (
            O => \N__40415\,
            I => \c0.n10782\
        );

    \I__9203\ : Odrv12
    port map (
            O => \N__40412\,
            I => \c0.n10782\
        );

    \I__9202\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40403\
        );

    \I__9201\ : CascadeMux
    port map (
            O => \N__40406\,
            I => \N__40400\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40397\
        );

    \I__9199\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40393\
        );

    \I__9198\ : IoSpan4Mux
    port map (
            O => \N__40397\,
            I => \N__40390\
        );

    \I__9197\ : InMux
    port map (
            O => \N__40396\,
            I => \N__40386\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__40393\,
            I => \N__40381\
        );

    \I__9195\ : IoSpan4Mux
    port map (
            O => \N__40390\,
            I => \N__40381\
        );

    \I__9194\ : InMux
    port map (
            O => \N__40389\,
            I => \N__40378\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__40386\,
            I => data_out_frame2_14_1
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__40381\,
            I => data_out_frame2_14_1
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__40378\,
            I => data_out_frame2_14_1
        );

    \I__9190\ : InMux
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__40368\,
            I => \c0.n17862\
        );

    \I__9188\ : CascadeMux
    port map (
            O => \N__40365\,
            I => \c0.n17862_cascade_\
        );

    \I__9187\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40359\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__40359\,
            I => \N__40356\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__40356\,
            I => \N__40352\
        );

    \I__9184\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40349\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__40352\,
            I => \c0.n17841\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__40349\,
            I => \c0.n17841\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__40344\,
            I => \c0.n12_adj_2410_cascade_\
        );

    \I__9180\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__40338\,
            I => \N__40335\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__40335\,
            I => \N__40331\
        );

    \I__9177\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40328\
        );

    \I__9176\ : Odrv4
    port map (
            O => \N__40331\,
            I => \c0.n17718\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__40328\,
            I => \c0.n17718\
        );

    \I__9174\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40319\
        );

    \I__9173\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40316\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__40319\,
            I => \c0.n17829\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__40316\,
            I => \c0.n17829\
        );

    \I__9170\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40306\
        );

    \I__9169\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40303\
        );

    \I__9168\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40300\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__40306\,
            I => \N__40297\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__40303\,
            I => \N__40294\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__40300\,
            I => \N__40291\
        );

    \I__9164\ : Span4Mux_v
    port map (
            O => \N__40297\,
            I => \N__40286\
        );

    \I__9163\ : Span4Mux_h
    port map (
            O => \N__40294\,
            I => \N__40286\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__40291\,
            I => \c0.data_out_10_4\
        );

    \I__9161\ : Odrv4
    port map (
            O => \N__40286\,
            I => \c0.data_out_10_4\
        );

    \I__9160\ : InMux
    port map (
            O => \N__40281\,
            I => \N__40278\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__40278\,
            I => \N__40274\
        );

    \I__9158\ : InMux
    port map (
            O => \N__40277\,
            I => \N__40271\
        );

    \I__9157\ : Span4Mux_v
    port map (
            O => \N__40274\,
            I => \N__40267\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40264\
        );

    \I__9155\ : InMux
    port map (
            O => \N__40270\,
            I => \N__40261\
        );

    \I__9154\ : Span4Mux_h
    port map (
            O => \N__40267\,
            I => \N__40258\
        );

    \I__9153\ : Span4Mux_h
    port map (
            O => \N__40264\,
            I => \N__40255\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__40261\,
            I => \N__40252\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__40258\,
            I => n2837
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__40255\,
            I => n2837
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__40252\,
            I => n2837
        );

    \I__9148\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40239\
        );

    \I__9147\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40239\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__40239\,
            I => data_out_3_0
        );

    \I__9145\ : InMux
    port map (
            O => \N__40236\,
            I => \N__40233\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__40233\,
            I => \N__40230\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__40230\,
            I => \c0.n2_adj_2221\
        );

    \I__9142\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40221\
        );

    \I__9141\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40221\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__40221\,
            I => data_out_2_0
        );

    \I__9139\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__40215\,
            I => \N__40212\
        );

    \I__9137\ : Span4Mux_s0_v
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__9136\ : Span4Mux_h
    port map (
            O => \N__40209\,
            I => \N__40206\
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__40206\,
            I => \c0.n5_adj_2433\
        );

    \I__9134\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__40200\,
            I => \N__40194\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40189\
        );

    \I__9131\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40189\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40186\
        );

    \I__9129\ : Span4Mux_s2_v
    port map (
            O => \N__40194\,
            I => \N__40183\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__40189\,
            I => \N__40180\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__40186\,
            I => data_out_frame2_14_7
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__40183\,
            I => data_out_frame2_14_7
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__40180\,
            I => data_out_frame2_14_7
        );

    \I__9124\ : InMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__40170\,
            I => \c0.n17899\
        );

    \I__9122\ : CascadeMux
    port map (
            O => \N__40167\,
            I => \c0.n17899_cascade_\
        );

    \I__9121\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40161\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__40161\,
            I => \N__40158\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__9118\ : Span4Mux_s0_v
    port map (
            O => \N__40155\,
            I => \N__40152\
        );

    \I__9117\ : Odrv4
    port map (
            O => \N__40152\,
            I => \c0.n34\
        );

    \I__9116\ : InMux
    port map (
            O => \N__40149\,
            I => \N__40143\
        );

    \I__9115\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40140\
        );

    \I__9114\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40137\
        );

    \I__9113\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40134\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__40143\,
            I => \N__40131\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__40140\,
            I => \N__40126\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__40137\,
            I => \N__40126\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__40134\,
            I => \N__40122\
        );

    \I__9108\ : Span4Mux_h
    port map (
            O => \N__40131\,
            I => \N__40119\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__40126\,
            I => \N__40116\
        );

    \I__9106\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40113\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__40122\,
            I => \N__40110\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__40119\,
            I => rand_data_30
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__40116\,
            I => rand_data_30
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__40113\,
            I => rand_data_30
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__40110\,
            I => rand_data_30
        );

    \I__9100\ : InMux
    port map (
            O => \N__40101\,
            I => n16607
        );

    \I__9099\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40093\
        );

    \I__9098\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40089\
        );

    \I__9097\ : InMux
    port map (
            O => \N__40096\,
            I => \N__40086\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__40093\,
            I => \N__40083\
        );

    \I__9095\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40080\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__40089\,
            I => \N__40077\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__40086\,
            I => \N__40073\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__40083\,
            I => \N__40070\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__40080\,
            I => \N__40067\
        );

    \I__9090\ : Span4Mux_s3_v
    port map (
            O => \N__40077\,
            I => \N__40064\
        );

    \I__9089\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40061\
        );

    \I__9088\ : Span4Mux_v
    port map (
            O => \N__40073\,
            I => \N__40058\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__40070\,
            I => \N__40051\
        );

    \I__9086\ : Span4Mux_v
    port map (
            O => \N__40067\,
            I => \N__40051\
        );

    \I__9085\ : Span4Mux_v
    port map (
            O => \N__40064\,
            I => \N__40051\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__40061\,
            I => rand_data_31
        );

    \I__9083\ : Odrv4
    port map (
            O => \N__40058\,
            I => rand_data_31
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__40051\,
            I => rand_data_31
        );

    \I__9081\ : InMux
    port map (
            O => \N__40044\,
            I => n16608
        );

    \I__9080\ : InMux
    port map (
            O => \N__40041\,
            I => \N__40037\
        );

    \I__9079\ : CascadeMux
    port map (
            O => \N__40040\,
            I => \N__40034\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__40037\,
            I => \N__40031\
        );

    \I__9077\ : InMux
    port map (
            O => \N__40034\,
            I => \N__40028\
        );

    \I__9076\ : Odrv4
    port map (
            O => \N__40031\,
            I => rand_setpoint_13
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__40028\,
            I => rand_setpoint_13
        );

    \I__9074\ : CascadeMux
    port map (
            O => \N__40023\,
            I => \N__40020\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40017\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__40017\,
            I => \N__40014\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__40014\,
            I => \c0.n18234\
        );

    \I__9070\ : InMux
    port map (
            O => \N__40011\,
            I => \N__40007\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__40010\,
            I => \N__40004\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__40007\,
            I => \N__40001\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39998\
        );

    \I__9066\ : Odrv12
    port map (
            O => \N__40001\,
            I => rand_setpoint_1
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__39998\,
            I => rand_setpoint_1
        );

    \I__9064\ : CascadeMux
    port map (
            O => \N__39993\,
            I => \N__39990\
        );

    \I__9063\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39987\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39981\
        );

    \I__9061\ : InMux
    port map (
            O => \N__39986\,
            I => \N__39978\
        );

    \I__9060\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39973\
        );

    \I__9059\ : InMux
    port map (
            O => \N__39984\,
            I => \N__39973\
        );

    \I__9058\ : Span4Mux_v
    port map (
            O => \N__39981\,
            I => \N__39969\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__39978\,
            I => \N__39966\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__39973\,
            I => \N__39963\
        );

    \I__9055\ : InMux
    port map (
            O => \N__39972\,
            I => \N__39960\
        );

    \I__9054\ : Span4Mux_v
    port map (
            O => \N__39969\,
            I => \N__39957\
        );

    \I__9053\ : Span4Mux_h
    port map (
            O => \N__39966\,
            I => \N__39954\
        );

    \I__9052\ : Span4Mux_h
    port map (
            O => \N__39963\,
            I => \N__39951\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__39960\,
            I => \c0.data_out_8_1\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__39957\,
            I => \c0.data_out_8_1\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__39954\,
            I => \c0.data_out_8_1\
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__39951\,
            I => \c0.data_out_8_1\
        );

    \I__9047\ : InMux
    port map (
            O => \N__39942\,
            I => \N__39938\
        );

    \I__9046\ : InMux
    port map (
            O => \N__39941\,
            I => \N__39935\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__39938\,
            I => \N__39932\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__39935\,
            I => \N__39927\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__39932\,
            I => \N__39924\
        );

    \I__9042\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39919\
        );

    \I__9041\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39919\
        );

    \I__9040\ : Span4Mux_h
    port map (
            O => \N__39927\,
            I => \N__39916\
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__39924\,
            I => \c0.data_out_7_5\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__39919\,
            I => \c0.data_out_7_5\
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__39916\,
            I => \c0.data_out_7_5\
        );

    \I__9036\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39904\
        );

    \I__9035\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39901\
        );

    \I__9034\ : InMux
    port map (
            O => \N__39907\,
            I => \N__39897\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__39904\,
            I => \N__39894\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__39901\,
            I => \N__39890\
        );

    \I__9031\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39887\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__39897\,
            I => \N__39884\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__39894\,
            I => \N__39881\
        );

    \I__9028\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39878\
        );

    \I__9027\ : Span4Mux_h
    port map (
            O => \N__39890\,
            I => \N__39875\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__39887\,
            I => \c0.data_out_7_7\
        );

    \I__9025\ : Odrv12
    port map (
            O => \N__39884\,
            I => \c0.data_out_7_7\
        );

    \I__9024\ : Odrv4
    port map (
            O => \N__39881\,
            I => \c0.data_out_7_7\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__39878\,
            I => \c0.data_out_7_7\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__39875\,
            I => \c0.data_out_7_7\
        );

    \I__9021\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39861\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__39858\,
            I => \c0.n10533\
        );

    \I__9018\ : InMux
    port map (
            O => \N__39855\,
            I => \N__39851\
        );

    \I__9017\ : CascadeMux
    port map (
            O => \N__39854\,
            I => \N__39848\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__39851\,
            I => \N__39845\
        );

    \I__9015\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__39845\,
            I => rand_setpoint_26
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__39842\,
            I => rand_setpoint_26
        );

    \I__9012\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39831\
        );

    \I__9011\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39826\
        );

    \I__9010\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39826\
        );

    \I__9009\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39823\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__39831\,
            I => \N__39816\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__39826\,
            I => \N__39816\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__39823\,
            I => \N__39813\
        );

    \I__9005\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39810\
        );

    \I__9004\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39807\
        );

    \I__9003\ : Span4Mux_h
    port map (
            O => \N__39816\,
            I => \N__39804\
        );

    \I__9002\ : Span4Mux_h
    port map (
            O => \N__39813\,
            I => \N__39801\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__39810\,
            I => \c0.data_out_5_2\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__39807\,
            I => \c0.data_out_5_2\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__39804\,
            I => \c0.data_out_5_2\
        );

    \I__8998\ : Odrv4
    port map (
            O => \N__39801\,
            I => \c0.data_out_5_2\
        );

    \I__8997\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39788\
        );

    \I__8996\ : CascadeMux
    port map (
            O => \N__39791\,
            I => \N__39785\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__39788\,
            I => \N__39782\
        );

    \I__8994\ : InMux
    port map (
            O => \N__39785\,
            I => \N__39779\
        );

    \I__8993\ : Odrv4
    port map (
            O => \N__39782\,
            I => rand_setpoint_30
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__39779\,
            I => rand_setpoint_30
        );

    \I__8991\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39770\
        );

    \I__8990\ : CascadeMux
    port map (
            O => \N__39773\,
            I => \N__39767\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__39770\,
            I => \N__39764\
        );

    \I__8988\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39761\
        );

    \I__8987\ : Odrv4
    port map (
            O => \N__39764\,
            I => rand_setpoint_27
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__39761\,
            I => rand_setpoint_27
        );

    \I__8985\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39752\
        );

    \I__8984\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39747\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__39752\,
            I => \N__39744\
        );

    \I__8982\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39736\
        );

    \I__8981\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39736\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39733\
        );

    \I__8979\ : Span4Mux_v
    port map (
            O => \N__39744\,
            I => \N__39730\
        );

    \I__8978\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39727\
        );

    \I__8977\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39722\
        );

    \I__8976\ : InMux
    port map (
            O => \N__39741\,
            I => \N__39722\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__39736\,
            I => \N__39719\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__39733\,
            I => \N__39716\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__39730\,
            I => \c0.data_out_5_3\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__39727\,
            I => \c0.data_out_5_3\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__39722\,
            I => \c0.data_out_5_3\
        );

    \I__8970\ : Odrv4
    port map (
            O => \N__39719\,
            I => \c0.data_out_5_3\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__39716\,
            I => \c0.data_out_5_3\
        );

    \I__8968\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39701\
        );

    \I__8967\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39696\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__39701\,
            I => \N__39693\
        );

    \I__8965\ : InMux
    port map (
            O => \N__39700\,
            I => \N__39690\
        );

    \I__8964\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39687\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__39696\,
            I => \N__39684\
        );

    \I__8962\ : Span4Mux_v
    port map (
            O => \N__39693\,
            I => \N__39681\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__39690\,
            I => \N__39677\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__39687\,
            I => \N__39674\
        );

    \I__8959\ : Span4Mux_h
    port map (
            O => \N__39684\,
            I => \N__39669\
        );

    \I__8958\ : Span4Mux_h
    port map (
            O => \N__39681\,
            I => \N__39669\
        );

    \I__8957\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39666\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__39677\,
            I => \N__39661\
        );

    \I__8955\ : Span4Mux_v
    port map (
            O => \N__39674\,
            I => \N__39661\
        );

    \I__8954\ : Odrv4
    port map (
            O => \N__39669\,
            I => rand_data_22
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__39666\,
            I => rand_data_22
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__39661\,
            I => rand_data_22
        );

    \I__8951\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39650\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__39653\,
            I => \N__39647\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__39650\,
            I => \N__39644\
        );

    \I__8948\ : InMux
    port map (
            O => \N__39647\,
            I => \N__39641\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__39644\,
            I => rand_setpoint_22
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__39641\,
            I => rand_setpoint_22
        );

    \I__8945\ : InMux
    port map (
            O => \N__39636\,
            I => n16599
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__39633\,
            I => \N__39629\
        );

    \I__8943\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39626\
        );

    \I__8942\ : InMux
    port map (
            O => \N__39629\,
            I => \N__39621\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__39626\,
            I => \N__39618\
        );

    \I__8940\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39615\
        );

    \I__8939\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39612\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__39621\,
            I => \N__39609\
        );

    \I__8937\ : Span4Mux_h
    port map (
            O => \N__39618\,
            I => \N__39606\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__39615\,
            I => \N__39603\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__39612\,
            I => \N__39599\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__39609\,
            I => \N__39596\
        );

    \I__8933\ : Span4Mux_v
    port map (
            O => \N__39606\,
            I => \N__39591\
        );

    \I__8932\ : Span4Mux_v
    port map (
            O => \N__39603\,
            I => \N__39591\
        );

    \I__8931\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39588\
        );

    \I__8930\ : Span4Mux_v
    port map (
            O => \N__39599\,
            I => \N__39585\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__39596\,
            I => rand_data_23
        );

    \I__8928\ : Odrv4
    port map (
            O => \N__39591\,
            I => rand_data_23
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__39588\,
            I => rand_data_23
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__39585\,
            I => rand_data_23
        );

    \I__8925\ : CascadeMux
    port map (
            O => \N__39576\,
            I => \N__39572\
        );

    \I__8924\ : CascadeMux
    port map (
            O => \N__39575\,
            I => \N__39569\
        );

    \I__8923\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39566\
        );

    \I__8922\ : InMux
    port map (
            O => \N__39569\,
            I => \N__39563\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__39566\,
            I => rand_setpoint_23
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__39563\,
            I => rand_setpoint_23
        );

    \I__8919\ : InMux
    port map (
            O => \N__39558\,
            I => n16600
        );

    \I__8918\ : InMux
    port map (
            O => \N__39555\,
            I => \N__39549\
        );

    \I__8917\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39546\
        );

    \I__8916\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39543\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__39552\,
            I => \N__39540\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__39549\,
            I => \N__39534\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39534\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39531\
        );

    \I__8911\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39528\
        );

    \I__8910\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39525\
        );

    \I__8909\ : Span4Mux_h
    port map (
            O => \N__39534\,
            I => \N__39520\
        );

    \I__8908\ : Span4Mux_v
    port map (
            O => \N__39531\,
            I => \N__39520\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__39528\,
            I => rand_data_24
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39525\,
            I => rand_data_24
        );

    \I__8905\ : Odrv4
    port map (
            O => \N__39520\,
            I => rand_data_24
        );

    \I__8904\ : InMux
    port map (
            O => \N__39513\,
            I => \bfn_14_12_0_\
        );

    \I__8903\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39507\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__39507\,
            I => \N__39504\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__39504\,
            I => \N__39499\
        );

    \I__8900\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39496\
        );

    \I__8899\ : InMux
    port map (
            O => \N__39502\,
            I => \N__39493\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__39499\,
            I => \N__39489\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__39496\,
            I => \N__39484\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__39493\,
            I => \N__39484\
        );

    \I__8895\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39481\
        );

    \I__8894\ : Sp12to4
    port map (
            O => \N__39489\,
            I => \N__39478\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__39484\,
            I => \N__39474\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__39481\,
            I => \N__39471\
        );

    \I__8891\ : Span12Mux_v
    port map (
            O => \N__39478\,
            I => \N__39468\
        );

    \I__8890\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39465\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__39474\,
            I => \N__39460\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__39471\,
            I => \N__39460\
        );

    \I__8887\ : Odrv12
    port map (
            O => \N__39468\,
            I => rand_data_25
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__39465\,
            I => rand_data_25
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__39460\,
            I => rand_data_25
        );

    \I__8884\ : CascadeMux
    port map (
            O => \N__39453\,
            I => \N__39450\
        );

    \I__8883\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39447\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__39447\,
            I => \N__39443\
        );

    \I__8881\ : CascadeMux
    port map (
            O => \N__39446\,
            I => \N__39440\
        );

    \I__8880\ : Span4Mux_v
    port map (
            O => \N__39443\,
            I => \N__39437\
        );

    \I__8879\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39434\
        );

    \I__8878\ : Odrv4
    port map (
            O => \N__39437\,
            I => rand_setpoint_25
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__39434\,
            I => rand_setpoint_25
        );

    \I__8876\ : InMux
    port map (
            O => \N__39429\,
            I => n16602
        );

    \I__8875\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39419\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39419\
        );

    \I__8873\ : InMux
    port map (
            O => \N__39424\,
            I => \N__39416\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39412\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__39416\,
            I => \N__39408\
        );

    \I__8870\ : InMux
    port map (
            O => \N__39415\,
            I => \N__39405\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__39412\,
            I => \N__39402\
        );

    \I__8868\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39399\
        );

    \I__8867\ : Span12Mux_s5_v
    port map (
            O => \N__39408\,
            I => \N__39394\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__39405\,
            I => \N__39394\
        );

    \I__8865\ : Odrv4
    port map (
            O => \N__39402\,
            I => rand_data_26
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__39399\,
            I => rand_data_26
        );

    \I__8863\ : Odrv12
    port map (
            O => \N__39394\,
            I => rand_data_26
        );

    \I__8862\ : InMux
    port map (
            O => \N__39387\,
            I => n16603
        );

    \I__8861\ : InMux
    port map (
            O => \N__39384\,
            I => n16604
        );

    \I__8860\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39378\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39375\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__39375\,
            I => \N__39371\
        );

    \I__8857\ : CascadeMux
    port map (
            O => \N__39374\,
            I => \N__39368\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__39371\,
            I => \N__39365\
        );

    \I__8855\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39362\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__39365\,
            I => rand_setpoint_28
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__39362\,
            I => rand_setpoint_28
        );

    \I__8852\ : InMux
    port map (
            O => \N__39357\,
            I => n16605
        );

    \I__8851\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39351\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39347\
        );

    \I__8849\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39344\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__39347\,
            I => \N__39337\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__39344\,
            I => \N__39337\
        );

    \I__8846\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39334\
        );

    \I__8845\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39331\
        );

    \I__8844\ : Span4Mux_h
    port map (
            O => \N__39337\,
            I => \N__39326\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__39334\,
            I => \N__39326\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__39331\,
            I => \N__39322\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__39326\,
            I => \N__39319\
        );

    \I__8840\ : InMux
    port map (
            O => \N__39325\,
            I => \N__39316\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__39322\,
            I => \N__39313\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__39319\,
            I => rand_data_29
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__39316\,
            I => rand_data_29
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__39313\,
            I => rand_data_29
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__39306\,
            I => \N__39302\
        );

    \I__8834\ : InMux
    port map (
            O => \N__39305\,
            I => \N__39299\
        );

    \I__8833\ : InMux
    port map (
            O => \N__39302\,
            I => \N__39296\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__39299\,
            I => rand_setpoint_29
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__39296\,
            I => rand_setpoint_29
        );

    \I__8830\ : InMux
    port map (
            O => \N__39291\,
            I => n16606
        );

    \I__8829\ : CascadeMux
    port map (
            O => \N__39288\,
            I => \N__39284\
        );

    \I__8828\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39279\
        );

    \I__8827\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39275\
        );

    \I__8826\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39272\
        );

    \I__8825\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39269\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__39279\,
            I => \N__39266\
        );

    \I__8823\ : InMux
    port map (
            O => \N__39278\,
            I => \N__39262\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__39275\,
            I => \N__39257\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__39272\,
            I => \N__39257\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39252\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__39266\,
            I => \N__39252\
        );

    \I__8818\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39249\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__39262\,
            I => \N__39244\
        );

    \I__8816\ : Sp12to4
    port map (
            O => \N__39257\,
            I => \N__39244\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__39252\,
            I => rand_data_14
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__39249\,
            I => rand_data_14
        );

    \I__8813\ : Odrv12
    port map (
            O => \N__39244\,
            I => rand_data_14
        );

    \I__8812\ : InMux
    port map (
            O => \N__39237\,
            I => n16591
        );

    \I__8811\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39225\
        );

    \I__8810\ : InMux
    port map (
            O => \N__39233\,
            I => \N__39225\
        );

    \I__8809\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39222\
        );

    \I__8808\ : InMux
    port map (
            O => \N__39231\,
            I => \N__39219\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__39230\,
            I => \N__39216\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39213\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39208\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__39219\,
            I => \N__39208\
        );

    \I__8803\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39204\
        );

    \I__8802\ : Span4Mux_h
    port map (
            O => \N__39213\,
            I => \N__39201\
        );

    \I__8801\ : Span4Mux_h
    port map (
            O => \N__39208\,
            I => \N__39198\
        );

    \I__8800\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39195\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__39204\,
            I => \N__39192\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__39201\,
            I => rand_data_15
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__39198\,
            I => rand_data_15
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__39195\,
            I => rand_data_15
        );

    \I__8795\ : Odrv12
    port map (
            O => \N__39192\,
            I => rand_data_15
        );

    \I__8794\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__39180\,
            I => \N__39177\
        );

    \I__8792\ : Span4Mux_h
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8791\ : Span4Mux_v
    port map (
            O => \N__39174\,
            I => \N__39170\
        );

    \I__8790\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39167\
        );

    \I__8789\ : Odrv4
    port map (
            O => \N__39170\,
            I => rand_setpoint_15
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__39167\,
            I => rand_setpoint_15
        );

    \I__8787\ : InMux
    port map (
            O => \N__39162\,
            I => n16592
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__8785\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39152\
        );

    \I__8784\ : InMux
    port map (
            O => \N__39155\,
            I => \N__39149\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__39152\,
            I => \N__39143\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39143\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39140\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__39143\,
            I => \N__39137\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39140\,
            I => \N__39132\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__39137\,
            I => \N__39129\
        );

    \I__8777\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39126\
        );

    \I__8776\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39123\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__39132\,
            I => \N__39120\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__39129\,
            I => rand_data_16
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__39126\,
            I => rand_data_16
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__39123\,
            I => rand_data_16
        );

    \I__8771\ : Odrv4
    port map (
            O => \N__39120\,
            I => rand_data_16
        );

    \I__8770\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__39108\,
            I => \N__39104\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__39107\,
            I => \N__39101\
        );

    \I__8767\ : Span4Mux_v
    port map (
            O => \N__39104\,
            I => \N__39098\
        );

    \I__8766\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39095\
        );

    \I__8765\ : Odrv4
    port map (
            O => \N__39098\,
            I => rand_setpoint_16
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__39095\,
            I => rand_setpoint_16
        );

    \I__8763\ : InMux
    port map (
            O => \N__39090\,
            I => \bfn_14_11_0_\
        );

    \I__8762\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39082\
        );

    \I__8761\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39079\
        );

    \I__8760\ : InMux
    port map (
            O => \N__39085\,
            I => \N__39076\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__39082\,
            I => \N__39071\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39071\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8756\ : Span4Mux_v
    port map (
            O => \N__39071\,
            I => \N__39064\
        );

    \I__8755\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39061\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__39067\,
            I => \N__39056\
        );

    \I__8753\ : Span4Mux_s2_v
    port map (
            O => \N__39064\,
            I => \N__39056\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39052\
        );

    \I__8751\ : Span4Mux_h
    port map (
            O => \N__39056\,
            I => \N__39049\
        );

    \I__8750\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39046\
        );

    \I__8749\ : Span4Mux_v
    port map (
            O => \N__39052\,
            I => \N__39043\
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__39049\,
            I => rand_data_17
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__39046\,
            I => rand_data_17
        );

    \I__8746\ : Odrv4
    port map (
            O => \N__39043\,
            I => rand_data_17
        );

    \I__8745\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8743\ : Span4Mux_v
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__39027\,
            I => \N__39023\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__8739\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__39017\,
            I => rand_setpoint_17
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__39014\,
            I => rand_setpoint_17
        );

    \I__8736\ : InMux
    port map (
            O => \N__39009\,
            I => n16594
        );

    \I__8735\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39003\,
            I => \N__38999\
        );

    \I__8733\ : CascadeMux
    port map (
            O => \N__39002\,
            I => \N__38996\
        );

    \I__8732\ : Span4Mux_h
    port map (
            O => \N__38999\,
            I => \N__38993\
        );

    \I__8731\ : InMux
    port map (
            O => \N__38996\,
            I => \N__38990\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__38993\,
            I => rand_setpoint_18
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__38990\,
            I => rand_setpoint_18
        );

    \I__8728\ : InMux
    port map (
            O => \N__38985\,
            I => n16595
        );

    \I__8727\ : InMux
    port map (
            O => \N__38982\,
            I => \N__38976\
        );

    \I__8726\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38973\
        );

    \I__8725\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38970\
        );

    \I__8724\ : InMux
    port map (
            O => \N__38979\,
            I => \N__38967\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__38976\,
            I => \N__38964\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__38973\,
            I => \N__38961\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38957\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__38967\,
            I => \N__38954\
        );

    \I__8719\ : Span4Mux_v
    port map (
            O => \N__38964\,
            I => \N__38951\
        );

    \I__8718\ : Span4Mux_v
    port map (
            O => \N__38961\,
            I => \N__38948\
        );

    \I__8717\ : InMux
    port map (
            O => \N__38960\,
            I => \N__38945\
        );

    \I__8716\ : Span4Mux_v
    port map (
            O => \N__38957\,
            I => \N__38940\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__38954\,
            I => \N__38940\
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__38951\,
            I => rand_data_19
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__38948\,
            I => rand_data_19
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__38945\,
            I => rand_data_19
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__38940\,
            I => rand_data_19
        );

    \I__8710\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__38928\,
            I => \N__38924\
        );

    \I__8708\ : CascadeMux
    port map (
            O => \N__38927\,
            I => \N__38921\
        );

    \I__8707\ : Span4Mux_h
    port map (
            O => \N__38924\,
            I => \N__38918\
        );

    \I__8706\ : InMux
    port map (
            O => \N__38921\,
            I => \N__38915\
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__38918\,
            I => rand_setpoint_19
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__38915\,
            I => rand_setpoint_19
        );

    \I__8703\ : InMux
    port map (
            O => \N__38910\,
            I => n16596
        );

    \I__8702\ : InMux
    port map (
            O => \N__38907\,
            I => \N__38901\
        );

    \I__8701\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38898\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__38905\,
            I => \N__38895\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__38904\,
            I => \N__38892\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__38901\,
            I => \N__38888\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__38898\,
            I => \N__38885\
        );

    \I__8696\ : InMux
    port map (
            O => \N__38895\,
            I => \N__38880\
        );

    \I__8695\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38880\
        );

    \I__8694\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38877\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__38888\,
            I => \N__38872\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__38885\,
            I => \N__38872\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__38880\,
            I => rand_data_20
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__38877\,
            I => rand_data_20
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__38872\,
            I => rand_data_20
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__38865\,
            I => \N__38861\
        );

    \I__8687\ : InMux
    port map (
            O => \N__38864\,
            I => \N__38858\
        );

    \I__8686\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38855\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__38858\,
            I => rand_setpoint_20
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__38855\,
            I => rand_setpoint_20
        );

    \I__8683\ : InMux
    port map (
            O => \N__38850\,
            I => n16597
        );

    \I__8682\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38843\
        );

    \I__8681\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38840\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__38843\,
            I => \N__38835\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__38840\,
            I => \N__38832\
        );

    \I__8678\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38829\
        );

    \I__8677\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38826\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__38835\,
            I => \N__38823\
        );

    \I__8675\ : Span4Mux_v
    port map (
            O => \N__38832\,
            I => \N__38820\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__38829\,
            I => \N__38817\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__38826\,
            I => \N__38813\
        );

    \I__8672\ : Span4Mux_h
    port map (
            O => \N__38823\,
            I => \N__38810\
        );

    \I__8671\ : Span4Mux_h
    port map (
            O => \N__38820\,
            I => \N__38805\
        );

    \I__8670\ : Span4Mux_v
    port map (
            O => \N__38817\,
            I => \N__38805\
        );

    \I__8669\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38802\
        );

    \I__8668\ : Span4Mux_v
    port map (
            O => \N__38813\,
            I => \N__38799\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__38810\,
            I => rand_data_21
        );

    \I__8666\ : Odrv4
    port map (
            O => \N__38805\,
            I => rand_data_21
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__38802\,
            I => rand_data_21
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__38799\,
            I => rand_data_21
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__38790\,
            I => \N__38786\
        );

    \I__8662\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38783\
        );

    \I__8661\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38780\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__38783\,
            I => rand_setpoint_21
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__38780\,
            I => rand_setpoint_21
        );

    \I__8658\ : InMux
    port map (
            O => \N__38775\,
            I => n16598
        );

    \I__8657\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38769\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__38769\,
            I => \N__38766\
        );

    \I__8655\ : Span4Mux_v
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__8654\ : Span4Mux_v
    port map (
            O => \N__38763\,
            I => \N__38759\
        );

    \I__8653\ : InMux
    port map (
            O => \N__38762\,
            I => \N__38756\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__38759\,
            I => rand_setpoint_6
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__38756\,
            I => rand_setpoint_6
        );

    \I__8650\ : InMux
    port map (
            O => \N__38751\,
            I => n16583
        );

    \I__8649\ : InMux
    port map (
            O => \N__38748\,
            I => \N__38745\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__8646\ : Span4Mux_h
    port map (
            O => \N__38739\,
            I => \N__38735\
        );

    \I__8645\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38732\
        );

    \I__8644\ : Odrv4
    port map (
            O => \N__38735\,
            I => rand_setpoint_7
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__38732\,
            I => rand_setpoint_7
        );

    \I__8642\ : InMux
    port map (
            O => \N__38727\,
            I => n16584
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__38724\,
            I => \N__38721\
        );

    \I__8640\ : InMux
    port map (
            O => \N__38721\,
            I => \N__38716\
        );

    \I__8639\ : InMux
    port map (
            O => \N__38720\,
            I => \N__38712\
        );

    \I__8638\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38709\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38706\
        );

    \I__8636\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38703\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__38712\,
            I => \N__38699\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__38709\,
            I => \N__38694\
        );

    \I__8633\ : Span4Mux_s1_v
    port map (
            O => \N__38706\,
            I => \N__38694\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38690\
        );

    \I__8631\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38687\
        );

    \I__8630\ : Span4Mux_h
    port map (
            O => \N__38699\,
            I => \N__38684\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__38694\,
            I => \N__38681\
        );

    \I__8628\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38678\
        );

    \I__8627\ : Sp12to4
    port map (
            O => \N__38690\,
            I => \N__38673\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38673\
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__38684\,
            I => rand_data_8
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__38681\,
            I => rand_data_8
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__38678\,
            I => rand_data_8
        );

    \I__8622\ : Odrv12
    port map (
            O => \N__38673\,
            I => rand_data_8
        );

    \I__8621\ : InMux
    port map (
            O => \N__38664\,
            I => \bfn_14_10_0_\
        );

    \I__8620\ : InMux
    port map (
            O => \N__38661\,
            I => \N__38657\
        );

    \I__8619\ : InMux
    port map (
            O => \N__38660\,
            I => \N__38654\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__38657\,
            I => \N__38651\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38646\
        );

    \I__8616\ : Span4Mux_s1_v
    port map (
            O => \N__38651\,
            I => \N__38643\
        );

    \I__8615\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38640\
        );

    \I__8614\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38636\
        );

    \I__8613\ : Span4Mux_s2_v
    port map (
            O => \N__38646\,
            I => \N__38633\
        );

    \I__8612\ : Span4Mux_h
    port map (
            O => \N__38643\,
            I => \N__38630\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__38640\,
            I => \N__38627\
        );

    \I__8610\ : InMux
    port map (
            O => \N__38639\,
            I => \N__38623\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__38636\,
            I => \N__38620\
        );

    \I__8608\ : Span4Mux_h
    port map (
            O => \N__38633\,
            I => \N__38617\
        );

    \I__8607\ : Span4Mux_v
    port map (
            O => \N__38630\,
            I => \N__38612\
        );

    \I__8606\ : Span4Mux_h
    port map (
            O => \N__38627\,
            I => \N__38612\
        );

    \I__8605\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38609\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__38623\,
            I => \N__38604\
        );

    \I__8603\ : Span4Mux_v
    port map (
            O => \N__38620\,
            I => \N__38604\
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__38617\,
            I => rand_data_9
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__38612\,
            I => rand_data_9
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__38609\,
            I => rand_data_9
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__38604\,
            I => rand_data_9
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__38595\,
            I => \N__38592\
        );

    \I__8597\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38589\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__38589\,
            I => \N__38585\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__38588\,
            I => \N__38582\
        );

    \I__8594\ : Span4Mux_v
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__8593\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38576\
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__38579\,
            I => rand_setpoint_9
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__38576\,
            I => rand_setpoint_9
        );

    \I__8590\ : InMux
    port map (
            O => \N__38571\,
            I => n16586
        );

    \I__8589\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38560\
        );

    \I__8587\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38557\
        );

    \I__8586\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38553\
        );

    \I__8585\ : Span4Mux_v
    port map (
            O => \N__38560\,
            I => \N__38549\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__38557\,
            I => \N__38546\
        );

    \I__8583\ : CascadeMux
    port map (
            O => \N__38556\,
            I => \N__38543\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__38553\,
            I => \N__38539\
        );

    \I__8581\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38536\
        );

    \I__8580\ : Span4Mux_h
    port map (
            O => \N__38549\,
            I => \N__38533\
        );

    \I__8579\ : Span4Mux_v
    port map (
            O => \N__38546\,
            I => \N__38530\
        );

    \I__8578\ : InMux
    port map (
            O => \N__38543\,
            I => \N__38527\
        );

    \I__8577\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38524\
        );

    \I__8576\ : Span12Mux_h
    port map (
            O => \N__38539\,
            I => \N__38519\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__38536\,
            I => \N__38519\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__38533\,
            I => rand_data_10
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__38530\,
            I => rand_data_10
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__38527\,
            I => rand_data_10
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__38524\,
            I => rand_data_10
        );

    \I__8570\ : Odrv12
    port map (
            O => \N__38519\,
            I => rand_data_10
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__38508\,
            I => \N__38504\
        );

    \I__8568\ : InMux
    port map (
            O => \N__38507\,
            I => \N__38501\
        );

    \I__8567\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38498\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__38501\,
            I => rand_setpoint_10
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__38498\,
            I => rand_setpoint_10
        );

    \I__8564\ : InMux
    port map (
            O => \N__38493\,
            I => n16587
        );

    \I__8563\ : InMux
    port map (
            O => \N__38490\,
            I => n16588
        );

    \I__8562\ : InMux
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__38484\,
            I => \N__38481\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__38481\,
            I => \N__38477\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__38480\,
            I => \N__38474\
        );

    \I__8558\ : Span4Mux_v
    port map (
            O => \N__38477\,
            I => \N__38471\
        );

    \I__8557\ : InMux
    port map (
            O => \N__38474\,
            I => \N__38468\
        );

    \I__8556\ : Odrv4
    port map (
            O => \N__38471\,
            I => rand_setpoint_12
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__38468\,
            I => rand_setpoint_12
        );

    \I__8554\ : InMux
    port map (
            O => \N__38463\,
            I => n16589
        );

    \I__8553\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38454\
        );

    \I__8552\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38454\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__38454\,
            I => \N__38451\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__38451\,
            I => \N__38446\
        );

    \I__8549\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38442\
        );

    \I__8548\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38438\
        );

    \I__8547\ : Span4Mux_h
    port map (
            O => \N__38446\,
            I => \N__38435\
        );

    \I__8546\ : InMux
    port map (
            O => \N__38445\,
            I => \N__38432\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__38442\,
            I => \N__38429\
        );

    \I__8544\ : InMux
    port map (
            O => \N__38441\,
            I => \N__38426\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__38438\,
            I => \N__38423\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__38435\,
            I => rand_data_13
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__38432\,
            I => rand_data_13
        );

    \I__8540\ : Odrv12
    port map (
            O => \N__38429\,
            I => rand_data_13
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__38426\,
            I => rand_data_13
        );

    \I__8538\ : Odrv12
    port map (
            O => \N__38423\,
            I => rand_data_13
        );

    \I__8537\ : InMux
    port map (
            O => \N__38412\,
            I => n16590
        );

    \I__8536\ : InMux
    port map (
            O => \N__38409\,
            I => n16575
        );

    \I__8535\ : InMux
    port map (
            O => \N__38406\,
            I => n16576
        );

    \I__8534\ : InMux
    port map (
            O => \N__38403\,
            I => n16577
        );

    \I__8533\ : InMux
    port map (
            O => \N__38400\,
            I => \N__38396\
        );

    \I__8532\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38393\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__38396\,
            I => \N__38389\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38385\
        );

    \I__8529\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38382\
        );

    \I__8528\ : Span4Mux_v
    port map (
            O => \N__38389\,
            I => \N__38378\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__38388\,
            I => \N__38375\
        );

    \I__8526\ : Span4Mux_v
    port map (
            O => \N__38385\,
            I => \N__38370\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__38382\,
            I => \N__38370\
        );

    \I__8524\ : InMux
    port map (
            O => \N__38381\,
            I => \N__38366\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__38378\,
            I => \N__38363\
        );

    \I__8522\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38360\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__38370\,
            I => \N__38357\
        );

    \I__8520\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38354\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__38366\,
            I => \N__38351\
        );

    \I__8518\ : Odrv4
    port map (
            O => \N__38363\,
            I => rand_data_0
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__38360\,
            I => rand_data_0
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__38357\,
            I => rand_data_0
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__38354\,
            I => rand_data_0
        );

    \I__8514\ : Odrv12
    port map (
            O => \N__38351\,
            I => rand_data_0
        );

    \I__8513\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__38337\,
            I => \N__38332\
        );

    \I__8511\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38329\
        );

    \I__8510\ : InMux
    port map (
            O => \N__38335\,
            I => \N__38326\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__38332\,
            I => \N__38321\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__38329\,
            I => \N__38321\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__38326\,
            I => \N__38317\
        );

    \I__8506\ : Span4Mux_v
    port map (
            O => \N__38321\,
            I => \N__38313\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__38320\,
            I => \N__38310\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__38317\,
            I => \N__38306\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38303\
        );

    \I__8502\ : Sp12to4
    port map (
            O => \N__38313\,
            I => \N__38300\
        );

    \I__8501\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38297\
        );

    \I__8500\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38294\
        );

    \I__8499\ : Sp12to4
    port map (
            O => \N__38306\,
            I => \N__38289\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__38303\,
            I => \N__38289\
        );

    \I__8497\ : Odrv12
    port map (
            O => \N__38300\,
            I => rand_data_1
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__38297\,
            I => rand_data_1
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__38294\,
            I => rand_data_1
        );

    \I__8494\ : Odrv12
    port map (
            O => \N__38289\,
            I => rand_data_1
        );

    \I__8493\ : InMux
    port map (
            O => \N__38280\,
            I => n16578
        );

    \I__8492\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38272\
        );

    \I__8491\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38268\
        );

    \I__8490\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38265\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__38272\,
            I => \N__38262\
        );

    \I__8488\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38258\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38255\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__38265\,
            I => \N__38252\
        );

    \I__8485\ : Sp12to4
    port map (
            O => \N__38262\,
            I => \N__38248\
        );

    \I__8484\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38245\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__38258\,
            I => \N__38242\
        );

    \I__8482\ : Span4Mux_h
    port map (
            O => \N__38255\,
            I => \N__38239\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__38252\,
            I => \N__38236\
        );

    \I__8480\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38233\
        );

    \I__8479\ : Span12Mux_h
    port map (
            O => \N__38248\,
            I => \N__38228\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38228\
        );

    \I__8477\ : Odrv12
    port map (
            O => \N__38242\,
            I => rand_data_2
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__38239\,
            I => rand_data_2
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__38236\,
            I => rand_data_2
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__38233\,
            I => rand_data_2
        );

    \I__8473\ : Odrv12
    port map (
            O => \N__38228\,
            I => rand_data_2
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__8471\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38211\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__38211\,
            I => \N__38208\
        );

    \I__8469\ : Span4Mux_h
    port map (
            O => \N__38208\,
            I => \N__38204\
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__38207\,
            I => \N__38201\
        );

    \I__8467\ : Sp12to4
    port map (
            O => \N__38204\,
            I => \N__38198\
        );

    \I__8466\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38195\
        );

    \I__8465\ : Odrv12
    port map (
            O => \N__38198\,
            I => rand_setpoint_2
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38195\,
            I => rand_setpoint_2
        );

    \I__8463\ : InMux
    port map (
            O => \N__38190\,
            I => n16579
        );

    \I__8462\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38183\
        );

    \I__8461\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38179\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__38183\,
            I => \N__38176\
        );

    \I__8459\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38171\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__38179\,
            I => \N__38168\
        );

    \I__8457\ : Span4Mux_v
    port map (
            O => \N__38176\,
            I => \N__38165\
        );

    \I__8456\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38161\
        );

    \I__8455\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38158\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__38171\,
            I => \N__38155\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__38168\,
            I => \N__38150\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__38165\,
            I => \N__38150\
        );

    \I__8451\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38147\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__38161\,
            I => \N__38144\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__38158\,
            I => rand_data_3
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__38155\,
            I => rand_data_3
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__38150\,
            I => rand_data_3
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__38147\,
            I => rand_data_3
        );

    \I__8445\ : Odrv12
    port map (
            O => \N__38144\,
            I => rand_data_3
        );

    \I__8444\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38126\
        );

    \I__8442\ : CascadeMux
    port map (
            O => \N__38129\,
            I => \N__38123\
        );

    \I__8441\ : Span4Mux_v
    port map (
            O => \N__38126\,
            I => \N__38120\
        );

    \I__8440\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38117\
        );

    \I__8439\ : Odrv4
    port map (
            O => \N__38120\,
            I => rand_setpoint_3
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__38117\,
            I => rand_setpoint_3
        );

    \I__8437\ : InMux
    port map (
            O => \N__38112\,
            I => n16580
        );

    \I__8436\ : InMux
    port map (
            O => \N__38109\,
            I => \N__38104\
        );

    \I__8435\ : InMux
    port map (
            O => \N__38108\,
            I => \N__38101\
        );

    \I__8434\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38098\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38091\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__38101\,
            I => \N__38091\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__38098\,
            I => \N__38091\
        );

    \I__8430\ : Span4Mux_v
    port map (
            O => \N__38091\,
            I => \N__38087\
        );

    \I__8429\ : CascadeMux
    port map (
            O => \N__38090\,
            I => \N__38084\
        );

    \I__8428\ : Sp12to4
    port map (
            O => \N__38087\,
            I => \N__38079\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38076\
        );

    \I__8426\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38073\
        );

    \I__8425\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38070\
        );

    \I__8424\ : Span12Mux_h
    port map (
            O => \N__38079\,
            I => \N__38065\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__38076\,
            I => \N__38065\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__38073\,
            I => rand_data_4
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__38070\,
            I => rand_data_4
        );

    \I__8420\ : Odrv12
    port map (
            O => \N__38065\,
            I => rand_data_4
        );

    \I__8419\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__38055\,
            I => \N__38052\
        );

    \I__8417\ : Span4Mux_h
    port map (
            O => \N__38052\,
            I => \N__38049\
        );

    \I__8416\ : Span4Mux_v
    port map (
            O => \N__38049\,
            I => \N__38045\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38042\
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__38045\,
            I => rand_setpoint_4
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38042\,
            I => rand_setpoint_4
        );

    \I__8412\ : InMux
    port map (
            O => \N__38037\,
            I => n16581
        );

    \I__8411\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38031\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__8409\ : Span4Mux_v
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__38025\,
            I => \N__38021\
        );

    \I__8407\ : InMux
    port map (
            O => \N__38024\,
            I => \N__38018\
        );

    \I__8406\ : Odrv4
    port map (
            O => \N__38021\,
            I => rand_setpoint_5
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__38018\,
            I => rand_setpoint_5
        );

    \I__8404\ : InMux
    port map (
            O => \N__38013\,
            I => n16582
        );

    \I__8403\ : InMux
    port map (
            O => \N__38010\,
            I => n16566
        );

    \I__8402\ : InMux
    port map (
            O => \N__38007\,
            I => n16567
        );

    \I__8401\ : InMux
    port map (
            O => \N__38004\,
            I => n16568
        );

    \I__8400\ : InMux
    port map (
            O => \N__38001\,
            I => n16569
        );

    \I__8399\ : InMux
    port map (
            O => \N__37998\,
            I => \bfn_14_8_0_\
        );

    \I__8398\ : InMux
    port map (
            O => \N__37995\,
            I => n16571
        );

    \I__8397\ : InMux
    port map (
            O => \N__37992\,
            I => n16572
        );

    \I__8396\ : InMux
    port map (
            O => \N__37989\,
            I => n16573
        );

    \I__8395\ : InMux
    port map (
            O => \N__37986\,
            I => n16574
        );

    \I__8394\ : InMux
    port map (
            O => \N__37983\,
            I => n16557
        );

    \I__8393\ : InMux
    port map (
            O => \N__37980\,
            I => n16558
        );

    \I__8392\ : InMux
    port map (
            O => \N__37977\,
            I => n16559
        );

    \I__8391\ : InMux
    port map (
            O => \N__37974\,
            I => n16560
        );

    \I__8390\ : InMux
    port map (
            O => \N__37971\,
            I => n16561
        );

    \I__8389\ : InMux
    port map (
            O => \N__37968\,
            I => \bfn_14_7_0_\
        );

    \I__8388\ : InMux
    port map (
            O => \N__37965\,
            I => n16563
        );

    \I__8387\ : InMux
    port map (
            O => \N__37962\,
            I => n16564
        );

    \I__8386\ : InMux
    port map (
            O => \N__37959\,
            I => n16565
        );

    \I__8385\ : InMux
    port map (
            O => \N__37956\,
            I => n16548
        );

    \I__8384\ : InMux
    port map (
            O => \N__37953\,
            I => n16549
        );

    \I__8383\ : InMux
    port map (
            O => \N__37950\,
            I => n16550
        );

    \I__8382\ : InMux
    port map (
            O => \N__37947\,
            I => n16551
        );

    \I__8381\ : InMux
    port map (
            O => \N__37944\,
            I => n16552
        );

    \I__8380\ : InMux
    port map (
            O => \N__37941\,
            I => n16553
        );

    \I__8379\ : InMux
    port map (
            O => \N__37938\,
            I => \bfn_14_6_0_\
        );

    \I__8378\ : InMux
    port map (
            O => \N__37935\,
            I => n16555
        );

    \I__8377\ : InMux
    port map (
            O => \N__37932\,
            I => n16556
        );

    \I__8376\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37923\
        );

    \I__8374\ : Span4Mux_s2_v
    port map (
            O => \N__37923\,
            I => \N__37920\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__37920\,
            I => \N__37917\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__37917\,
            I => \c0.n18681\
        );

    \I__8371\ : InMux
    port map (
            O => \N__37914\,
            I => \bfn_14_5_0_\
        );

    \I__8370\ : InMux
    port map (
            O => \N__37911\,
            I => n16547
        );

    \I__8369\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__37905\,
            I => \c0.n17783\
        );

    \I__8367\ : CascadeMux
    port map (
            O => \N__37902\,
            I => \c0.n15_adj_2414_cascade_\
        );

    \I__8366\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37896\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__37896\,
            I => \N__37893\
        );

    \I__8364\ : Span4Mux_s1_v
    port map (
            O => \N__37893\,
            I => \N__37890\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__37890\,
            I => \c0.data_out_frame2_20_1\
        );

    \I__8362\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__37884\,
            I => \N__37881\
        );

    \I__8360\ : Span4Mux_v
    port map (
            O => \N__37881\,
            I => \N__37878\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__37878\,
            I => \c0.n31\
        );

    \I__8358\ : CascadeMux
    port map (
            O => \N__37875\,
            I => \c0.n32_cascade_\
        );

    \I__8357\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37869\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__37869\,
            I => \N__37866\
        );

    \I__8355\ : Span12Mux_s2_v
    port map (
            O => \N__37866\,
            I => \N__37863\
        );

    \I__8354\ : Odrv12
    port map (
            O => \N__37863\,
            I => \c0.data_out_frame2_19_7\
        );

    \I__8353\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37855\
        );

    \I__8352\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37850\
        );

    \I__8351\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37850\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__37855\,
            I => \N__37847\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__37850\,
            I => \N__37844\
        );

    \I__8348\ : Span4Mux_s2_v
    port map (
            O => \N__37847\,
            I => \N__37839\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__37844\,
            I => \N__37836\
        );

    \I__8346\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37831\
        );

    \I__8345\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37831\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__37839\,
            I => \N__37828\
        );

    \I__8343\ : Odrv4
    port map (
            O => \N__37836\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__37831\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__37828\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__8340\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37818\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__8338\ : Odrv12
    port map (
            O => \N__37815\,
            I => \c0.n17777\
        );

    \I__8337\ : InMux
    port map (
            O => \N__37812\,
            I => \N__37809\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__37809\,
            I => \c0.n6_adj_2430\
        );

    \I__8335\ : CascadeMux
    port map (
            O => \N__37806\,
            I => \c0.n17777_cascade_\
        );

    \I__8334\ : InMux
    port map (
            O => \N__37803\,
            I => \N__37799\
        );

    \I__8333\ : InMux
    port map (
            O => \N__37802\,
            I => \N__37796\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__37799\,
            I => \N__37793\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__37796\,
            I => \N__37789\
        );

    \I__8330\ : Span4Mux_s3_v
    port map (
            O => \N__37793\,
            I => \N__37786\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__37792\,
            I => \N__37782\
        );

    \I__8328\ : Span4Mux_h
    port map (
            O => \N__37789\,
            I => \N__37779\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37776\
        );

    \I__8326\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37771\
        );

    \I__8325\ : InMux
    port map (
            O => \N__37782\,
            I => \N__37771\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__37779\,
            I => data_out_frame2_5_5
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__37776\,
            I => data_out_frame2_5_5
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__37771\,
            I => data_out_frame2_5_5
        );

    \I__8321\ : CascadeMux
    port map (
            O => \N__37764\,
            I => \c0.n10617_cascade_\
        );

    \I__8320\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37758\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__37758\,
            I => \N__37755\
        );

    \I__8318\ : Span4Mux_s2_v
    port map (
            O => \N__37755\,
            I => \N__37751\
        );

    \I__8317\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37748\
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__37751\,
            I => \c0.n17765\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__37748\,
            I => \c0.n17765\
        );

    \I__8314\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37737\
        );

    \I__8313\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37734\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__37741\,
            I => \N__37731\
        );

    \I__8311\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37728\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37725\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37722\
        );

    \I__8308\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37718\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37715\
        );

    \I__8306\ : Span4Mux_s2_v
    port map (
            O => \N__37725\,
            I => \N__37710\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__37722\,
            I => \N__37710\
        );

    \I__8304\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37707\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__37718\,
            I => \N__37702\
        );

    \I__8302\ : Span4Mux_h
    port map (
            O => \N__37715\,
            I => \N__37702\
        );

    \I__8301\ : Span4Mux_h
    port map (
            O => \N__37710\,
            I => \N__37699\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37707\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__37702\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__37699\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__37692\,
            I => \c0.n18759_cascade_\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__8295\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37683\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__37683\,
            I => \N__37680\
        );

    \I__8293\ : Span4Mux_s0_v
    port map (
            O => \N__37680\,
            I => \N__37676\
        );

    \I__8292\ : CascadeMux
    port map (
            O => \N__37679\,
            I => \N__37672\
        );

    \I__8291\ : Span4Mux_v
    port map (
            O => \N__37676\,
            I => \N__37668\
        );

    \I__8290\ : InMux
    port map (
            O => \N__37675\,
            I => \N__37663\
        );

    \I__8289\ : InMux
    port map (
            O => \N__37672\,
            I => \N__37663\
        );

    \I__8288\ : InMux
    port map (
            O => \N__37671\,
            I => \N__37660\
        );

    \I__8287\ : Odrv4
    port map (
            O => \N__37668\,
            I => data_out_frame2_6_0
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__37663\,
            I => data_out_frame2_6_0
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__37660\,
            I => data_out_frame2_6_0
        );

    \I__8284\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__37650\,
            I => \N__37647\
        );

    \I__8282\ : Odrv12
    port map (
            O => \N__37647\,
            I => \c0.n10920\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__37644\,
            I => \c0.n17783_cascade_\
        );

    \I__8280\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37638\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__37638\,
            I => \N__37634\
        );

    \I__8278\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37631\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__37634\,
            I => \c0.n10849\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__37631\,
            I => \c0.n10849\
        );

    \I__8275\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37623\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37619\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__37622\,
            I => \N__37616\
        );

    \I__8272\ : Span4Mux_s1_v
    port map (
            O => \N__37619\,
            I => \N__37613\
        );

    \I__8271\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37610\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__37613\,
            I => \c0.n17859\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__37610\,
            I => \c0.n17859\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__37605\,
            I => \c0.n15_cascade_\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__37602\,
            I => \N__37599\
        );

    \I__8266\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37596\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__8263\ : Odrv4
    port map (
            O => \N__37590\,
            I => \c0.data_out_frame2_19_0\
        );

    \I__8262\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37580\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__37583\,
            I => \N__37577\
        );

    \I__8259\ : Sp12to4
    port map (
            O => \N__37580\,
            I => \N__37574\
        );

    \I__8258\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37571\
        );

    \I__8257\ : Span12Mux_s2_v
    port map (
            O => \N__37574\,
            I => \N__37566\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__37571\,
            I => \N__37566\
        );

    \I__8255\ : Odrv12
    port map (
            O => \N__37566\,
            I => \c0.n10688\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__37563\,
            I => \c0.n10813_cascade_\
        );

    \I__8253\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37556\
        );

    \I__8252\ : InMux
    port map (
            O => \N__37559\,
            I => \N__37553\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__37556\,
            I => \N__37550\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__37553\,
            I => \c0.n10577\
        );

    \I__8249\ : Odrv4
    port map (
            O => \N__37550\,
            I => \c0.n10577\
        );

    \I__8248\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37541\
        );

    \I__8247\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37538\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37529\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37529\
        );

    \I__8244\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37526\
        );

    \I__8243\ : InMux
    port map (
            O => \N__37536\,
            I => \N__37523\
        );

    \I__8242\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37518\
        );

    \I__8241\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37518\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__37529\,
            I => \N__37515\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__37526\,
            I => \N__37512\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__37523\,
            I => data_out_6_0
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__37518\,
            I => data_out_6_0
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__37515\,
            I => data_out_6_0
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__37512\,
            I => data_out_6_0
        );

    \I__8234\ : CascadeMux
    port map (
            O => \N__37503\,
            I => \N__37500\
        );

    \I__8233\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__37497\,
            I => \c0.n10680\
        );

    \I__8231\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37491\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__37491\,
            I => \c0.n17816\
        );

    \I__8229\ : CascadeMux
    port map (
            O => \N__37488\,
            I => \c0.n10680_cascade_\
        );

    \I__8228\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37479\
        );

    \I__8227\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37476\
        );

    \I__8226\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37473\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37470\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37464\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37464\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37461\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37470\,
            I => \N__37458\
        );

    \I__8220\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37455\
        );

    \I__8219\ : Span4Mux_v
    port map (
            O => \N__37464\,
            I => \N__37452\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__37461\,
            I => \c0.data_out_5_5\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__37458\,
            I => \c0.data_out_5_5\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__37455\,
            I => \c0.data_out_5_5\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__37452\,
            I => \c0.data_out_5_5\
        );

    \I__8214\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37438\
        );

    \I__8213\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37435\
        );

    \I__8212\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37430\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__37438\,
            I => \N__37427\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__37435\,
            I => \N__37424\
        );

    \I__8209\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37419\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37419\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37412\
        );

    \I__8206\ : Span4Mux_v
    port map (
            O => \N__37427\,
            I => \N__37412\
        );

    \I__8205\ : Span4Mux_v
    port map (
            O => \N__37424\,
            I => \N__37412\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__37419\,
            I => data_out_8_6
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__37412\,
            I => data_out_8_6
        );

    \I__8202\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37404\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37400\
        );

    \I__8200\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37397\
        );

    \I__8199\ : Span4Mux_v
    port map (
            O => \N__37400\,
            I => \N__37394\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__37397\,
            I => \N__37391\
        );

    \I__8197\ : Span4Mux_h
    port map (
            O => \N__37394\,
            I => \N__37383\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__37391\,
            I => \N__37383\
        );

    \I__8195\ : InMux
    port map (
            O => \N__37390\,
            I => \N__37378\
        );

    \I__8194\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37378\
        );

    \I__8193\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37375\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__37383\,
            I => data_out_8_5
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__37378\,
            I => data_out_8_5
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__37375\,
            I => data_out_8_5
        );

    \I__8189\ : CascadeMux
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37358\
        );

    \I__8186\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37355\
        );

    \I__8185\ : Span4Mux_v
    port map (
            O => \N__37358\,
            I => \N__37352\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37349\
        );

    \I__8183\ : Span4Mux_v
    port map (
            O => \N__37352\,
            I => \N__37346\
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__37349\,
            I => \c0.n17771\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__37346\,
            I => \c0.n17771\
        );

    \I__8180\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37337\
        );

    \I__8179\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37332\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37329\
        );

    \I__8177\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37326\
        );

    \I__8176\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37323\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__37332\,
            I => \N__37320\
        );

    \I__8174\ : Span4Mux_v
    port map (
            O => \N__37329\,
            I => \N__37317\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__37326\,
            I => \N__37314\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__37323\,
            I => \N__37310\
        );

    \I__8171\ : Span4Mux_v
    port map (
            O => \N__37320\,
            I => \N__37307\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__37317\,
            I => \N__37304\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__37314\,
            I => \N__37301\
        );

    \I__8168\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37298\
        );

    \I__8167\ : Span4Mux_h
    port map (
            O => \N__37310\,
            I => \N__37295\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__37307\,
            I => data_out_5_1
        );

    \I__8165\ : Odrv4
    port map (
            O => \N__37304\,
            I => data_out_5_1
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__37301\,
            I => data_out_5_1
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__37298\,
            I => data_out_5_1
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__37295\,
            I => data_out_5_1
        );

    \I__8161\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37279\
        );

    \I__8160\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37272\
        );

    \I__8159\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37269\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__37279\,
            I => \N__37266\
        );

    \I__8157\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37261\
        );

    \I__8156\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37261\
        );

    \I__8155\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37256\
        );

    \I__8154\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37256\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__37272\,
            I => \N__37253\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__37269\,
            I => \N__37250\
        );

    \I__8151\ : Span4Mux_v
    port map (
            O => \N__37266\,
            I => \N__37246\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__37261\,
            I => \N__37243\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37240\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__37253\,
            I => \N__37235\
        );

    \I__8147\ : Span4Mux_h
    port map (
            O => \N__37250\,
            I => \N__37235\
        );

    \I__8146\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37232\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__37246\,
            I => \c0.data_out_5_4\
        );

    \I__8144\ : Odrv12
    port map (
            O => \N__37243\,
            I => \c0.data_out_5_4\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__37240\,
            I => \c0.data_out_5_4\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__37235\,
            I => \c0.data_out_5_4\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__37232\,
            I => \c0.data_out_5_4\
        );

    \I__8140\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37217\
        );

    \I__8139\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37214\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37209\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37206\
        );

    \I__8136\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37203\
        );

    \I__8135\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37200\
        );

    \I__8134\ : Span12Mux_h
    port map (
            O => \N__37209\,
            I => \N__37193\
        );

    \I__8133\ : Span12Mux_h
    port map (
            O => \N__37206\,
            I => \N__37193\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__37203\,
            I => \N__37193\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__37200\,
            I => data_out_frame2_13_2
        );

    \I__8130\ : Odrv12
    port map (
            O => \N__37193\,
            I => data_out_frame2_13_2
        );

    \I__8129\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37184\
        );

    \I__8128\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37180\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__37184\,
            I => \N__37175\
        );

    \I__8126\ : InMux
    port map (
            O => \N__37183\,
            I => \N__37172\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__37180\,
            I => \N__37169\
        );

    \I__8124\ : InMux
    port map (
            O => \N__37179\,
            I => \N__37166\
        );

    \I__8123\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37163\
        );

    \I__8122\ : Span4Mux_h
    port map (
            O => \N__37175\,
            I => \N__37160\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37157\
        );

    \I__8120\ : Span4Mux_s0_v
    port map (
            O => \N__37169\,
            I => \N__37154\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__37166\,
            I => \N__37151\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__37163\,
            I => data_out_frame2_16_0
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__37160\,
            I => data_out_frame2_16_0
        );

    \I__8116\ : Odrv4
    port map (
            O => \N__37157\,
            I => data_out_frame2_16_0
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__37154\,
            I => data_out_frame2_16_0
        );

    \I__8114\ : Odrv12
    port map (
            O => \N__37151\,
            I => data_out_frame2_16_0
        );

    \I__8113\ : InMux
    port map (
            O => \N__37140\,
            I => \N__37135\
        );

    \I__8112\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37130\
        );

    \I__8111\ : InMux
    port map (
            O => \N__37138\,
            I => \N__37130\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__37135\,
            I => \N__37125\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37122\
        );

    \I__8108\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37119\
        );

    \I__8107\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37116\
        );

    \I__8106\ : Span4Mux_h
    port map (
            O => \N__37125\,
            I => \N__37113\
        );

    \I__8105\ : Span4Mux_h
    port map (
            O => \N__37122\,
            I => \N__37110\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__37119\,
            I => data_out_frame2_8_6
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__37116\,
            I => data_out_frame2_8_6
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__37113\,
            I => data_out_frame2_8_6
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__37110\,
            I => data_out_frame2_8_6
        );

    \I__8100\ : InMux
    port map (
            O => \N__37101\,
            I => \N__37098\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__37098\,
            I => \N__37094\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37089\
        );

    \I__8097\ : Span4Mux_h
    port map (
            O => \N__37094\,
            I => \N__37086\
        );

    \I__8096\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37083\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37080\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__37089\,
            I => data_out_10_6
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__37086\,
            I => data_out_10_6
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__37083\,
            I => data_out_10_6
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__37080\,
            I => data_out_10_6
        );

    \I__8090\ : InMux
    port map (
            O => \N__37071\,
            I => \N__37067\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37070\,
            I => \N__37063\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__37067\,
            I => \N__37060\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37066\,
            I => \N__37057\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__37063\,
            I => \N__37052\
        );

    \I__8085\ : Span4Mux_v
    port map (
            O => \N__37060\,
            I => \N__37052\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__37057\,
            I => \c0.data_out_7_2\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__37052\,
            I => \c0.data_out_7_2\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__37047\,
            I => \N__37044\
        );

    \I__8081\ : InMux
    port map (
            O => \N__37044\,
            I => \N__37040\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37037\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37040\,
            I => \N__37031\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37031\
        );

    \I__8077\ : CascadeMux
    port map (
            O => \N__37036\,
            I => \N__37028\
        );

    \I__8076\ : Span4Mux_v
    port map (
            O => \N__37031\,
            I => \N__37025\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__8074\ : Odrv4
    port map (
            O => \N__37025\,
            I => \c0.data_out_9_1\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37022\,
            I => \c0.data_out_9_1\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__37014\,
            I => \N__37011\
        );

    \I__8070\ : Span4Mux_h
    port map (
            O => \N__37011\,
            I => \N__37008\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__37008\,
            I => \c0.n17730\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37005\,
            I => \N__37001\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37004\,
            I => \N__36998\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__37001\,
            I => \c0.n17835\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__36998\,
            I => \c0.n17835\
        );

    \I__8064\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__36990\,
            I => \N__36986\
        );

    \I__8062\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36983\
        );

    \I__8061\ : Span12Mux_v
    port map (
            O => \N__36986\,
            I => \N__36980\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__8059\ : Odrv12
    port map (
            O => \N__36980\,
            I => \c0.n17844\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__36977\,
            I => \c0.n17844\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__36972\,
            I => \c0.n17730_cascade_\
        );

    \I__8056\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36965\
        );

    \I__8055\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36962\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__36965\,
            I => \N__36959\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__36962\,
            I => n17758
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__36959\,
            I => n17758
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__36954\,
            I => \c0.n14_adj_2363_cascade_\
        );

    \I__8050\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36948\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__36945\,
            I => \c0.n13\
        );

    \I__8047\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36939\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__36939\,
            I => \N__36934\
        );

    \I__8045\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36930\
        );

    \I__8044\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36927\
        );

    \I__8043\ : Span4Mux_h
    port map (
            O => \N__36934\,
            I => \N__36924\
        );

    \I__8042\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36921\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__36930\,
            I => \c0.data_out_9_3\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__36927\,
            I => \c0.data_out_9_3\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__36924\,
            I => \c0.data_out_9_3\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__36921\,
            I => \c0.data_out_9_3\
        );

    \I__8037\ : CascadeMux
    port map (
            O => \N__36912\,
            I => \c0.n17816_cascade_\
        );

    \I__8036\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36905\
        );

    \I__8035\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36902\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__36905\,
            I => \c0.n17877\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__36902\,
            I => \c0.n17877\
        );

    \I__8032\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36894\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__36894\,
            I => \c0.n12\
        );

    \I__8030\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36887\
        );

    \I__8029\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36884\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__36887\,
            I => \N__36881\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36878\
        );

    \I__8026\ : Span4Mux_h
    port map (
            O => \N__36881\,
            I => \N__36875\
        );

    \I__8025\ : Odrv4
    port map (
            O => \N__36878\,
            I => \c0.n17786\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__36875\,
            I => \c0.n17786\
        );

    \I__8023\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36867\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36864\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__36864\,
            I => \N__36861\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__36861\,
            I => \c0.n18184\
        );

    \I__8019\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36855\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__36855\,
            I => \N__36850\
        );

    \I__8017\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36847\
        );

    \I__8016\ : InMux
    port map (
            O => \N__36853\,
            I => \N__36844\
        );

    \I__8015\ : Span4Mux_h
    port map (
            O => \N__36850\,
            I => \N__36841\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36838\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__36844\,
            I => \c0.data_out_7_1\
        );

    \I__8012\ : Odrv4
    port map (
            O => \N__36841\,
            I => \c0.data_out_7_1\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__36838\,
            I => \c0.data_out_7_1\
        );

    \I__8010\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36824\
        );

    \I__8009\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36824\
        );

    \I__8008\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36821\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36818\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__36821\,
            I => \N__36815\
        );

    \I__8005\ : Odrv4
    port map (
            O => \N__36818\,
            I => \c0.n10537\
        );

    \I__8004\ : Odrv4
    port map (
            O => \N__36815\,
            I => \c0.n10537\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__36810\,
            I => \c0.n18238_cascade_\
        );

    \I__8002\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36804\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36799\
        );

    \I__8000\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36794\
        );

    \I__7999\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36794\
        );

    \I__7998\ : Span4Mux_v
    port map (
            O => \N__36799\,
            I => \N__36791\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__36794\,
            I => \c0.data_out_6_4\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__36791\,
            I => \c0.data_out_6_4\
        );

    \I__7995\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36783\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__36783\,
            I => \N__36780\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__36780\,
            I => \c0.n6_adj_2276\
        );

    \I__7992\ : InMux
    port map (
            O => \N__36777\,
            I => \N__36773\
        );

    \I__7991\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36770\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__36773\,
            I => \N__36766\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36763\
        );

    \I__7988\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36760\
        );

    \I__7987\ : Span4Mux_h
    port map (
            O => \N__36766\,
            I => \N__36757\
        );

    \I__7986\ : Span12Mux_v
    port map (
            O => \N__36763\,
            I => \N__36754\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__36760\,
            I => \c0.data_out_6_7\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__36757\,
            I => \c0.data_out_6_7\
        );

    \I__7983\ : Odrv12
    port map (
            O => \N__36754\,
            I => \c0.data_out_6_7\
        );

    \I__7982\ : InMux
    port map (
            O => \N__36747\,
            I => \N__36742\
        );

    \I__7981\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36739\
        );

    \I__7980\ : InMux
    port map (
            O => \N__36745\,
            I => \N__36736\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__36742\,
            I => \N__36728\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__36739\,
            I => \N__36728\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__36736\,
            I => \N__36728\
        );

    \I__7976\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36725\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__36728\,
            I => \N__36722\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__36725\,
            I => \c0.data_out_6_5\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__36722\,
            I => \c0.data_out_6_5\
        );

    \I__7972\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36713\
        );

    \I__7971\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36710\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__36713\,
            I => \N__36705\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__36710\,
            I => \N__36702\
        );

    \I__7968\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36699\
        );

    \I__7967\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36696\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__36705\,
            I => \N__36689\
        );

    \I__7965\ : Span4Mux_v
    port map (
            O => \N__36702\,
            I => \N__36689\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__36699\,
            I => \N__36689\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__36696\,
            I => data_out_8_4
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__36689\,
            I => data_out_8_4
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__36684\,
            I => \N__36681\
        );

    \I__7960\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__36678\,
            I => \c0.n17745\
        );

    \I__7958\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36672\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36669\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__36669\,
            I => \c0.n10542\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__36666\,
            I => \c0.n17745_cascade_\
        );

    \I__7954\ : CascadeMux
    port map (
            O => \N__36663\,
            I => \N__36660\
        );

    \I__7953\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36656\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__36659\,
            I => \N__36653\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36650\
        );

    \I__7950\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36647\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__36650\,
            I => \N__36641\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__36647\,
            I => \N__36641\
        );

    \I__7947\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36638\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36635\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__36638\,
            I => \c0.data_out_10_7\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__36635\,
            I => \c0.data_out_10_7\
        );

    \I__7943\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36627\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__36627\,
            I => \N__36620\
        );

    \I__7941\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36615\
        );

    \I__7940\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36615\
        );

    \I__7939\ : InMux
    port map (
            O => \N__36624\,
            I => \N__36610\
        );

    \I__7938\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36610\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__36620\,
            I => data_out_8_3
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__36615\,
            I => data_out_8_3
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__36610\,
            I => data_out_8_3
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__36603\,
            I => \N__36600\
        );

    \I__7933\ : InMux
    port map (
            O => \N__36600\,
            I => \N__36597\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__36597\,
            I => \N__36594\
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__36594\,
            I => \c0.n8_adj_2219\
        );

    \I__7930\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36588\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36585\
        );

    \I__7928\ : Span4Mux_h
    port map (
            O => \N__36585\,
            I => \N__36581\
        );

    \I__7927\ : InMux
    port map (
            O => \N__36584\,
            I => \N__36578\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__36581\,
            I => \N__36575\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__36578\,
            I => data_out_0_3
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__36575\,
            I => data_out_0_3
        );

    \I__7923\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36567\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__36567\,
            I => \N__36564\
        );

    \I__7921\ : Span4Mux_h
    port map (
            O => \N__36564\,
            I => \N__36561\
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__36561\,
            I => \c0.n18376\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__36558\,
            I => \N__36554\
        );

    \I__7918\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36550\
        );

    \I__7917\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36547\
        );

    \I__7916\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36544\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__36550\,
            I => \N__36541\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__36547\,
            I => \N__36536\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__36544\,
            I => \N__36533\
        );

    \I__7912\ : Span4Mux_h
    port map (
            O => \N__36541\,
            I => \N__36530\
        );

    \I__7911\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36525\
        );

    \I__7910\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36525\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__36536\,
            I => data_out_8_2
        );

    \I__7908\ : Odrv4
    port map (
            O => \N__36533\,
            I => data_out_8_2
        );

    \I__7907\ : Odrv4
    port map (
            O => \N__36530\,
            I => data_out_8_2
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__36525\,
            I => data_out_8_2
        );

    \I__7905\ : CEMux
    port map (
            O => \N__36516\,
            I => \N__36513\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__36513\,
            I => \N__36509\
        );

    \I__7903\ : CEMux
    port map (
            O => \N__36512\,
            I => \N__36506\
        );

    \I__7902\ : Span4Mux_v
    port map (
            O => \N__36509\,
            I => \N__36503\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36500\
        );

    \I__7900\ : Span4Mux_h
    port map (
            O => \N__36503\,
            I => \N__36495\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__36500\,
            I => \N__36495\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__36495\,
            I => \c0.n11056\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__36492\,
            I => \c0.n18199_cascade_\
        );

    \I__7896\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36486\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36482\
        );

    \I__7894\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__7893\ : Span4Mux_v
    port map (
            O => \N__36482\,
            I => \N__36476\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36473\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__36476\,
            I => \N__36468\
        );

    \I__7890\ : Span4Mux_v
    port map (
            O => \N__36473\,
            I => \N__36468\
        );

    \I__7889\ : Odrv4
    port map (
            O => \N__36468\,
            I => \c0.n17832\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__36465\,
            I => \c0.n18242_cascade_\
        );

    \I__7887\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36459\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__36459\,
            I => \N__36455\
        );

    \I__7885\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36452\
        );

    \I__7884\ : Span4Mux_v
    port map (
            O => \N__36455\,
            I => \N__36449\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__36452\,
            I => \c0.data_out_6_6\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__36449\,
            I => \c0.data_out_6_6\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__7880\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36438\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__36438\,
            I => \c0.n5\
        );

    \I__7878\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__36432\,
            I => \c0.n18247\
        );

    \I__7876\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36423\
        );

    \I__7875\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36420\
        );

    \I__7874\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36417\
        );

    \I__7873\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36414\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36407\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__36420\,
            I => \N__36407\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__36417\,
            I => \N__36407\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__36414\,
            I => data_out_frame2_15_3
        );

    \I__7868\ : Odrv12
    port map (
            O => \N__36407\,
            I => data_out_frame2_15_3
        );

    \I__7867\ : CascadeMux
    port map (
            O => \N__36402\,
            I => \c0.n6_adj_2422_cascade_\
        );

    \I__7866\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36393\
        );

    \I__7865\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36393\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__36393\,
            I => data_out_frame2_18_4
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__36390\,
            I => \c0.n10870_cascade_\
        );

    \I__7862\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36384\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__36384\,
            I => \N__36381\
        );

    \I__7860\ : Span4Mux_v
    port map (
            O => \N__36381\,
            I => \N__36378\
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__36378\,
            I => \c0.n27_adj_2428\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__36375\,
            I => \N__36372\
        );

    \I__7857\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36369\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__36369\,
            I => \c0.n5_adj_2274\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__36366\,
            I => \c0.n18879_cascade_\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__36363\,
            I => \N__36360\
        );

    \I__7853\ : InMux
    port map (
            O => \N__36360\,
            I => \N__36357\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__36357\,
            I => \N__36354\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__36354\,
            I => \N__36351\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__36351\,
            I => \c0.n10852\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__36348\,
            I => \N__36345\
        );

    \I__7848\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36342\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N__36339\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__36339\,
            I => \N__36336\
        );

    \I__7845\ : Span4Mux_h
    port map (
            O => \N__36336\,
            I => \N__36332\
        );

    \I__7844\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36329\
        );

    \I__7843\ : IoSpan4Mux
    port map (
            O => \N__36332\,
            I => \N__36326\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36323\
        );

    \I__7841\ : Span4Mux_s1_v
    port map (
            O => \N__36326\,
            I => \N__36320\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__36323\,
            I => \c0.n10867\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__36320\,
            I => \c0.n10867\
        );

    \I__7838\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36310\
        );

    \I__7837\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36307\
        );

    \I__7836\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36303\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__36310\,
            I => \N__36300\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__36307\,
            I => \N__36297\
        );

    \I__7833\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36294\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__36303\,
            I => data_out_frame2_8_5
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__36300\,
            I => data_out_frame2_8_5
        );

    \I__7830\ : Odrv4
    port map (
            O => \N__36297\,
            I => data_out_frame2_8_5
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__36294\,
            I => data_out_frame2_8_5
        );

    \I__7828\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36282\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__36282\,
            I => \c0.n14_adj_2447\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__7825\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36273\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__36273\,
            I => \N__36270\
        );

    \I__7823\ : Span12Mux_v
    port map (
            O => \N__36270\,
            I => \N__36267\
        );

    \I__7822\ : Odrv12
    port map (
            O => \N__36267\,
            I => \c0.data_out_frame2_19_4\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__36264\,
            I => \N__36261\
        );

    \I__7820\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36258\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__36258\,
            I => \c0.n10_adj_2440\
        );

    \I__7818\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36252\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__36252\,
            I => \N__36249\
        );

    \I__7816\ : Span4Mux_s2_v
    port map (
            O => \N__36249\,
            I => \N__36246\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__36246\,
            I => \c0.n6_adj_2357\
        );

    \I__7814\ : InMux
    port map (
            O => \N__36243\,
            I => \N__36240\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__36240\,
            I => \N__36236\
        );

    \I__7812\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36233\
        );

    \I__7811\ : Odrv12
    port map (
            O => \N__36236\,
            I => \c0.n10864\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__36233\,
            I => \c0.n10864\
        );

    \I__7809\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36224\
        );

    \I__7808\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36221\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36217\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__36221\,
            I => \N__36213\
        );

    \I__7805\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36210\
        );

    \I__7804\ : Span4Mux_h
    port map (
            O => \N__36217\,
            I => \N__36207\
        );

    \I__7803\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36204\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__36213\,
            I => \N__36201\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__36210\,
            I => data_out_frame2_6_4
        );

    \I__7800\ : Odrv4
    port map (
            O => \N__36207\,
            I => data_out_frame2_6_4
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__36204\,
            I => data_out_frame2_6_4
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__36201\,
            I => data_out_frame2_6_4
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__36192\,
            I => \c0.n10720_cascade_\
        );

    \I__7796\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36186\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__36180\
        );

    \I__7794\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36177\
        );

    \I__7793\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36174\
        );

    \I__7792\ : InMux
    port map (
            O => \N__36183\,
            I => \N__36171\
        );

    \I__7791\ : Span4Mux_h
    port map (
            O => \N__36180\,
            I => \N__36168\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36165\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__36174\,
            I => \N__36162\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__36171\,
            I => data_out_frame2_10_2
        );

    \I__7787\ : Odrv4
    port map (
            O => \N__36168\,
            I => data_out_frame2_10_2
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__36165\,
            I => data_out_frame2_10_2
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__36162\,
            I => data_out_frame2_10_2
        );

    \I__7784\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36150\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__36150\,
            I => \N__36146\
        );

    \I__7782\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36143\
        );

    \I__7781\ : Odrv4
    port map (
            O => \N__36146\,
            I => \c0.n10819\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__36143\,
            I => \c0.n10819\
        );

    \I__7779\ : InMux
    port map (
            O => \N__36138\,
            I => \N__36135\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36131\
        );

    \I__7777\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36128\
        );

    \I__7776\ : Span12Mux_s1_v
    port map (
            O => \N__36131\,
            I => \N__36125\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__36128\,
            I => \N__36122\
        );

    \I__7774\ : Odrv12
    port map (
            O => \N__36125\,
            I => \c0.n17886\
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__36122\,
            I => \c0.n17886\
        );

    \I__7772\ : InMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36111\
        );

    \I__7770\ : Odrv12
    port map (
            O => \N__36111\,
            I => \c0.n20_adj_2442\
        );

    \I__7769\ : CascadeMux
    port map (
            O => \N__36108\,
            I => \c0.n16_cascade_\
        );

    \I__7768\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36101\
        );

    \I__7767\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36098\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__36101\,
            I => \N__36093\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__36098\,
            I => \N__36093\
        );

    \I__7764\ : Span4Mux_s3_v
    port map (
            O => \N__36093\,
            I => \N__36090\
        );

    \I__7763\ : Odrv4
    port map (
            O => \N__36090\,
            I => \c0.n17795\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__7761\ : InMux
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__36081\,
            I => \N__36078\
        );

    \I__7759\ : Span4Mux_h
    port map (
            O => \N__36078\,
            I => \N__36075\
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__36075\,
            I => \c0.data_out_frame2_19_5\
        );

    \I__7757\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36063\
        );

    \I__7756\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36063\
        );

    \I__7755\ : InMux
    port map (
            O => \N__36070\,
            I => \N__36063\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__36063\,
            I => \c0.n10839\
        );

    \I__7753\ : InMux
    port map (
            O => \N__36060\,
            I => \N__36057\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__36057\,
            I => \N__36054\
        );

    \I__7751\ : Odrv4
    port map (
            O => \N__36054\,
            I => \c0.n10890\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36046\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36043\
        );

    \I__7748\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36040\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36036\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__36043\,
            I => \N__36033\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__36040\,
            I => \N__36030\
        );

    \I__7744\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36027\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__36036\,
            I => \N__36024\
        );

    \I__7742\ : Span4Mux_s3_v
    port map (
            O => \N__36033\,
            I => \N__36019\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__36030\,
            I => \N__36019\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__36027\,
            I => data_out_frame2_10_5
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__36024\,
            I => data_out_frame2_10_5
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__36019\,
            I => data_out_frame2_10_5
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__36012\,
            I => \N__36008\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36011\,
            I => \N__36005\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36008\,
            I => \N__36002\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__36005\,
            I => \N__35999\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__36002\,
            I => \N__35996\
        );

    \I__7732\ : Span4Mux_v
    port map (
            O => \N__35999\,
            I => \N__35993\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__35996\,
            I => \c0.n10816\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__35993\,
            I => \c0.n10816\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__35988\,
            I => \c0.n12_adj_2446_cascade_\
        );

    \I__7728\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35981\
        );

    \I__7727\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35976\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__35981\,
            I => \N__35973\
        );

    \I__7725\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35968\
        );

    \I__7724\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35968\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__35976\,
            I => data_out_frame2_15_1
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__35973\,
            I => data_out_frame2_15_1
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__35968\,
            I => data_out_frame2_15_1
        );

    \I__7720\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35958\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__35958\,
            I => \N__35955\
        );

    \I__7718\ : Span4Mux_s0_v
    port map (
            O => \N__35955\,
            I => \N__35952\
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__35952\,
            I => \c0.n10829\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__35949\,
            I => \c0.n10890_cascade_\
        );

    \I__7715\ : InMux
    port map (
            O => \N__35946\,
            I => \N__35943\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__35943\,
            I => \N__35940\
        );

    \I__7713\ : Span4Mux_h
    port map (
            O => \N__35940\,
            I => \N__35937\
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__35937\,
            I => \c0.n17_adj_2449\
        );

    \I__7711\ : CascadeMux
    port map (
            O => \N__35934\,
            I => \c0.n16_adj_2448_cascade_\
        );

    \I__7710\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35927\
        );

    \I__7709\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35924\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35919\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35919\
        );

    \I__7706\ : Span4Mux_s1_v
    port map (
            O => \N__35919\,
            I => \N__35916\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__35916\,
            I => \c0.n17911\
        );

    \I__7704\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35910\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__35910\,
            I => \c0.n15_adj_2445\
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__35907\,
            I => \c0.n14_adj_2444_cascade_\
        );

    \I__7701\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35901\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__35901\,
            I => \N__35894\
        );

    \I__7699\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35889\
        );

    \I__7698\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35889\
        );

    \I__7697\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35884\
        );

    \I__7696\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35884\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__35894\,
            I => data_out_frame2_16_1
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__35889\,
            I => data_out_frame2_16_1
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__35884\,
            I => data_out_frame2_16_1
        );

    \I__7692\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35874\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__35874\,
            I => \N__35871\
        );

    \I__7690\ : Odrv12
    port map (
            O => \N__35871\,
            I => \c0.data_out_frame2_20_5\
        );

    \I__7689\ : CascadeMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__7688\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__35862\,
            I => \c0.n16_adj_2358\
        );

    \I__7686\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35854\
        );

    \I__7685\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35847\
        );

    \I__7684\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35847\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35844\
        );

    \I__7682\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35841\
        );

    \I__7681\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35838\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35835\
        );

    \I__7679\ : Span4Mux_v
    port map (
            O => \N__35844\,
            I => \N__35830\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__35841\,
            I => \N__35830\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__35838\,
            I => \c0.data_out_7_4\
        );

    \I__7676\ : Odrv12
    port map (
            O => \N__35835\,
            I => \c0.data_out_7_4\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__35830\,
            I => \c0.data_out_7_4\
        );

    \I__7674\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35817\
        );

    \I__7673\ : InMux
    port map (
            O => \N__35822\,
            I => \N__35817\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__35817\,
            I => data_out_3_2
        );

    \I__7671\ : CascadeMux
    port map (
            O => \N__35814\,
            I => \N__35811\
        );

    \I__7670\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35805\
        );

    \I__7669\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35805\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__35805\,
            I => \c0.data_out_1_2\
        );

    \I__7667\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35799\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__35799\,
            I => \N__35796\
        );

    \I__7665\ : Odrv12
    port map (
            O => \N__35796\,
            I => \c0.n18223\
        );

    \I__7664\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35789\
        );

    \I__7663\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35786\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35783\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__35786\,
            I => data_out_2_2
        );

    \I__7660\ : Odrv4
    port map (
            O => \N__35783\,
            I => data_out_2_2
        );

    \I__7659\ : IoInMux
    port map (
            O => \N__35778\,
            I => \N__35775\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__7657\ : Span4Mux_s3_v
    port map (
            O => \N__35772\,
            I => \N__35769\
        );

    \I__7656\ : Sp12to4
    port map (
            O => \N__35769\,
            I => \N__35766\
        );

    \I__7655\ : Span12Mux_h
    port map (
            O => \N__35766\,
            I => \N__35763\
        );

    \I__7654\ : Odrv12
    port map (
            O => \N__35763\,
            I => \PIN_24_c_3\
        );

    \I__7653\ : CEMux
    port map (
            O => \N__35760\,
            I => \N__35757\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35754\
        );

    \I__7651\ : Span4Mux_v
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__35751\,
            I => \control.n6\
        );

    \I__7649\ : SRMux
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__35745\,
            I => \control.n17251\
        );

    \I__7647\ : IoInMux
    port map (
            O => \N__35742\,
            I => \N__35739\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__35739\,
            I => \N__35736\
        );

    \I__7645\ : Span12Mux_s10_v
    port map (
            O => \N__35736\,
            I => \N__35733\
        );

    \I__7644\ : Span12Mux_h
    port map (
            O => \N__35733\,
            I => \N__35730\
        );

    \I__7643\ : Odrv12
    port map (
            O => \N__35730\,
            I => \PIN_23_c_4\
        );

    \I__7642\ : CEMux
    port map (
            O => \N__35727\,
            I => \N__35724\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__35724\,
            I => \N__35720\
        );

    \I__7640\ : CEMux
    port map (
            O => \N__35723\,
            I => \N__35717\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__35720\,
            I => \N__35714\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35711\
        );

    \I__7637\ : Span4Mux_h
    port map (
            O => \N__35714\,
            I => \N__35708\
        );

    \I__7636\ : Span4Mux_v
    port map (
            O => \N__35711\,
            I => \N__35705\
        );

    \I__7635\ : Odrv4
    port map (
            O => \N__35708\,
            I => \control.n6_adj_2460\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__35705\,
            I => \control.n6_adj_2460\
        );

    \I__7633\ : SRMux
    port map (
            O => \N__35700\,
            I => \N__35697\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__35697\,
            I => \N__35694\
        );

    \I__7631\ : Odrv12
    port map (
            O => \N__35694\,
            I => \control.n10490\
        );

    \I__7630\ : InMux
    port map (
            O => \N__35691\,
            I => \N__35686\
        );

    \I__7629\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35683\
        );

    \I__7628\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35680\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35676\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35672\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35669\
        );

    \I__7624\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35666\
        );

    \I__7623\ : Span4Mux_h
    port map (
            O => \N__35676\,
            I => \N__35660\
        );

    \I__7622\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35657\
        );

    \I__7621\ : Span4Mux_v
    port map (
            O => \N__35672\,
            I => \N__35649\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__35669\,
            I => \N__35649\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N__35649\
        );

    \I__7618\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35646\
        );

    \I__7617\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35643\
        );

    \I__7616\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35640\
        );

    \I__7615\ : Span4Mux_h
    port map (
            O => \N__35660\,
            I => \N__35633\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35633\
        );

    \I__7613\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35630\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__35649\,
            I => \N__35625\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35625\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__35643\,
            I => \N__35620\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__35640\,
            I => \N__35620\
        );

    \I__7608\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35617\
        );

    \I__7607\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35614\
        );

    \I__7606\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35611\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35608\
        );

    \I__7604\ : Span4Mux_h
    port map (
            O => \N__35625\,
            I => \N__35603\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__35620\,
            I => \N__35603\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__35617\,
            I => \N__35600\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__35614\,
            I => \N__35593\
        );

    \I__7600\ : Sp12to4
    port map (
            O => \N__35611\,
            I => \N__35593\
        );

    \I__7599\ : Sp12to4
    port map (
            O => \N__35608\,
            I => \N__35593\
        );

    \I__7598\ : Span4Mux_h
    port map (
            O => \N__35603\,
            I => \N__35588\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__35600\,
            I => \N__35588\
        );

    \I__7596\ : Span12Mux_s9_v
    port map (
            O => \N__35593\,
            I => \N__35585\
        );

    \I__7595\ : Span4Mux_v
    port map (
            O => \N__35588\,
            I => \N__35582\
        );

    \I__7594\ : Odrv12
    port map (
            O => \N__35585\,
            I => hall3
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__35582\,
            I => hall3
        );

    \I__7592\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35571\
        );

    \I__7591\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35568\
        );

    \I__7590\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35563\
        );

    \I__7589\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35560\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__35571\,
            I => \N__35556\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35553\
        );

    \I__7586\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35550\
        );

    \I__7585\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35547\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35542\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__35560\,
            I => \N__35539\
        );

    \I__7582\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35536\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__35556\,
            I => \N__35527\
        );

    \I__7580\ : Span4Mux_v
    port map (
            O => \N__35553\,
            I => \N__35527\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__35550\,
            I => \N__35527\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35527\
        );

    \I__7577\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35524\
        );

    \I__7576\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35521\
        );

    \I__7575\ : Span4Mux_v
    port map (
            O => \N__35542\,
            I => \N__35516\
        );

    \I__7574\ : Span4Mux_v
    port map (
            O => \N__35539\,
            I => \N__35516\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__35536\,
            I => \N__35513\
        );

    \I__7572\ : Span4Mux_h
    port map (
            O => \N__35527\,
            I => \N__35508\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35505\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35502\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__35516\,
            I => \N__35497\
        );

    \I__7568\ : Span4Mux_v
    port map (
            O => \N__35513\,
            I => \N__35497\
        );

    \I__7567\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35494\
        );

    \I__7566\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35491\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__35508\,
            I => \N__35486\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__35505\,
            I => \N__35486\
        );

    \I__7563\ : Span12Mux_h
    port map (
            O => \N__35502\,
            I => \N__35477\
        );

    \I__7562\ : Sp12to4
    port map (
            O => \N__35497\,
            I => \N__35477\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__35494\,
            I => \N__35477\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35477\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__35486\,
            I => hall2
        );

    \I__7558\ : Odrv12
    port map (
            O => \N__35477\,
            I => hall2
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__35472\,
            I => \N__35467\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__35471\,
            I => \N__35464\
        );

    \I__7555\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35458\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35455\
        );

    \I__7553\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35451\
        );

    \I__7552\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35448\
        );

    \I__7551\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35445\
        );

    \I__7550\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35438\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35433\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__35455\,
            I => \N__35433\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__35454\,
            I => \N__35430\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__35451\,
            I => \N__35423\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__35448\,
            I => \N__35423\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__35445\,
            I => \N__35423\
        );

    \I__7543\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35420\
        );

    \I__7542\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35415\
        );

    \I__7541\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35415\
        );

    \I__7540\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35412\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__35438\,
            I => \N__35408\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__35433\,
            I => \N__35405\
        );

    \I__7537\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35402\
        );

    \I__7536\ : Span4Mux_v
    port map (
            O => \N__35423\,
            I => \N__35399\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__35420\,
            I => \N__35392\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__35415\,
            I => \N__35392\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__35412\,
            I => \N__35392\
        );

    \I__7532\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35389\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__35408\,
            I => \N__35386\
        );

    \I__7530\ : Span4Mux_h
    port map (
            O => \N__35405\,
            I => \N__35383\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__35402\,
            I => \N__35380\
        );

    \I__7528\ : Span4Mux_h
    port map (
            O => \N__35399\,
            I => \N__35375\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__35392\,
            I => \N__35375\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__35389\,
            I => \N__35372\
        );

    \I__7525\ : Sp12to4
    port map (
            O => \N__35386\,
            I => \N__35369\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__35383\,
            I => \N__35364\
        );

    \I__7523\ : Span4Mux_v
    port map (
            O => \N__35380\,
            I => \N__35364\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__35375\,
            I => \N__35359\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__35372\,
            I => \N__35359\
        );

    \I__7520\ : Odrv12
    port map (
            O => \N__35369\,
            I => hall1
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__35364\,
            I => hall1
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__35359\,
            I => hall1
        );

    \I__7517\ : SRMux
    port map (
            O => \N__35352\,
            I => \N__35348\
        );

    \I__7516\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35344\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__35348\,
            I => \N__35341\
        );

    \I__7514\ : SRMux
    port map (
            O => \N__35347\,
            I => \N__35338\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35334\
        );

    \I__7512\ : Span4Mux_v
    port map (
            O => \N__35341\,
            I => \N__35329\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__35338\,
            I => \N__35329\
        );

    \I__7510\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35326\
        );

    \I__7509\ : Span4Mux_v
    port map (
            O => \N__35334\,
            I => \N__35321\
        );

    \I__7508\ : Span4Mux_h
    port map (
            O => \N__35329\,
            I => \N__35316\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35316\
        );

    \I__7506\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35312\
        );

    \I__7505\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35309\
        );

    \I__7504\ : Span4Mux_h
    port map (
            O => \N__35321\,
            I => \N__35304\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__35316\,
            I => \N__35304\
        );

    \I__7502\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35301\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__35312\,
            I => \control.PHASES_5__N_2160\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__35309\,
            I => \control.PHASES_5__N_2160\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__35304\,
            I => \control.PHASES_5__N_2160\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__35301\,
            I => \control.PHASES_5__N_2160\
        );

    \I__7497\ : IoInMux
    port map (
            O => \N__35292\,
            I => \N__35289\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__35289\,
            I => \N__35286\
        );

    \I__7495\ : Span12Mux_s3_v
    port map (
            O => \N__35286\,
            I => \N__35283\
        );

    \I__7494\ : Span12Mux_h
    port map (
            O => \N__35283\,
            I => \N__35280\
        );

    \I__7493\ : Odrv12
    port map (
            O => \N__35280\,
            I => \control.PHASES_5_N_2130_5\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__35277\,
            I => \N__35274\
        );

    \I__7491\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35271\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35268\
        );

    \I__7489\ : Span12Mux_h
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__7488\ : Odrv12
    port map (
            O => \N__35265\,
            I => \c0.n17748\
        );

    \I__7487\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35259\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35256\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__35256\,
            I => \c0.n18191\
        );

    \I__7484\ : CascadeMux
    port map (
            O => \N__35253\,
            I => \c0.n18867_cascade_\
        );

    \I__7483\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35240\
        );

    \I__7482\ : InMux
    port map (
            O => \N__35249\,
            I => \N__35240\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__35248\,
            I => \N__35237\
        );

    \I__7480\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35227\
        );

    \I__7479\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35224\
        );

    \I__7478\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35221\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35213\
        );

    \I__7476\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35208\
        );

    \I__7475\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35208\
        );

    \I__7474\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35203\
        );

    \I__7473\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35203\
        );

    \I__7472\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35196\
        );

    \I__7471\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35196\
        );

    \I__7470\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35196\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35187\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35180\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__35224\,
            I => \N__35180\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__35221\,
            I => \N__35180\
        );

    \I__7465\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35177\
        );

    \I__7464\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35168\
        );

    \I__7463\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35168\
        );

    \I__7462\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35168\
        );

    \I__7461\ : InMux
    port map (
            O => \N__35216\,
            I => \N__35168\
        );

    \I__7460\ : Span4Mux_h
    port map (
            O => \N__35213\,
            I => \N__35165\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__35208\,
            I => \N__35162\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35157\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__35196\,
            I => \N__35157\
        );

    \I__7456\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35154\
        );

    \I__7455\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35145\
        );

    \I__7454\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35145\
        );

    \I__7453\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35145\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35145\
        );

    \I__7451\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35141\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__35187\,
            I => \N__35134\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__35180\,
            I => \N__35134\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35134\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35127\
        );

    \I__7446\ : Span4Mux_v
    port map (
            O => \N__35165\,
            I => \N__35127\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__35162\,
            I => \N__35127\
        );

    \I__7444\ : Span12Mux_h
    port map (
            O => \N__35157\,
            I => \N__35120\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__35154\,
            I => \N__35120\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__35145\,
            I => \N__35120\
        );

    \I__7441\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35117\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__35141\,
            I => byte_transmit_counter_2
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__35134\,
            I => byte_transmit_counter_2
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__35127\,
            I => byte_transmit_counter_2
        );

    \I__7437\ : Odrv12
    port map (
            O => \N__35120\,
            I => byte_transmit_counter_2
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__35117\,
            I => byte_transmit_counter_2
        );

    \I__7435\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__35100\,
            I => n10_adj_2505
        );

    \I__7432\ : CascadeMux
    port map (
            O => \N__35097\,
            I => \n18870_cascade_\
        );

    \I__7431\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35089\
        );

    \I__7430\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35085\
        );

    \I__7429\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35082\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__35089\,
            I => \N__35077\
        );

    \I__7427\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35074\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__35085\,
            I => \N__35066\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35066\
        );

    \I__7424\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35063\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35060\
        );

    \I__7422\ : Span4Mux_h
    port map (
            O => \N__35077\,
            I => \N__35055\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__35074\,
            I => \N__35055\
        );

    \I__7420\ : InMux
    port map (
            O => \N__35073\,
            I => \N__35050\
        );

    \I__7419\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35050\
        );

    \I__7418\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35046\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__35066\,
            I => \N__35041\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35041\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__35060\,
            I => \N__35038\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__35055\,
            I => \N__35033\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35033\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35049\,
            I => \N__35030\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35046\,
            I => byte_transmit_counter_3
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__35041\,
            I => byte_transmit_counter_3
        );

    \I__7409\ : Odrv12
    port map (
            O => \N__35038\,
            I => byte_transmit_counter_3
        );

    \I__7408\ : Odrv4
    port map (
            O => \N__35033\,
            I => byte_transmit_counter_3
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__35030\,
            I => byte_transmit_counter_3
        );

    \I__7406\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35016\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__35016\,
            I => n10_adj_2530
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__35013\,
            I => \N__35010\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35007\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__35007\,
            I => \c0.n5_adj_2214\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35004\,
            I => \N__35000\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34997\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35000\,
            I => \N__34994\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__34997\,
            I => \c0.data_out_1_4\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__34994\,
            I => \c0.data_out_1_4\
        );

    \I__7396\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__34986\,
            I => \c0.n18190\
        );

    \I__7394\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34977\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__34977\,
            I => \c0.n2_adj_2348\
        );

    \I__7391\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34971\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__34971\,
            I => \c0.n18334\
        );

    \I__7389\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__34965\,
            I => \c0.n17819\
        );

    \I__7387\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34959\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__34959\,
            I => \c0.n6_adj_2277\
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__34956\,
            I => \N__34952\
        );

    \I__7384\ : CascadeMux
    port map (
            O => \N__34955\,
            I => \N__34949\
        );

    \I__7383\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34945\
        );

    \I__7382\ : InMux
    port map (
            O => \N__34949\,
            I => \N__34942\
        );

    \I__7381\ : InMux
    port map (
            O => \N__34948\,
            I => \N__34939\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__34945\,
            I => \c0.data_out_9_4\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__34942\,
            I => \c0.data_out_9_4\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__34939\,
            I => \c0.data_out_9_4\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__34932\,
            I => \c0.n8_adj_2211_cascade_\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__34929\,
            I => \c0.n18222_cascade_\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__34926\,
            I => \c0.n18693_cascade_\
        );

    \I__7374\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__34917\,
            I => n18696
        );

    \I__7371\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34905\
        );

    \I__7370\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34905\
        );

    \I__7369\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34900\
        );

    \I__7368\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34900\
        );

    \I__7367\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34897\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__34905\,
            I => \N__34890\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__34900\,
            I => \N__34890\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__34897\,
            I => \N__34890\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__34890\,
            I => \N__34887\
        );

    \I__7362\ : Odrv4
    port map (
            O => \N__34887\,
            I => \c0.data_out_6_2\
        );

    \I__7361\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34881\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__34881\,
            I => \c0.n5_adj_2347\
        );

    \I__7359\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34873\
        );

    \I__7358\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34862\
        );

    \I__7357\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34862\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__34873\,
            I => \N__34859\
        );

    \I__7355\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34853\
        );

    \I__7354\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34848\
        );

    \I__7353\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34845\
        );

    \I__7352\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34839\
        );

    \I__7351\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34839\
        );

    \I__7350\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34836\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34829\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__34859\,
            I => \N__34826\
        );

    \I__7347\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34823\
        );

    \I__7346\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34820\
        );

    \I__7345\ : CascadeMux
    port map (
            O => \N__34856\,
            I => \N__34817\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34814\
        );

    \I__7343\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34811\
        );

    \I__7342\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34808\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34805\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34802\
        );

    \I__7339\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34799\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34796\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N__34793\
        );

    \I__7336\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34784\
        );

    \I__7335\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34784\
        );

    \I__7334\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34784\
        );

    \I__7333\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34784\
        );

    \I__7332\ : Sp12to4
    port map (
            O => \N__34829\,
            I => \N__34775\
        );

    \I__7331\ : Sp12to4
    port map (
            O => \N__34826\,
            I => \N__34775\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__34823\,
            I => \N__34775\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34775\
        );

    \I__7328\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34771\
        );

    \I__7327\ : Span12Mux_v
    port map (
            O => \N__34814\,
            I => \N__34768\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__34811\,
            I => \N__34763\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__34808\,
            I => \N__34763\
        );

    \I__7324\ : Span4Mux_v
    port map (
            O => \N__34805\,
            I => \N__34760\
        );

    \I__7323\ : Span4Mux_v
    port map (
            O => \N__34802\,
            I => \N__34753\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__34799\,
            I => \N__34753\
        );

    \I__7321\ : Span4Mux_h
    port map (
            O => \N__34796\,
            I => \N__34753\
        );

    \I__7320\ : Span12Mux_v
    port map (
            O => \N__34793\,
            I => \N__34746\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__34784\,
            I => \N__34746\
        );

    \I__7318\ : Span12Mux_h
    port map (
            O => \N__34775\,
            I => \N__34746\
        );

    \I__7317\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34743\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__34771\,
            I => byte_transmit_counter_1
        );

    \I__7315\ : Odrv12
    port map (
            O => \N__34768\,
            I => byte_transmit_counter_1
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__34763\,
            I => byte_transmit_counter_1
        );

    \I__7313\ : Odrv4
    port map (
            O => \N__34760\,
            I => byte_transmit_counter_1
        );

    \I__7312\ : Odrv4
    port map (
            O => \N__34753\,
            I => byte_transmit_counter_1
        );

    \I__7311\ : Odrv12
    port map (
            O => \N__34746\,
            I => byte_transmit_counter_1
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__34743\,
            I => byte_transmit_counter_1
        );

    \I__7309\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34725\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__34725\,
            I => \N__34720\
        );

    \I__7307\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34715\
        );

    \I__7306\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34715\
        );

    \I__7305\ : Odrv4
    port map (
            O => \N__34720\,
            I => \c0.data_out_9_7\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__34715\,
            I => \c0.data_out_9_7\
        );

    \I__7303\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34707\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__34707\,
            I => \c0.n17774\
        );

    \I__7301\ : CascadeMux
    port map (
            O => \N__34704\,
            I => \c0.n17774_cascade_\
        );

    \I__7300\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34691\
        );

    \I__7299\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34691\
        );

    \I__7298\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34691\
        );

    \I__7297\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34688\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__34691\,
            I => \c0.data_out_10_3\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__34688\,
            I => \c0.data_out_10_3\
        );

    \I__7294\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34680\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34674\
        );

    \I__7292\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34669\
        );

    \I__7291\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34669\
        );

    \I__7290\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34666\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__34674\,
            I => \N__34661\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34661\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__34666\,
            I => \c0.data_out_10_5\
        );

    \I__7286\ : Odrv4
    port map (
            O => \N__34661\,
            I => \c0.data_out_10_5\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__34653\,
            I => \N__34650\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__34650\,
            I => \c0.n6_adj_2314\
        );

    \I__7282\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34641\
        );

    \I__7281\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34641\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34638\
        );

    \I__7279\ : Odrv12
    port map (
            O => \N__34638\,
            I => \c0.n17883\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__34635\,
            I => \c0.n10801_cascade_\
        );

    \I__7277\ : InMux
    port map (
            O => \N__34632\,
            I => \N__34627\
        );

    \I__7276\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34624\
        );

    \I__7275\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34621\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__34627\,
            I => \N__34618\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__34624\,
            I => \N__34613\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__34621\,
            I => \N__34613\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__34618\,
            I => \c0.data_out_10_0\
        );

    \I__7270\ : Odrv12
    port map (
            O => \N__34613\,
            I => \c0.data_out_10_0\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34604\
        );

    \I__7268\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34601\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__34604\,
            I => \c0.n17768\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__34601\,
            I => \c0.n17768\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__34596\,
            I => \c0.n10_adj_2366_cascade_\
        );

    \I__7264\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34585\
        );

    \I__7263\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34585\
        );

    \I__7262\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34582\
        );

    \I__7261\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34579\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34576\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__34582\,
            I => \c0.data_out_10_1\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__34579\,
            I => \c0.data_out_10_1\
        );

    \I__7257\ : Odrv4
    port map (
            O => \N__34576\,
            I => \c0.data_out_10_1\
        );

    \I__7256\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34566\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__34566\,
            I => \N__34560\
        );

    \I__7254\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34557\
        );

    \I__7253\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34554\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34551\
        );

    \I__7251\ : Span4Mux_v
    port map (
            O => \N__34560\,
            I => \N__34542\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__34557\,
            I => \N__34542\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__34554\,
            I => \N__34542\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34542\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__34542\,
            I => \N__34539\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__34539\,
            I => \c0.data_out_6_1\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__34536\,
            I => \c0.n6_adj_2318_cascade_\
        );

    \I__7244\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34529\
        );

    \I__7243\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34526\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__34529\,
            I => \N__34520\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__34526\,
            I => \N__34520\
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__34525\,
            I => \N__34516\
        );

    \I__7239\ : Span4Mux_v
    port map (
            O => \N__34520\,
            I => \N__34513\
        );

    \I__7238\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34510\
        );

    \I__7237\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34507\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__34513\,
            I => \N__34504\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__34510\,
            I => \N__34499\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__34507\,
            I => \N__34499\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__34504\,
            I => \c0.data_out_9_0\
        );

    \I__7232\ : Odrv12
    port map (
            O => \N__34499\,
            I => \c0.data_out_9_0\
        );

    \I__7231\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34489\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__34493\,
            I => \N__34486\
        );

    \I__7229\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34482\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__34489\,
            I => \N__34479\
        );

    \I__7227\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34476\
        );

    \I__7226\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34473\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34470\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__34479\,
            I => \N__34467\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__34476\,
            I => \c0.data_out_9_6\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__34473\,
            I => \c0.data_out_9_6\
        );

    \I__7221\ : Odrv12
    port map (
            O => \N__34470\,
            I => \c0.data_out_9_6\
        );

    \I__7220\ : Odrv4
    port map (
            O => \N__34467\,
            I => \c0.data_out_9_6\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34455\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__34455\,
            I => \c0.n6_adj_2367\
        );

    \I__7217\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34449\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34449\,
            I => \c0.n17850\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__7214\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34440\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__34440\,
            I => \N__34436\
        );

    \I__7212\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34433\
        );

    \I__7211\ : Span4Mux_v
    port map (
            O => \N__34436\,
            I => \N__34428\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34428\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__34428\,
            I => \c0.n10749\
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__34425\,
            I => \c0.data_out_9__2__N_367_cascade_\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__34422\,
            I => \c0.n15_adj_2319_cascade_\
        );

    \I__7206\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34416\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__34416\,
            I => \N__34413\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__34413\,
            I => \c0.n14_adj_2320\
        );

    \I__7203\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34405\
        );

    \I__7202\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34400\
        );

    \I__7201\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34400\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__34405\,
            I => \c0.data_out_10_2\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__34400\,
            I => \c0.data_out_10_2\
        );

    \I__7198\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34389\
        );

    \I__7197\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34389\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__34386\,
            I => \c0.n17826\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__34383\,
            I => \c0.n17761_cascade_\
        );

    \I__7193\ : InMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34373\
        );

    \I__7191\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34370\
        );

    \I__7190\ : Odrv4
    port map (
            O => \N__34373\,
            I => n9_adj_2477
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34370\,
            I => n9_adj_2477
        );

    \I__7188\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34362\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__34362\,
            I => \c0.n17761\
        );

    \I__7186\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__34353\,
            I => \c0.n18747\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__34350\,
            I => \c0.n17807_cascade_\
        );

    \I__7182\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34344\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__34344\,
            I => \N__34338\
        );

    \I__7180\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34333\
        );

    \I__7179\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34328\
        );

    \I__7178\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34328\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__34338\,
            I => \N__34325\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34322\
        );

    \I__7175\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34319\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__34333\,
            I => data_out_9_2
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__34328\,
            I => data_out_9_2
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__34325\,
            I => data_out_9_2
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__34322\,
            I => data_out_9_2
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__34319\,
            I => data_out_9_2
        );

    \I__7169\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34305\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__34302\,
            I => \N__34298\
        );

    \I__7166\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34294\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34291\
        );

    \I__7164\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34288\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__34294\,
            I => data_in_3_1
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__34291\,
            I => data_in_3_1
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__34288\,
            I => data_in_3_1
        );

    \I__7160\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34277\
        );

    \I__7159\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34274\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34268\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34268\
        );

    \I__7156\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34265\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__34268\,
            I => \N__34262\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__34265\,
            I => data_in_2_1
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__34262\,
            I => data_in_2_1
        );

    \I__7152\ : InMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__34254\,
            I => \N__34251\
        );

    \I__7150\ : Span4Mux_h
    port map (
            O => \N__34251\,
            I => \N__34247\
        );

    \I__7149\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34243\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__34247\,
            I => \N__34240\
        );

    \I__7147\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__34243\,
            I => data_in_3_3
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__34240\,
            I => data_in_3_3
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__34237\,
            I => data_in_3_3
        );

    \I__7143\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34222\
        );

    \I__7142\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34222\
        );

    \I__7141\ : CascadeMux
    port map (
            O => \N__34228\,
            I => \N__34213\
        );

    \I__7140\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34205\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__34222\,
            I => \N__34202\
        );

    \I__7138\ : CascadeMux
    port map (
            O => \N__34221\,
            I => \N__34199\
        );

    \I__7137\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34189\
        );

    \I__7136\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34172\
        );

    \I__7135\ : InMux
    port map (
            O => \N__34218\,
            I => \N__34172\
        );

    \I__7134\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34172\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34165\
        );

    \I__7132\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34165\
        );

    \I__7131\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34165\
        );

    \I__7130\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34156\
        );

    \I__7129\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34156\
        );

    \I__7128\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34156\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34156\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34153\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__34202\,
            I => \N__34150\
        );

    \I__7124\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34143\
        );

    \I__7123\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34143\
        );

    \I__7122\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34143\
        );

    \I__7121\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34132\
        );

    \I__7120\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34132\
        );

    \I__7119\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34132\
        );

    \I__7118\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34132\
        );

    \I__7117\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34132\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34129\
        );

    \I__7115\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34123\
        );

    \I__7114\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34118\
        );

    \I__7113\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34118\
        );

    \I__7112\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34113\
        );

    \I__7111\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34113\
        );

    \I__7110\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34106\
        );

    \I__7109\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34106\
        );

    \I__7108\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34106\
        );

    \I__7107\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34101\
        );

    \I__7106\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34101\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__34172\,
            I => \N__34098\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__34165\,
            I => \N__34093\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__34156\,
            I => \N__34093\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__34153\,
            I => \N__34090\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__34150\,
            I => \N__34087\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__34143\,
            I => \N__34080\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__34132\,
            I => \N__34080\
        );

    \I__7098\ : Span4Mux_h
    port map (
            O => \N__34129\,
            I => \N__34080\
        );

    \I__7097\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34073\
        );

    \I__7096\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34073\
        );

    \I__7095\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34073\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__34123\,
            I => rx_data_ready
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__34118\,
            I => rx_data_ready
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__34113\,
            I => rx_data_ready
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__34106\,
            I => rx_data_ready
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__34101\,
            I => rx_data_ready
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__34098\,
            I => rx_data_ready
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__34093\,
            I => rx_data_ready
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__34090\,
            I => rx_data_ready
        );

    \I__7086\ : Odrv4
    port map (
            O => \N__34087\,
            I => rx_data_ready
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__34080\,
            I => rx_data_ready
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__34073\,
            I => rx_data_ready
        );

    \I__7083\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34045\
        );

    \I__7082\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34042\
        );

    \I__7081\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34039\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__34045\,
            I => \N__34036\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__34042\,
            I => \N__34033\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__34039\,
            I => \N__34030\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__34036\,
            I => \N__34024\
        );

    \I__7076\ : Span4Mux_h
    port map (
            O => \N__34033\,
            I => \N__34024\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__34030\,
            I => \N__34021\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34018\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__34024\,
            I => \N__34013\
        );

    \I__7072\ : Span4Mux_h
    port map (
            O => \N__34021\,
            I => \N__34013\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34018\,
            I => data_in_2_3
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__34013\,
            I => data_in_2_3
        );

    \I__7069\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__34002\,
            I => \c0.n18365\
        );

    \I__7066\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33996\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33993\
        );

    \I__7064\ : Span4Mux_s1_v
    port map (
            O => \N__33993\,
            I => \N__33990\
        );

    \I__7063\ : Span4Mux_v
    port map (
            O => \N__33990\,
            I => \N__33986\
        );

    \I__7062\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33983\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__33986\,
            I => \N__33980\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__33983\,
            I => data_out_frame2_18_5
        );

    \I__7059\ : Odrv4
    port map (
            O => \N__33980\,
            I => data_out_frame2_18_5
        );

    \I__7058\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33972\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__33972\,
            I => n1
        );

    \I__7056\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33966\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__33963\,
            I => \N__33960\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__33960\,
            I => n24_adj_2523
        );

    \I__7052\ : InMux
    port map (
            O => \N__33957\,
            I => \N__33954\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__33954\,
            I => n18_adj_2526
        );

    \I__7050\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__7048\ : Odrv4
    port map (
            O => \N__33945\,
            I => \c0.n5_adj_2436\
        );

    \I__7047\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33931\
        );

    \I__7046\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33931\
        );

    \I__7045\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33928\
        );

    \I__7044\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33925\
        );

    \I__7043\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33918\
        );

    \I__7042\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33918\
        );

    \I__7041\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33918\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33915\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33911\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33906\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__33918\,
            I => \N__33906\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__33915\,
            I => \N__33903\
        );

    \I__7035\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33900\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__33911\,
            I => \N__33895\
        );

    \I__7033\ : Span4Mux_v
    port map (
            O => \N__33906\,
            I => \N__33895\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__33903\,
            I => \N__33892\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__33900\,
            I => \r_Bit_Index_0_adj_2519\
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__33895\,
            I => \r_Bit_Index_0_adj_2519\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__33892\,
            I => \r_Bit_Index_0_adj_2519\
        );

    \I__7028\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33877\
        );

    \I__7027\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33877\
        );

    \I__7026\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33874\
        );

    \I__7025\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33871\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33866\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33866\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33861\
        );

    \I__7021\ : Span4Mux_v
    port map (
            O => \N__33866\,
            I => \N__33861\
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__33861\,
            I => \r_Bit_Index_1_adj_2518\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__33858\,
            I => \N__33854\
        );

    \I__7018\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33847\
        );

    \I__7017\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33844\
        );

    \I__7016\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33835\
        );

    \I__7015\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33835\
        );

    \I__7014\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33835\
        );

    \I__7013\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33835\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33831\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__33844\,
            I => \N__33826\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33826\
        );

    \I__7009\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33823\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__33831\,
            I => \N__33818\
        );

    \I__7007\ : Span4Mux_h
    port map (
            O => \N__33826\,
            I => \N__33818\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__33823\,
            I => \tx_transmit_N_1947_3\
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__33818\,
            I => \tx_transmit_N_1947_3\
        );

    \I__7004\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__33807\,
            I => \N__33803\
        );

    \I__7001\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33800\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__33803\,
            I => \c0.n85\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__33800\,
            I => \c0.n85\
        );

    \I__6998\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33791\
        );

    \I__6997\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33784\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33781\
        );

    \I__6995\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33772\
        );

    \I__6994\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33772\
        );

    \I__6993\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33772\
        );

    \I__6992\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33772\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__33784\,
            I => \c0.n14068\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__33781\,
            I => \c0.n14068\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__33772\,
            I => \c0.n14068\
        );

    \I__6988\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__33759\,
            I => \N__33756\
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__33756\,
            I => \c0.n18259\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__33753\,
            I => \N__33749\
        );

    \I__6983\ : InMux
    port map (
            O => \N__33752\,
            I => \N__33743\
        );

    \I__6982\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33743\
        );

    \I__6981\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33740\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__33743\,
            I => \N__33737\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__33740\,
            I => \N__33734\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__33737\,
            I => \N__33731\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__33734\,
            I => \N__33728\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__33731\,
            I => n18014
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__33728\,
            I => n18014
        );

    \I__6974\ : CascadeMux
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6973\ : InMux
    port map (
            O => \N__33720\,
            I => \N__33717\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__33717\,
            I => \N__33714\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__33714\,
            I => \N__33711\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__33711\,
            I => n4_adj_2472
        );

    \I__6969\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33701\
        );

    \I__6968\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33701\
        );

    \I__6967\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33698\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__33701\,
            I => \N__33695\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__33698\,
            I => \N__33692\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__33695\,
            I => \N__33689\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__33692\,
            I => \N__33686\
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__33689\,
            I => n11545
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__33686\,
            I => n11545
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__33681\,
            I => \N__33676\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33673\
        );

    \I__6958\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33668\
        );

    \I__6957\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33668\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__33673\,
            I => \N__33664\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33661\
        );

    \I__6954\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33658\
        );

    \I__6953\ : Span4Mux_v
    port map (
            O => \N__33664\,
            I => \N__33655\
        );

    \I__6952\ : Span4Mux_h
    port map (
            O => \N__33661\,
            I => \N__33652\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__33658\,
            I => \r_Bit_Index_2_adj_2517\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__33655\,
            I => \r_Bit_Index_2_adj_2517\
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__33652\,
            I => \r_Bit_Index_2_adj_2517\
        );

    \I__6948\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33641\
        );

    \I__6947\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33638\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__33641\,
            I => \N__33635\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33632\
        );

    \I__6944\ : Span4Mux_s2_v
    port map (
            O => \N__33635\,
            I => \N__33629\
        );

    \I__6943\ : Span12Mux_s8_v
    port map (
            O => \N__33632\,
            I => \N__33626\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__33629\,
            I => \N__33623\
        );

    \I__6941\ : Odrv12
    port map (
            O => \N__33626\,
            I => \c0.n17715\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__33623\,
            I => \c0.n17715\
        );

    \I__6939\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33614\
        );

    \I__6938\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33611\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__33614\,
            I => \N__33608\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__33611\,
            I => \c0.delay_counter_3\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__33608\,
            I => \c0.delay_counter_3\
        );

    \I__6934\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33599\
        );

    \I__6933\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33596\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__33599\,
            I => \c0.delay_counter_8\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__33596\,
            I => \c0.delay_counter_8\
        );

    \I__6930\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__33588\,
            I => \c0.n18\
        );

    \I__6928\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33581\
        );

    \I__6927\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33578\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33581\,
            I => \c0.delay_counter_10\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__33578\,
            I => \c0.delay_counter_10\
        );

    \I__6924\ : CascadeMux
    port map (
            O => \N__33573\,
            I => \N__33570\
        );

    \I__6923\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33566\
        );

    \I__6922\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33563\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__33566\,
            I => \c0.delay_counter_0\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__33563\,
            I => \c0.delay_counter_0\
        );

    \I__6919\ : CascadeMux
    port map (
            O => \N__33558\,
            I => \N__33554\
        );

    \I__6918\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33551\
        );

    \I__6917\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__33551\,
            I => \c0.delay_counter_13\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__33548\,
            I => \c0.delay_counter_13\
        );

    \I__6914\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33539\
        );

    \I__6913\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33536\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__33539\,
            I => \c0.delay_counter_6\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__33536\,
            I => \c0.delay_counter_6\
        );

    \I__6910\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__6908\ : Span4Mux_s2_v
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__33519\,
            I => \c0.n18810\
        );

    \I__6905\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33511\
        );

    \I__6904\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33508\
        );

    \I__6903\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33505\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__33511\,
            I => \N__33502\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__33508\,
            I => \N__33497\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33497\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__33502\,
            I => \c0.tx_transmit_N_1947_0\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__33497\,
            I => \c0.tx_transmit_N_1947_0\
        );

    \I__6897\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33487\
        );

    \I__6896\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33484\
        );

    \I__6895\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33481\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__33487\,
            I => \N__33478\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__33484\,
            I => \c0.tx_transmit_N_1947_1\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__33481\,
            I => \c0.tx_transmit_N_1947_1\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__33478\,
            I => \c0.tx_transmit_N_1947_1\
        );

    \I__6890\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33466\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33463\
        );

    \I__6888\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33460\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33457\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__33463\,
            I => \c0.tx_transmit_N_1947_2\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__33460\,
            I => \c0.tx_transmit_N_1947_2\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__33457\,
            I => \c0.tx_transmit_N_1947_2\
        );

    \I__6883\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33447\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33442\
        );

    \I__6881\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33437\
        );

    \I__6880\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33437\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__33442\,
            I => \c0.n155\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__33437\,
            I => \c0.n155\
        );

    \I__6877\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33428\
        );

    \I__6876\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33425\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__33428\,
            I => \c0.delay_counter_9\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__33425\,
            I => \c0.delay_counter_9\
        );

    \I__6873\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33416\
        );

    \I__6872\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33413\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__33416\,
            I => \c0.delay_counter_1\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__33413\,
            I => \c0.delay_counter_1\
        );

    \I__6869\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__33405\,
            I => \c0.n22\
        );

    \I__6867\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__33393\,
            I => n25_adj_2468
        );

    \I__6863\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__33387\,
            I => \c0.n18807\
        );

    \I__6861\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33379\
        );

    \I__6860\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33376\
        );

    \I__6859\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33373\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__33379\,
            I => \N__33369\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__33376\,
            I => \N__33366\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33363\
        );

    \I__6855\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33360\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__33369\,
            I => \N__33357\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__33366\,
            I => \N__33354\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__33363\,
            I => data_out_frame2_6_7
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__33360\,
            I => data_out_frame2_6_7
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__33357\,
            I => data_out_frame2_6_7
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__33354\,
            I => data_out_frame2_6_7
        );

    \I__6848\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33341\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33338\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__33341\,
            I => data_out_frame2_18_0
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__33338\,
            I => data_out_frame2_18_0
        );

    \I__6844\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33329\
        );

    \I__6843\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33325\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__33329\,
            I => \N__33321\
        );

    \I__6841\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33317\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33314\
        );

    \I__6839\ : InMux
    port map (
            O => \N__33324\,
            I => \N__33311\
        );

    \I__6838\ : Span4Mux_s2_v
    port map (
            O => \N__33321\,
            I => \N__33308\
        );

    \I__6837\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33305\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__33317\,
            I => data_out_frame2_12_1
        );

    \I__6835\ : Odrv4
    port map (
            O => \N__33314\,
            I => data_out_frame2_12_1
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__33311\,
            I => data_out_frame2_12_1
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__33308\,
            I => data_out_frame2_12_1
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__33305\,
            I => data_out_frame2_12_1
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__33294\,
            I => \c0.n10829_cascade_\
        );

    \I__6830\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33284\
        );

    \I__6829\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33284\
        );

    \I__6828\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33278\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33274\
        );

    \I__6826\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33271\
        );

    \I__6825\ : CascadeMux
    port map (
            O => \N__33282\,
            I => \N__33268\
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__33281\,
            I => \N__33265\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33260\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__33277\,
            I => \N__33256\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__33274\,
            I => \N__33250\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__33271\,
            I => \N__33250\
        );

    \I__6819\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33241\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33241\
        );

    \I__6817\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33241\
        );

    \I__6816\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33241\
        );

    \I__6815\ : Span4Mux_v
    port map (
            O => \N__33260\,
            I => \N__33238\
        );

    \I__6814\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33230\
        );

    \I__6813\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33230\
        );

    \I__6812\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33230\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__33250\,
            I => \N__33225\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33225\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__33238\,
            I => \N__33222\
        );

    \I__6808\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33219\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__33230\,
            I => \N__33216\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__33225\,
            I => \N__33213\
        );

    \I__6805\ : Sp12to4
    port map (
            O => \N__33222\,
            I => \N__33210\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33207\
        );

    \I__6803\ : Span4Mux_h
    port map (
            O => \N__33216\,
            I => \N__33204\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__33213\,
            I => \N__33201\
        );

    \I__6801\ : Odrv12
    port map (
            O => \N__33210\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__33207\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__33204\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__33201\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6797\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__33186\,
            I => \c0.n14161\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__33183\,
            I => \N__33171\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33160\
        );

    \I__6792\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33160\
        );

    \I__6791\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33160\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33160\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33157\
        );

    \I__6788\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33154\
        );

    \I__6787\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33151\
        );

    \I__6786\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33146\
        );

    \I__6785\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33146\
        );

    \I__6784\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33143\
        );

    \I__6783\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33137\
        );

    \I__6782\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33137\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33134\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__33157\,
            I => \N__33131\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__33154\,
            I => \N__33124\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__33151\,
            I => \N__33124\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__33146\,
            I => \N__33124\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33121\
        );

    \I__6775\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33118\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__33137\,
            I => \N__33113\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__33134\,
            I => \N__33113\
        );

    \I__6772\ : Span4Mux_v
    port map (
            O => \N__33131\,
            I => \N__33108\
        );

    \I__6771\ : Span4Mux_v
    port map (
            O => \N__33124\,
            I => \N__33108\
        );

    \I__6770\ : Span12Mux_h
    port map (
            O => \N__33121\,
            I => \N__33103\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33103\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__33113\,
            I => \N__33100\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__33108\,
            I => \N__33097\
        );

    \I__6766\ : Odrv12
    port map (
            O => \N__33103\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__33100\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__33097\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33084\
        );

    \I__6762\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33076\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33076\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33076\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33073\
        );

    \I__6758\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33070\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__33073\,
            I => \N__33062\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33062\
        );

    \I__6754\ : Span4Mux_s3_v
    port map (
            O => \N__33067\,
            I => \N__33052\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__33062\,
            I => \N__33052\
        );

    \I__6752\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33041\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33041\
        );

    \I__6750\ : InMux
    port map (
            O => \N__33059\,
            I => \N__33041\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33041\
        );

    \I__6748\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33041\
        );

    \I__6747\ : Span4Mux_h
    port map (
            O => \N__33052\,
            I => \N__33038\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__33041\,
            I => \c0.n50\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__33038\,
            I => \c0.n50\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__33033\,
            I => \n11114_cascade_\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33027\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33027\,
            I => \c0.n17874\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__33021\,
            I => \c0.n17908\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33015\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__6737\ : Odrv12
    port map (
            O => \N__33012\,
            I => \c0.n18_adj_2423\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__33009\,
            I => \c0.n17908_cascade_\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__33003\,
            I => \c0.n28_adj_2425\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__33000\,
            I => \c0.n30_adj_2424_cascade_\
        );

    \I__6732\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__32994\,
            I => \c0.n29_adj_2427\
        );

    \I__6730\ : InMux
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__6728\ : Span4Mux_s2_v
    port map (
            O => \N__32985\,
            I => \N__32981\
        );

    \I__6727\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32978\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__32981\,
            I => \N__32975\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__32978\,
            I => data_out_frame2_17_5
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__32975\,
            I => data_out_frame2_17_5
        );

    \I__6723\ : CascadeMux
    port map (
            O => \N__32970\,
            I => \c0.n18639_cascade_\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \c0.n10700_cascade_\
        );

    \I__6721\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__32961\,
            I => \c0.n21\
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__32958\,
            I => \N__32955\
        );

    \I__6718\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__32952\,
            I => \c0.n17804\
        );

    \I__6716\ : CascadeMux
    port map (
            O => \N__32949\,
            I => \n11017_cascade_\
        );

    \I__6715\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32942\
        );

    \I__6714\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32939\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__32942\,
            I => data_out_0_0
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__32939\,
            I => data_out_0_0
        );

    \I__6711\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32928\
        );

    \I__6710\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32928\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__32928\,
            I => data_out_3_4
        );

    \I__6708\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32918\
        );

    \I__6706\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32915\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__32918\,
            I => \N__32910\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__32915\,
            I => \N__32910\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__32910\,
            I => \control.PHASES_5_N_2152_1\
        );

    \I__6702\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32901\
        );

    \I__6701\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32897\
        );

    \I__6700\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32894\
        );

    \I__6699\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32891\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32888\
        );

    \I__6697\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32885\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__32897\,
            I => \N__32882\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__32894\,
            I => \N__32877\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__32891\,
            I => \N__32877\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__32888\,
            I => \N__32874\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__32885\,
            I => \N__32867\
        );

    \I__6691\ : Span4Mux_v
    port map (
            O => \N__32882\,
            I => \N__32867\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__32877\,
            I => \N__32867\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__32874\,
            I => \control.pwm_delay_9\
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__32867\,
            I => \control.pwm_delay_9\
        );

    \I__6687\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__32859\,
            I => \N__32853\
        );

    \I__6685\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32850\
        );

    \I__6684\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32847\
        );

    \I__6683\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32844\
        );

    \I__6682\ : Sp12to4
    port map (
            O => \N__32853\,
            I => \N__32839\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__32850\,
            I => \N__32839\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__32847\,
            I => \N__32834\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32834\
        );

    \I__6678\ : Span12Mux_s10_v
    port map (
            O => \N__32839\,
            I => \N__32831\
        );

    \I__6677\ : Span12Mux_s10_v
    port map (
            O => \N__32834\,
            I => \N__32828\
        );

    \I__6676\ : Odrv12
    port map (
            O => \N__32831\,
            I => \control.n18\
        );

    \I__6675\ : Odrv12
    port map (
            O => \N__32828\,
            I => \control.n18\
        );

    \I__6674\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32820\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__32820\,
            I => \control.n17926\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__32817\,
            I => \control.PHASES_5__N_2160_cascade_\
        );

    \I__6671\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32810\
        );

    \I__6670\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32807\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__32810\,
            I => \control.n5\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__32807\,
            I => \control.n5\
        );

    \I__6667\ : CascadeMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__6666\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32796\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__32796\,
            I => \control.n17950\
        );

    \I__6664\ : CEMux
    port map (
            O => \N__32793\,
            I => \N__32790\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__6662\ : Span4Mux_s3_v
    port map (
            O => \N__32787\,
            I => \N__32784\
        );

    \I__6661\ : Span4Mux_h
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__32781\,
            I => \N__32778\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__32778\,
            I => \N__32775\
        );

    \I__6658\ : Odrv4
    port map (
            O => \N__32775\,
            I => \control.n9\
        );

    \I__6657\ : CascadeMux
    port map (
            O => \N__32772\,
            I => \c0.n1_cascade_\
        );

    \I__6656\ : CascadeMux
    port map (
            O => \N__32769\,
            I => \N__32766\
        );

    \I__6655\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32763\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32760\
        );

    \I__6653\ : Odrv12
    port map (
            O => \N__32760\,
            I => n22
        );

    \I__6652\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32754\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__32754\,
            I => \c0.n18849\
        );

    \I__6650\ : CascadeMux
    port map (
            O => \N__32751\,
            I => \n18852_cascade_\
        );

    \I__6649\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32745\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__32745\,
            I => n10
        );

    \I__6647\ : CascadeMux
    port map (
            O => \N__32742\,
            I => \N__32739\
        );

    \I__6646\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32736\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__32736\,
            I => \c0.n18264\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__32733\,
            I => \N__32730\
        );

    \I__6643\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32727\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__32727\,
            I => \c0.n8\
        );

    \I__6641\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32721\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__32721\,
            I => n10_adj_2527
        );

    \I__6639\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__32715\,
            I => \c0.n18322\
        );

    \I__6637\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32708\
        );

    \I__6636\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32705\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32702\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__32705\,
            I => data_out_0_1
        );

    \I__6633\ : Odrv12
    port map (
            O => \N__32702\,
            I => data_out_0_1
        );

    \I__6632\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32694\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__32694\,
            I => \c0.n17742\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__32691\,
            I => \N__32688\
        );

    \I__6629\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32685\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__32685\,
            I => \c0.n10558\
        );

    \I__6627\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32678\
        );

    \I__6626\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32675\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__32678\,
            I => \N__32671\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__32675\,
            I => \N__32668\
        );

    \I__6623\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32665\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__32671\,
            I => \c0.data_out_9_5\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__32668\,
            I => \c0.data_out_9_5\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__32665\,
            I => \c0.data_out_9_5\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__32658\,
            I => \c0.n6_adj_2365_cascade_\
        );

    \I__6618\ : CascadeMux
    port map (
            O => \N__32655\,
            I => \N__32652\
        );

    \I__6617\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32649\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__32649\,
            I => \c0.n5_adj_2220\
        );

    \I__6615\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32642\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__32645\,
            I => \N__32639\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__32642\,
            I => \N__32636\
        );

    \I__6612\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32633\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__32636\,
            I => \N__32630\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__32633\,
            I => \r_Tx_Data_4\
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__32630\,
            I => \r_Tx_Data_4\
        );

    \I__6608\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__32622\,
            I => \c0.n18265\
        );

    \I__6606\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \N__32615\
        );

    \I__6605\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32608\
        );

    \I__6604\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32608\
        );

    \I__6603\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32605\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__32613\,
            I => \N__32602\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32595\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__32605\,
            I => \N__32595\
        );

    \I__6599\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32592\
        );

    \I__6598\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32589\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__32600\,
            I => \N__32586\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__32595\,
            I => \N__32580\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32580\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32577\
        );

    \I__6593\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32574\
        );

    \I__6592\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32571\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32567\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__32577\,
            I => \N__32564\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__32574\,
            I => \N__32561\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__32571\,
            I => \N__32558\
        );

    \I__6587\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32555\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__32567\,
            I => \N__32552\
        );

    \I__6585\ : Span4Mux_h
    port map (
            O => \N__32564\,
            I => \N__32549\
        );

    \I__6584\ : Span4Mux_h
    port map (
            O => \N__32561\,
            I => \N__32542\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__32558\,
            I => \N__32542\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32542\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__32552\,
            I => n9667
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__32549\,
            I => n9667
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__32542\,
            I => n9667
        );

    \I__6578\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32526\
        );

    \I__6576\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32520\
        );

    \I__6575\ : InMux
    port map (
            O => \N__32530\,
            I => \N__32517\
        );

    \I__6574\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32514\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32510\
        );

    \I__6572\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32507\
        );

    \I__6571\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32503\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32500\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32493\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__32517\,
            I => \N__32493\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__32514\,
            I => \N__32493\
        );

    \I__6566\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32490\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__32510\,
            I => \N__32485\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32485\
        );

    \I__6563\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32481\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__32503\,
            I => \N__32474\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__32500\,
            I => \N__32474\
        );

    \I__6560\ : Span4Mux_v
    port map (
            O => \N__32493\,
            I => \N__32474\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__32490\,
            I => \N__32469\
        );

    \I__6558\ : Span4Mux_v
    port map (
            O => \N__32485\,
            I => \N__32469\
        );

    \I__6557\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32466\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32481\,
            I => byte_transmit_counter_4
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__32474\,
            I => byte_transmit_counter_4
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__32469\,
            I => byte_transmit_counter_4
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__32466\,
            I => byte_transmit_counter_4
        );

    \I__6552\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32450\
        );

    \I__6550\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32447\
        );

    \I__6549\ : Span4Mux_v
    port map (
            O => \N__32450\,
            I => \N__32444\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__32447\,
            I => \r_Tx_Data_0\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__32444\,
            I => \r_Tx_Data_0\
        );

    \I__6546\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32435\
        );

    \I__6545\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32432\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32429\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32432\,
            I => \c0.n10524\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__32429\,
            I => \c0.n10524\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32420\
        );

    \I__6540\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32417\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__32420\,
            I => \c0.n10550\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__32417\,
            I => \c0.n10550\
        );

    \I__6537\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32409\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__6534\ : Span4Mux_h
    port map (
            O => \N__32403\,
            I => \N__32400\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__32400\,
            I => \c0.n10746\
        );

    \I__6532\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__32394\,
            I => \c0.n6_adj_2361\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \c0.n10746_cascade_\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__32388\,
            I => \n17758_cascade_\
        );

    \I__6528\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32382\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__32382\,
            I => \c0.n10734\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__6525\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__32373\,
            I => \c0.n8_adj_2232\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__6522\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__32361\,
            I => n10_adj_2461
        );

    \I__6519\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32354\
        );

    \I__6518\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32349\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32346\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32343\
        );

    \I__6515\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32340\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__32349\,
            I => data_out_8_7
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__32346\,
            I => data_out_8_7
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__32343\,
            I => data_out_8_7
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__32340\,
            I => data_out_8_7
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__32331\,
            I => \c0.n17742_cascade_\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__32328\,
            I => \n18864_cascade_\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__32325\,
            I => \n10_adj_2529_cascade_\
        );

    \I__6507\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32318\
        );

    \I__6506\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32315\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__32318\,
            I => \N__32312\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__32315\,
            I => \r_Tx_Data_3\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__32312\,
            I => \r_Tx_Data_3\
        );

    \I__6502\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32304\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__32304\,
            I => n10_adj_2499
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__32301\,
            I => \c0.n10550_cascade_\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__32298\,
            I => \n17978_cascade_\
        );

    \I__6498\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32288\
        );

    \I__6497\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32288\
        );

    \I__6496\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32285\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__32288\,
            I => \UART_TRANSMITTER_state_7_N_1223_1\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__32285\,
            I => \UART_TRANSMITTER_state_7_N_1223_1\
        );

    \I__6493\ : InMux
    port map (
            O => \N__32280\,
            I => \N__32277\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__32277\,
            I => n18202
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__6490\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32265\
        );

    \I__6489\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32265\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__32265\,
            I => n574
        );

    \I__6487\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32259\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32253\
        );

    \I__6485\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32246\
        );

    \I__6484\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32246\
        );

    \I__6483\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32246\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__32253\,
            I => n4
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__32246\,
            I => n4
        );

    \I__6480\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32238\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__32238\,
            I => n22_adj_2522
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__6477\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32229\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__32229\,
            I => \c0.n18226\
        );

    \I__6475\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__32223\,
            I => n21_adj_2524
        );

    \I__6473\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__32217\,
            I => n6_adj_2470
        );

    \I__6471\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__32211\,
            I => n18368
        );

    \I__6469\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \c0.n18861_cascade_\
        );

    \I__6468\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32202\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32199\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__32199\,
            I => \N__32196\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__32196\,
            I => \c0.n18377\
        );

    \I__6464\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32190\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__32190\,
            I => \c0.n18019\
        );

    \I__6462\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32184\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__32184\,
            I => n129
        );

    \I__6460\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32175\
        );

    \I__6459\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32172\
        );

    \I__6458\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32169\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__32178\,
            I => \N__32165\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__32175\,
            I => \N__32161\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32172\,
            I => \N__32156\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__32169\,
            I => \N__32156\
        );

    \I__6453\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32153\
        );

    \I__6452\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32148\
        );

    \I__6451\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32148\
        );

    \I__6450\ : Odrv12
    port map (
            O => \N__32161\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__6449\ : Odrv4
    port map (
            O => \N__32156\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__32153\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__32148\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__32139\,
            I => \n129_cascade_\
        );

    \I__6445\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32133\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__32133\,
            I => \N__32126\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32121\
        );

    \I__6442\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32121\
        );

    \I__6441\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32115\
        );

    \I__6440\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32115\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__32126\,
            I => \N__32112\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__32121\,
            I => \N__32109\
        );

    \I__6437\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32106\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__32115\,
            I => \c0.tx_active\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__32112\,
            I => \c0.tx_active\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__32109\,
            I => \c0.tx_active\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__32106\,
            I => \c0.tx_active\
        );

    \I__6432\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32094\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__32091\,
            I => \c0.n1707\
        );

    \I__6429\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32084\
        );

    \I__6428\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32081\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__32084\,
            I => \c0.delay_counter_11\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__32081\,
            I => \c0.delay_counter_11\
        );

    \I__6425\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32072\
        );

    \I__6424\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32069\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__32072\,
            I => \c0.delay_counter_12\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__32069\,
            I => \c0.delay_counter_12\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__6420\ : InMux
    port map (
            O => \N__32061\,
            I => \N__32057\
        );

    \I__6419\ : InMux
    port map (
            O => \N__32060\,
            I => \N__32054\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__32057\,
            I => \N__32051\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__32054\,
            I => \c0.delay_counter_4\
        );

    \I__6416\ : Odrv12
    port map (
            O => \N__32051\,
            I => \c0.delay_counter_4\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32042\
        );

    \I__6414\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32039\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__32039\,
            I => \c0.delay_counter_7\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__32036\,
            I => \c0.delay_counter_7\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__32028\,
            I => \c0.n24\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__32025\,
            I => \N__32020\
        );

    \I__6407\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32016\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32011\
        );

    \I__6405\ : InMux
    port map (
            O => \N__32020\,
            I => \N__32011\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32008\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32003\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__32003\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__32008\,
            I => n12227
        );

    \I__6400\ : Odrv4
    port map (
            O => \N__32003\,
            I => n12227
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__31998\,
            I => \n574_cascade_\
        );

    \I__6398\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31992\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__31992\,
            I => \c0.n98\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__6395\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__31983\,
            I => \N__31980\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__31980\,
            I => \N__31977\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__31977\,
            I => \c0.n18230\
        );

    \I__6391\ : InMux
    port map (
            O => \N__31974\,
            I => \c0.n16640\
        );

    \I__6390\ : InMux
    port map (
            O => \N__31971\,
            I => \bfn_11_8_0_\
        );

    \I__6389\ : InMux
    port map (
            O => \N__31968\,
            I => \c0.n16642\
        );

    \I__6388\ : InMux
    port map (
            O => \N__31965\,
            I => \c0.n16643\
        );

    \I__6387\ : InMux
    port map (
            O => \N__31962\,
            I => \c0.n16644\
        );

    \I__6386\ : InMux
    port map (
            O => \N__31959\,
            I => \c0.n16645\
        );

    \I__6385\ : InMux
    port map (
            O => \N__31956\,
            I => \c0.n16646\
        );

    \I__6384\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31949\
        );

    \I__6383\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31946\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31943\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__31946\,
            I => \c0.delay_counter_2\
        );

    \I__6380\ : Odrv12
    port map (
            O => \N__31943\,
            I => \c0.delay_counter_2\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__31938\,
            I => \N__31935\
        );

    \I__6378\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31931\
        );

    \I__6377\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31928\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31925\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__31928\,
            I => \c0.delay_counter_5\
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__31925\,
            I => \c0.delay_counter_5\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__31920\,
            I => \N__31917\
        );

    \I__6372\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__31914\,
            I => n26_adj_2466
        );

    \I__6370\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31907\
        );

    \I__6369\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31904\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__31907\,
            I => \N__31900\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__31904\,
            I => \N__31897\
        );

    \I__6366\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31894\
        );

    \I__6365\ : Span4Mux_v
    port map (
            O => \N__31900\,
            I => \N__31889\
        );

    \I__6364\ : Span4Mux_h
    port map (
            O => \N__31897\,
            I => \N__31889\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__31894\,
            I => data_out_frame2_7_1
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__31889\,
            I => data_out_frame2_7_1
        );

    \I__6361\ : InMux
    port map (
            O => \N__31884\,
            I => \c0.n16634\
        );

    \I__6360\ : InMux
    port map (
            O => \N__31881\,
            I => \c0.n16635\
        );

    \I__6359\ : InMux
    port map (
            O => \N__31878\,
            I => \c0.n16636\
        );

    \I__6358\ : InMux
    port map (
            O => \N__31875\,
            I => \c0.n16637\
        );

    \I__6357\ : InMux
    port map (
            O => \N__31872\,
            I => \c0.n16638\
        );

    \I__6356\ : InMux
    port map (
            O => \N__31869\,
            I => \c0.n16639\
        );

    \I__6355\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31860\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__31860\,
            I => \c0.n17727\
        );

    \I__6352\ : InMux
    port map (
            O => \N__31857\,
            I => \N__31849\
        );

    \I__6351\ : InMux
    port map (
            O => \N__31856\,
            I => \N__31849\
        );

    \I__6350\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31846\
        );

    \I__6349\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31843\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31840\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__31846\,
            I => data_out_frame2_5_1
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__31843\,
            I => data_out_frame2_5_1
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__31840\,
            I => data_out_frame2_5_1
        );

    \I__6344\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31830\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__31830\,
            I => \c0.n18837\
        );

    \I__6342\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31824\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__31824\,
            I => \N__31820\
        );

    \I__6340\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31817\
        );

    \I__6339\ : Span4Mux_s0_v
    port map (
            O => \N__31820\,
            I => \N__31814\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__31817\,
            I => data_out_frame2_18_1
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__31814\,
            I => data_out_frame2_18_1
        );

    \I__6336\ : InMux
    port map (
            O => \N__31809\,
            I => \N__31806\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__31806\,
            I => \N__31802\
        );

    \I__6334\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31799\
        );

    \I__6333\ : Span4Mux_h
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__31799\,
            I => data_out_frame2_17_7
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__31796\,
            I => data_out_frame2_17_7
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__31791\,
            I => \c0.n10867_cascade_\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__31788\,
            I => \c0.n17739_cascade_\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31781\
        );

    \I__6327\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31776\
        );

    \I__6326\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31776\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__31776\,
            I => data_out_frame2_17_0
        );

    \I__6324\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__31770\,
            I => \c0.n18840\
        );

    \I__6322\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__31764\,
            I => \c0.n18795\
        );

    \I__6320\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31754\
        );

    \I__6318\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31751\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__31754\,
            I => \N__31748\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__31751\,
            I => data_out_frame2_18_7
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__31748\,
            I => data_out_frame2_18_7
        );

    \I__6314\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__31734\,
            I => \c0.n18360\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__6309\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__31722\,
            I => \c0.n18256\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__31719\,
            I => \c0.n14_adj_2359_cascade_\
        );

    \I__6305\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31713\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31713\,
            I => \c0.data_out_frame2_20_0\
        );

    \I__6303\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__31707\,
            I => \c0.n15_adj_2429\
        );

    \I__6301\ : InMux
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__31701\,
            I => \c0.n17847\
        );

    \I__6299\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31694\
        );

    \I__6298\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31691\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__31694\,
            I => \N__31688\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__31691\,
            I => data_out_2_5
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__31688\,
            I => data_out_2_5
        );

    \I__6294\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__6292\ : Odrv4
    port map (
            O => \N__31677\,
            I => \c0.n18335\
        );

    \I__6291\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31670\
        );

    \I__6290\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31667\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__31670\,
            I => \c0.data_out_2_3\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__31667\,
            I => \c0.data_out_2_3\
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__31662\,
            I => \c0.n19_cascade_\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__31659\,
            I => \N__31656\
        );

    \I__6285\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31653\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__31653\,
            I => \c0.data_out_frame2_19_1\
        );

    \I__6283\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__31647\,
            I => \c0.n20\
        );

    \I__6281\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31641\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__31641\,
            I => \N__31638\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__31638\,
            I => \c0.n18266\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__31635\,
            I => \n10_adj_2528_cascade_\
        );

    \I__6277\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31629\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__31629\,
            I => \N__31625\
        );

    \I__6275\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__31622\,
            I => \r_Tx_Data_2\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__31619\,
            I => \r_Tx_Data_2\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__31614\,
            I => \N__31611\
        );

    \I__6270\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31607\
        );

    \I__6269\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31604\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__31607\,
            I => data_out_3_5
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__31604\,
            I => data_out_3_5
        );

    \I__6266\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31595\
        );

    \I__6265\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31592\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__31595\,
            I => data_out_1_6
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__31592\,
            I => data_out_1_6
        );

    \I__6262\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31581\
        );

    \I__6261\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31581\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__31581\,
            I => \c0.data_out_0_6\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__31578\,
            I => \N__31575\
        );

    \I__6258\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31572\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__31572\,
            I => \N__31569\
        );

    \I__6256\ : Span4Mux_v
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__31566\,
            I => \c0.n1_adj_2272\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__6253\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__31557\,
            I => \c0.n5_adj_2241\
        );

    \I__6251\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31551\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__31551\,
            I => \c0.n18753\
        );

    \I__6249\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__31542\,
            I => \c0.n2\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__31539\,
            I => \N__31536\
        );

    \I__6245\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31533\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__31530\,
            I => \N__31527\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__31527\,
            I => \c0.n18189\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \n18876_cascade_\
        );

    \I__6240\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__31518\,
            I => n10_adj_2531
        );

    \I__6238\ : CascadeMux
    port map (
            O => \N__31515\,
            I => \c0.n5_adj_2196_cascade_\
        );

    \I__6237\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__31509\,
            I => \c0.n18873\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__31506\,
            I => \n5_cascade_\
        );

    \I__6234\ : CascadeMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__6233\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__31497\,
            I => \c0.n8_adj_2209\
        );

    \I__6231\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__31491\,
            I => n10_adj_2533
        );

    \I__6229\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31482\
        );

    \I__6228\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31479\
        );

    \I__6227\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31474\
        );

    \I__6226\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31474\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__31482\,
            I => \r_Bit_Index_1\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__31479\,
            I => \r_Bit_Index_1\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__31474\,
            I => \r_Bit_Index_1\
        );

    \I__6222\ : InMux
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__31464\,
            I => \c0.tx.n18167\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__31461\,
            I => \N__31456\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__31460\,
            I => \N__31452\
        );

    \I__6218\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31449\
        );

    \I__6217\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31446\
        );

    \I__6216\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31441\
        );

    \I__6215\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31441\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__31449\,
            I => \r_Bit_Index_2\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31446\,
            I => \r_Bit_Index_2\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__31441\,
            I => \r_Bit_Index_2\
        );

    \I__6211\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31431\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__31431\,
            I => \c0.tx.n18711\
        );

    \I__6209\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31424\
        );

    \I__6208\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31421\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31418\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__31421\,
            I => \r_Tx_Data_1\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__31418\,
            I => \r_Tx_Data_1\
        );

    \I__6204\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__31410\,
            I => \c0.tx.n18040\
        );

    \I__6202\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__31404\,
            I => \c0.n8_adj_2205\
        );

    \I__6200\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31392\
        );

    \I__6199\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31387\
        );

    \I__6198\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31387\
        );

    \I__6197\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31384\
        );

    \I__6196\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31381\
        );

    \I__6195\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31374\
        );

    \I__6194\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31374\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31365\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__31387\,
            I => \N__31365\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__31384\,
            I => \N__31365\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__31381\,
            I => \N__31365\
        );

    \I__6189\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31362\
        );

    \I__6188\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31359\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__31374\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__31365\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__31362\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__31359\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__6183\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31337\
        );

    \I__6182\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31337\
        );

    \I__6181\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31337\
        );

    \I__6180\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31334\
        );

    \I__6179\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31331\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__31345\,
            I => \N__31328\
        );

    \I__6177\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31322\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31315\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__31334\,
            I => \N__31315\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31315\
        );

    \I__6173\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31308\
        );

    \I__6172\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31308\
        );

    \I__6171\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31308\
        );

    \I__6170\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31305\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__31322\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__31315\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__31308\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__31305\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__31296\,
            I => \N__31286\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__31295\,
            I => \N__31282\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__31294\,
            I => \N__31279\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__31293\,
            I => \N__31276\
        );

    \I__6161\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31272\
        );

    \I__6160\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31269\
        );

    \I__6159\ : CascadeMux
    port map (
            O => \N__31290\,
            I => \N__31266\
        );

    \I__6158\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31261\
        );

    \I__6157\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31261\
        );

    \I__6156\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31258\
        );

    \I__6155\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31253\
        );

    \I__6154\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31253\
        );

    \I__6153\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31247\
        );

    \I__6152\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31247\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31242\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31242\
        );

    \I__6149\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31239\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__31261\,
            I => \N__31232\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__31258\,
            I => \N__31232\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31232\
        );

    \I__6145\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31229\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__31247\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__31242\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__31239\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__31232\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__31229\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__6139\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31208\
        );

    \I__6138\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31208\
        );

    \I__6137\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31202\
        );

    \I__6136\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31202\
        );

    \I__6135\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31197\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31197\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31194\
        );

    \I__6132\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31191\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__31202\,
            I => \N__31188\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31181\
        );

    \I__6129\ : Span4Mux_v
    port map (
            O => \N__31194\,
            I => \N__31181\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31181\
        );

    \I__6127\ : Span4Mux_v
    port map (
            O => \N__31188\,
            I => \N__31178\
        );

    \I__6126\ : Span4Mux_h
    port map (
            O => \N__31181\,
            I => \N__31175\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__31178\,
            I => \c0.tx.r_SM_Main_2_N_2031_1\
        );

    \I__6124\ : Odrv4
    port map (
            O => \N__31175\,
            I => \c0.tx.r_SM_Main_2_N_2031_1\
        );

    \I__6123\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31161\
        );

    \I__6122\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31161\
        );

    \I__6121\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31161\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__31158\,
            I => n18012
        );

    \I__6118\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31145\
        );

    \I__6117\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31142\
        );

    \I__6116\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31137\
        );

    \I__6115\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31137\
        );

    \I__6114\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31134\
        );

    \I__6113\ : InMux
    port map (
            O => \N__31150\,
            I => \N__31129\
        );

    \I__6112\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31129\
        );

    \I__6111\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31126\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__31145\,
            I => \N__31121\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31121\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__31137\,
            I => \r_Bit_Index_0\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__31134\,
            I => \r_Bit_Index_0\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__31129\,
            I => \r_Bit_Index_0\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__31126\,
            I => \r_Bit_Index_0\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__31121\,
            I => \r_Bit_Index_0\
        );

    \I__6103\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31104\
        );

    \I__6102\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31104\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__31104\,
            I => \r_Tx_Data_5\
        );

    \I__6100\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__31098\,
            I => \c0.tx.n18166\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__31095\,
            I => \n5440_cascade_\
        );

    \I__6097\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31089\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__31089\,
            I => n18016
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__31086\,
            I => \n18016_cascade_\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__31077\,
            I => \c0.n8_adj_2207\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31070\
        );

    \I__6090\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31067\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__31070\,
            I => \c0.tx.n13802\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__31067\,
            I => \c0.tx.n13802\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__31062\,
            I => \c0.tx.n13802_cascade_\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__31059\,
            I => \c0.tx.n6796_cascade_\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__31056\,
            I => \c0.n4_cascade_\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__31053\,
            I => \n5341_cascade_\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__31047\,
            I => \N__31043\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31040\
        );

    \I__6080\ : Odrv4
    port map (
            O => \N__31043\,
            I => \tx_transmit_N_1947_7\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__31040\,
            I => \tx_transmit_N_1947_7\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31031\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31028\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__31031\,
            I => \N__31025\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__31028\,
            I => byte_transmit_counter_7
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__31025\,
            I => byte_transmit_counter_7
        );

    \I__6073\ : InMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31013\
        );

    \I__6071\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31010\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__31013\,
            I => \c0.tx_transmit_N_1947_5\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__31010\,
            I => \c0.tx_transmit_N_1947_5\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__31005\,
            I => \N__30997\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__31004\,
            I => \N__30994\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__31003\,
            I => \N__30990\
        );

    \I__6065\ : CascadeMux
    port map (
            O => \N__31002\,
            I => \N__30986\
        );

    \I__6064\ : CascadeMux
    port map (
            O => \N__31001\,
            I => \N__30983\
        );

    \I__6063\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30979\
        );

    \I__6062\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30968\
        );

    \I__6061\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30968\
        );

    \I__6060\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30968\
        );

    \I__6059\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30968\
        );

    \I__6058\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30968\
        );

    \I__6057\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30961\
        );

    \I__6056\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30961\
        );

    \I__6055\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30961\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__30979\,
            I => n10973
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__30968\,
            I => n10973
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__30961\,
            I => n10973
        );

    \I__6051\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30943\
        );

    \I__6050\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30943\
        );

    \I__6049\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30932\
        );

    \I__6048\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30932\
        );

    \I__6047\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30932\
        );

    \I__6046\ : InMux
    port map (
            O => \N__30949\,
            I => \N__30932\
        );

    \I__6045\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30932\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__30943\,
            I => n5341
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__30932\,
            I => n5341
        );

    \I__6042\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30923\
        );

    \I__6041\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30920\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__30923\,
            I => \N__30917\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__30920\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__30917\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__6037\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__30909\,
            I => \c0.n17998\
        );

    \I__6035\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30903\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__30900\,
            I => \c0.tx.n17938\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__6031\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__30891\,
            I => n10_adj_2536
        );

    \I__6029\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30884\
        );

    \I__6028\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30881\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__30884\,
            I => byte_transmit_counter_6
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__30881\,
            I => byte_transmit_counter_6
        );

    \I__6025\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30870\
        );

    \I__6024\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30870\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__30870\,
            I => \tx_transmit_N_1947_6\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__30867\,
            I => \N__30863\
        );

    \I__6021\ : InMux
    port map (
            O => \N__30866\,
            I => \N__30858\
        );

    \I__6020\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30858\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__30858\,
            I => \tx_transmit_N_1947_4\
        );

    \I__6018\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30850\
        );

    \I__6017\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30847\
        );

    \I__6016\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30844\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__30850\,
            I => \N__30841\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__30847\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__30844\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__30841\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__30834\,
            I => \c0.tx2.n10_cascade_\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__30831\,
            I => \N__30826\
        );

    \I__6009\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30823\
        );

    \I__6008\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30820\
        );

    \I__6007\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30817\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__30823\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__30820\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__30817\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__6003\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30807\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__6001\ : Sp12to4
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__6000\ : Odrv12
    port map (
            O => \N__30801\,
            I => \c0.tx2.n12775\
        );

    \I__5999\ : InMux
    port map (
            O => \N__30798\,
            I => \N__30795\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__30795\,
            I => \N__30792\
        );

    \I__5997\ : Odrv12
    port map (
            O => \N__30792\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__5996\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30786\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__30786\,
            I => \c0.tx2.n18061\
        );

    \I__5994\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30778\
        );

    \I__5993\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30775\
        );

    \I__5992\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30770\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30766\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__30775\,
            I => \N__30763\
        );

    \I__5989\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30758\
        );

    \I__5988\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30755\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__30770\,
            I => \N__30752\
        );

    \I__5986\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30749\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__30766\,
            I => \N__30744\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__30763\,
            I => \N__30744\
        );

    \I__5983\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30739\
        );

    \I__5982\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30739\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__30758\,
            I => \r_SM_Main_2\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__30755\,
            I => \r_SM_Main_2\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__30752\,
            I => \r_SM_Main_2\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__30749\,
            I => \r_SM_Main_2\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__30744\,
            I => \r_SM_Main_2\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__30739\,
            I => \r_SM_Main_2\
        );

    \I__5975\ : CEMux
    port map (
            O => \N__30726\,
            I => \N__30721\
        );

    \I__5974\ : CEMux
    port map (
            O => \N__30725\,
            I => \N__30718\
        );

    \I__5973\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30715\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30712\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30709\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30706\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__30712\,
            I => n11096
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__30709\,
            I => n11096
        );

    \I__5967\ : Odrv12
    port map (
            O => \N__30706\,
            I => n11096
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__30699\,
            I => \c0.n18260_cascade_\
        );

    \I__5965\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__30693\,
            I => \c0.n130\
        );

    \I__5963\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__30687\,
            I => \c0.n3465\
        );

    \I__5961\ : SRMux
    port map (
            O => \N__30684\,
            I => \N__30681\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30678\
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__30678\,
            I => \c0.n4806\
        );

    \I__5958\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__30666\,
            I => \c0.n18362\
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__30663\,
            I => \N__30660\
        );

    \I__5953\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30654\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__30659\,
            I => \N__30651\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__30658\,
            I => \N__30647\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__30657\,
            I => \N__30644\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__30654\,
            I => \N__30639\
        );

    \I__5948\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30636\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__30650\,
            I => \N__30633\
        );

    \I__5946\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30630\
        );

    \I__5945\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30627\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__30643\,
            I => \N__30624\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__30642\,
            I => \N__30621\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__30639\,
            I => \N__30618\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30615\
        );

    \I__5940\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30612\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30607\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30607\
        );

    \I__5937\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30604\
        );

    \I__5936\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30601\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__30618\,
            I => \N__30592\
        );

    \I__5934\ : Span4Mux_s0_v
    port map (
            O => \N__30615\,
            I => \N__30592\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30592\
        );

    \I__5932\ : Span4Mux_s2_v
    port map (
            O => \N__30607\,
            I => \N__30587\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__30604\,
            I => \N__30587\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__30601\,
            I => \N__30584\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__30600\,
            I => \N__30581\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__30599\,
            I => \N__30578\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__30592\,
            I => \N__30575\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__30587\,
            I => \N__30570\
        );

    \I__5925\ : Span4Mux_v
    port map (
            O => \N__30584\,
            I => \N__30570\
        );

    \I__5924\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30567\
        );

    \I__5923\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30564\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__30575\,
            I => \c0.n12359\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__30570\,
            I => \c0.n12359\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__30567\,
            I => \c0.n12359\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__30564\,
            I => \c0.n12359\
        );

    \I__5918\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30548\
        );

    \I__5917\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30543\
        );

    \I__5916\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30540\
        );

    \I__5915\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30537\
        );

    \I__5914\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30534\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30531\
        );

    \I__5912\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30528\
        );

    \I__5911\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30525\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30520\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30520\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30512\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__30534\,
            I => \N__30512\
        );

    \I__5906\ : Span4Mux_s0_v
    port map (
            O => \N__30531\,
            I => \N__30505\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30505\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N__30505\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__30520\,
            I => \N__30502\
        );

    \I__5902\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30499\
        );

    \I__5901\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30496\
        );

    \I__5900\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30493\
        );

    \I__5899\ : Span12Mux_s4_v
    port map (
            O => \N__30512\,
            I => \N__30489\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__30505\,
            I => \N__30484\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__30502\,
            I => \N__30484\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__30499\,
            I => \N__30481\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30478\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__30493\,
            I => \N__30475\
        );

    \I__5893\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30472\
        );

    \I__5892\ : Odrv12
    port map (
            O => \N__30489\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__30484\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__30481\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__30478\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__30475\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__30472\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__5886\ : SRMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5884\ : Odrv12
    port map (
            O => \N__30453\,
            I => \c0.n4_adj_2204\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30444\
        );

    \I__5882\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30444\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__30444\,
            I => \c0.tx2.n13800\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__30441\,
            I => \N__30431\
        );

    \I__5879\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30427\
        );

    \I__5878\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30424\
        );

    \I__5877\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30417\
        );

    \I__5876\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30417\
        );

    \I__5875\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30417\
        );

    \I__5874\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30407\
        );

    \I__5873\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30407\
        );

    \I__5872\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30407\
        );

    \I__5871\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30407\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30404\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30399\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30399\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30396\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30393\
        );

    \I__5865\ : Span4Mux_v
    port map (
            O => \N__30404\,
            I => \N__30388\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__30399\,
            I => \N__30388\
        );

    \I__5863\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30385\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__30393\,
            I => \N__30382\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__30388\,
            I => \N__30379\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__30385\,
            I => \r_SM_Main_1\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__30382\,
            I => \r_SM_Main_1\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__30379\,
            I => \r_SM_Main_1\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30363\
        );

    \I__5855\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30360\
        );

    \I__5854\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30357\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30352\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__30363\,
            I => \N__30349\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__30360\,
            I => \N__30344\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__30357\,
            I => \N__30344\
        );

    \I__5849\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30341\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__30355\,
            I => \N__30336\
        );

    \I__5847\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30333\
        );

    \I__5846\ : Span4Mux_s2_v
    port map (
            O => \N__30349\,
            I => \N__30330\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__30344\,
            I => \N__30327\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30324\
        );

    \I__5843\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30317\
        );

    \I__5842\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30317\
        );

    \I__5841\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30317\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__30333\,
            I => \r_SM_Main_0\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__30330\,
            I => \r_SM_Main_0\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__30327\,
            I => \r_SM_Main_0\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__30324\,
            I => \r_SM_Main_0\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__30317\,
            I => \r_SM_Main_0\
        );

    \I__5835\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__30297\,
            I => n3
        );

    \I__5831\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30291\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__5829\ : Span12Mux_s7_v
    port map (
            O => \N__30288\,
            I => \N__30285\
        );

    \I__5828\ : Odrv12
    port map (
            O => \N__30285\,
            I => \c0.tx2.n18164\
        );

    \I__5827\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__30279\,
            I => \N__30276\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__30276\,
            I => \N__30273\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__30273\,
            I => \N__30270\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__30270\,
            I => \c0.tx2.n18163\
        );

    \I__5822\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__30264\,
            I => \c0.tx2.n18062\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__30261\,
            I => \c0.tx2.n18717_cascade_\
        );

    \I__5819\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__30255\,
            I => \c0.tx2.o_Tx_Serial_N_2062\
        );

    \I__5817\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30248\
        );

    \I__5816\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30245\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__30248\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__30245\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__5813\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30236\
        );

    \I__5812\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30233\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__30236\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__30233\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__30228\,
            I => \N__30224\
        );

    \I__5808\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30221\
        );

    \I__5807\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30218\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__30221\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__30218\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__5804\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30209\
        );

    \I__5803\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30206\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__30209\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__30206\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__5800\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__5798\ : Odrv4
    port map (
            O => \N__30195\,
            I => \c0.tx2.n10\
        );

    \I__5797\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30188\
        );

    \I__5796\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30185\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30181\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30178\
        );

    \I__5793\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30175\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__30181\,
            I => \N__30172\
        );

    \I__5791\ : Span4Mux_h
    port map (
            O => \N__30178\,
            I => \N__30169\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30175\,
            I => tx2_active
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__30172\,
            I => tx2_active
        );

    \I__5788\ : Odrv4
    port map (
            O => \N__30169\,
            I => tx2_active
        );

    \I__5787\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30158\
        );

    \I__5786\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30155\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__30158\,
            I => \N__30150\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__30155\,
            I => \N__30150\
        );

    \I__5783\ : Span4Mux_h
    port map (
            O => \N__30150\,
            I => \N__30146\
        );

    \I__5782\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30143\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__30146\,
            I => \c0.n14064\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__30143\,
            I => \c0.n14064\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__30138\,
            I => \c0.n12359_cascade_\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__30135\,
            I => \c0.n6_adj_2443_cascade_\
        );

    \I__5777\ : InMux
    port map (
            O => \N__30132\,
            I => \N__30128\
        );

    \I__5776\ : SRMux
    port map (
            O => \N__30131\,
            I => \N__30125\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__30128\,
            I => \N__30121\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30118\
        );

    \I__5773\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30115\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__30121\,
            I => \N__30105\
        );

    \I__5771\ : Sp12to4
    port map (
            O => \N__30118\,
            I => \N__30100\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__30115\,
            I => \N__30100\
        );

    \I__5769\ : InMux
    port map (
            O => \N__30114\,
            I => \N__30097\
        );

    \I__5768\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30090\
        );

    \I__5767\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30090\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30090\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30083\
        );

    \I__5764\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30083\
        );

    \I__5763\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30083\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__30105\,
            I => \c0.n10513\
        );

    \I__5761\ : Odrv12
    port map (
            O => \N__30100\,
            I => \c0.n10513\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__30097\,
            I => \c0.n10513\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__30090\,
            I => \c0.n10513\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__30083\,
            I => \c0.n10513\
        );

    \I__5757\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30061\
        );

    \I__5756\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30061\
        );

    \I__5755\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30058\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30051\
        );

    \I__5753\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30051\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30051\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__30066\,
            I => \N__30046\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__30061\,
            I => \N__30036\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__30036\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__30036\
        );

    \I__5747\ : InMux
    port map (
            O => \N__30050\,
            I => \N__30031\
        );

    \I__5746\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30026\
        );

    \I__5745\ : InMux
    port map (
            O => \N__30046\,
            I => \N__30026\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30023\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__30044\,
            I => \N__30018\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__30043\,
            I => \N__30015\
        );

    \I__5741\ : Span4Mux_h
    port map (
            O => \N__30036\,
            I => \N__30012\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30008\
        );

    \I__5739\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30004\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__29997\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__30026\,
            I => \N__29997\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__30023\,
            I => \N__29997\
        );

    \I__5735\ : InMux
    port map (
            O => \N__30022\,
            I => \N__29990\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30021\,
            I => \N__29990\
        );

    \I__5733\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29990\
        );

    \I__5732\ : InMux
    port map (
            O => \N__30015\,
            I => \N__29987\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__30012\,
            I => \N__29984\
        );

    \I__5730\ : InMux
    port map (
            O => \N__30011\,
            I => \N__29979\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30008\,
            I => \N__29974\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29974\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__30004\,
            I => \N__29967\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__29997\,
            I => \N__29967\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29967\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__29987\,
            I => \N__29962\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__29984\,
            I => \N__29962\
        );

    \I__5722\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29957\
        );

    \I__5721\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29957\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29950\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__29974\,
            I => \N__29950\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__29967\,
            I => \N__29950\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__29962\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__29957\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__29950\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__29943\,
            I => \N__29940\
        );

    \I__5713\ : InMux
    port map (
            O => \N__29940\,
            I => \N__29937\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__29937\,
            I => \N__29934\
        );

    \I__5711\ : Span12Mux_v
    port map (
            O => \N__29934\,
            I => \N__29931\
        );

    \I__5710\ : Odrv12
    port map (
            O => \N__29931\,
            I => \c0.n10958\
        );

    \I__5709\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29922\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__29927\,
            I => \N__29919\
        );

    \I__5707\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29913\
        );

    \I__5706\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29913\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29910\
        );

    \I__5704\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29907\
        );

    \I__5703\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29904\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__29913\,
            I => \N__29901\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__29910\,
            I => \N__29898\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__29907\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2213\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__29904\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2213\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__29901\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2213\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__29898\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2213\
        );

    \I__5696\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29886\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29883\
        );

    \I__5694\ : Span4Mux_s3_v
    port map (
            O => \N__29883\,
            I => \N__29880\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__29880\,
            I => n6707
        );

    \I__5692\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29873\
        );

    \I__5691\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29870\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__29873\,
            I => \N__29867\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__29870\,
            I => \N__29864\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__29867\,
            I => \N__29861\
        );

    \I__5687\ : Span12Mux_s7_v
    port map (
            O => \N__29864\,
            I => \N__29858\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__29861\,
            I => \N__29855\
        );

    \I__5685\ : Odrv12
    port map (
            O => \N__29858\,
            I => \c0.tx2.n12769\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__29855\,
            I => \c0.tx2.n12769\
        );

    \I__5683\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29846\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__29849\,
            I => \N__29843\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29838\
        );

    \I__5680\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29835\
        );

    \I__5679\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29832\
        );

    \I__5678\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29829\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__29838\,
            I => \N__29825\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29818\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29818\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__29829\,
            I => \N__29818\
        );

    \I__5673\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29815\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__29825\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__29818\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__29815\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__29808\,
            I => \r_SM_Main_2_N_2031_1_cascade_\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__29805\,
            I => \n18014_cascade_\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__29802\,
            I => \c0.n5_adj_2435_cascade_\
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__5665\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__29790\,
            I => \c0.n6_adj_2223\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__29787\,
            I => \c0.n18687_cascade_\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__5660\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__29775\,
            I => \c0.n18690\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__29772\,
            I => \N__29769\
        );

    \I__5656\ : InMux
    port map (
            O => \N__29769\,
            I => \N__29766\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__29763\,
            I => \N__29760\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__29757\,
            I => \c0.n5_adj_2197\
        );

    \I__5651\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__5649\ : Span12Mux_s3_v
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__5648\ : Odrv12
    port map (
            O => \N__29745\,
            I => \c0.n6\
        );

    \I__5647\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__29736\,
            I => \c0.n6_adj_2354\
        );

    \I__5644\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29730\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__29730\,
            I => \c0.n18855\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__29727\,
            I => \c0.n10893_cascade_\
        );

    \I__5641\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29720\
        );

    \I__5640\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29717\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__29720\,
            I => \N__29714\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__29717\,
            I => data_out_frame2_17_1
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__29714\,
            I => data_out_frame2_17_1
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__29709\,
            I => \c0.n18888_cascade_\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__29706\,
            I => \c0.n18789_cascade_\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__29703\,
            I => \c0.n18792_cascade_\
        );

    \I__5633\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29697\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__29697\,
            I => \c0.n22_adj_2270\
        );

    \I__5631\ : InMux
    port map (
            O => \N__29694\,
            I => \N__29691\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__29691\,
            I => \c0.n18885\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__29688\,
            I => \c0.n10861_cascade_\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__5627\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__29679\,
            I => \c0.n18798\
        );

    \I__5625\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29672\
        );

    \I__5624\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29669\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__29672\,
            I => \control.pwm_delay_2\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__29669\,
            I => \control.pwm_delay_2\
        );

    \I__5621\ : InMux
    port map (
            O => \N__29664\,
            I => \control.n16648\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__29661\,
            I => \N__29657\
        );

    \I__5619\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29654\
        );

    \I__5618\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29651\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__29654\,
            I => \control.pwm_delay_3\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__29651\,
            I => \control.pwm_delay_3\
        );

    \I__5615\ : InMux
    port map (
            O => \N__29646\,
            I => \control.n16649\
        );

    \I__5614\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29639\
        );

    \I__5613\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29636\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__29639\,
            I => \control.pwm_delay_4\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__29636\,
            I => \control.pwm_delay_4\
        );

    \I__5610\ : InMux
    port map (
            O => \N__29631\,
            I => \control.n16650\
        );

    \I__5609\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29624\
        );

    \I__5608\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29621\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__29624\,
            I => \control.pwm_delay_5\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__29621\,
            I => \control.pwm_delay_5\
        );

    \I__5605\ : InMux
    port map (
            O => \N__29616\,
            I => \control.n16651\
        );

    \I__5604\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29609\
        );

    \I__5603\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29606\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__29609\,
            I => \control.pwm_delay_6\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__29606\,
            I => \control.pwm_delay_6\
        );

    \I__5600\ : InMux
    port map (
            O => \N__29601\,
            I => \control.n16652\
        );

    \I__5599\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29594\
        );

    \I__5598\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29591\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__29594\,
            I => \control.pwm_delay_7\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__29591\,
            I => \control.pwm_delay_7\
        );

    \I__5595\ : InMux
    port map (
            O => \N__29586\,
            I => \control.n16653\
        );

    \I__5594\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29579\
        );

    \I__5593\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29576\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29573\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__29576\,
            I => \control.pwm_delay_8\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__29573\,
            I => \control.pwm_delay_8\
        );

    \I__5589\ : InMux
    port map (
            O => \N__29568\,
            I => \bfn_9_24_0_\
        );

    \I__5588\ : InMux
    port map (
            O => \N__29565\,
            I => \control.n16655\
        );

    \I__5587\ : CascadeMux
    port map (
            O => \N__29562\,
            I => \N__29559\
        );

    \I__5586\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29553\
        );

    \I__5585\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29553\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__29553\,
            I => data_out_3_7
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__5582\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29541\
        );

    \I__5581\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29541\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__29541\,
            I => data_out_2_7
        );

    \I__5579\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__29535\,
            I => \N__29532\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__29532\,
            I => \c0.n2_adj_2229\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__29529\,
            I => \n2837_cascade_\
        );

    \I__5575\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29522\
        );

    \I__5574\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29519\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__29522\,
            I => data_out_0_5
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__29519\,
            I => data_out_0_5
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__29514\,
            I => \control.n12_cascade_\
        );

    \I__5570\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__29508\,
            I => \control.n10\
        );

    \I__5568\ : InMux
    port map (
            O => \N__29505\,
            I => \bfn_9_23_0_\
        );

    \I__5567\ : InMux
    port map (
            O => \N__29502\,
            I => \N__29499\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__29499\,
            I => \control.n9_adj_2459\
        );

    \I__5565\ : InMux
    port map (
            O => \N__29496\,
            I => \control.n16647\
        );

    \I__5564\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__29490\,
            I => \N__29487\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__29487\,
            I => \c0.n18188\
        );

    \I__5561\ : CEMux
    port map (
            O => \N__29484\,
            I => \N__29480\
        );

    \I__5560\ : CEMux
    port map (
            O => \N__29483\,
            I => \N__29476\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__29480\,
            I => \N__29473\
        );

    \I__5558\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29469\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__29476\,
            I => \N__29466\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__29473\,
            I => \N__29463\
        );

    \I__5555\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29460\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__29469\,
            I => \N__29457\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__29466\,
            I => \N__29450\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__29463\,
            I => \N__29450\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29450\
        );

    \I__5550\ : Odrv12
    port map (
            O => \N__29457\,
            I => n5155
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__29450\,
            I => n5155
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__5547\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__29436\,
            I => \c0.n18354\
        );

    \I__5544\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__29430\,
            I => n18756
        );

    \I__5542\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29423\
        );

    \I__5541\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29420\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29417\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__29420\,
            I => \c0.data_out_3_6\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__29417\,
            I => \c0.data_out_3_6\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__29412\,
            I => \n10_adj_2532_cascade_\
        );

    \I__5536\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29403\
        );

    \I__5535\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29403\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__29403\,
            I => \r_Tx_Data_6\
        );

    \I__5533\ : InMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__29391\,
            I => \c0.tx.n17984\
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__29388\,
            I => \n10_adj_2537_cascade_\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__29385\,
            I => \n10_adj_2535_cascade_\
        );

    \I__5527\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29378\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29375\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__29378\,
            I => \r_Tx_Data_7\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__29375\,
            I => \r_Tx_Data_7\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__29370\,
            I => \n3_adj_2525_cascade_\
        );

    \I__5522\ : IoInMux
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__29364\,
            I => \N__29361\
        );

    \I__5520\ : Span4Mux_s3_h
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__29358\,
            I => \N__29355\
        );

    \I__5518\ : Span4Mux_v
    port map (
            O => \N__29355\,
            I => \N__29350\
        );

    \I__5517\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29347\
        );

    \I__5516\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29344\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__29350\,
            I => \N__29341\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__29347\,
            I => \N__29338\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29335\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__29341\,
            I => tx_o
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__29338\,
            I => tx_o
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__29335\,
            I => tx_o
        );

    \I__5509\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29325\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__29325\,
            I => \c0.tx.n17697\
        );

    \I__5507\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29318\
        );

    \I__5506\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29315\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__29318\,
            I => data_out_1_7
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__29315\,
            I => data_out_1_7
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__29310\,
            I => \c0.tx.n11030_cascade_\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__29304\,
            I => \c0.tx.n18041\
        );

    \I__5500\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__29298\,
            I => \c0.tx.o_Tx_Serial_N_2062\
        );

    \I__5498\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29292\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__29292\,
            I => n18750
        );

    \I__5496\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__29286\,
            I => \c0.tx_active_prev\
        );

    \I__5494\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__29280\,
            I => \N__29275\
        );

    \I__5492\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29271\
        );

    \I__5491\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29268\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__29275\,
            I => \N__29265\
        );

    \I__5489\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29262\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29257\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29257\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__29265\,
            I => data_in_1_1
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__29262\,
            I => data_in_1_1
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__29257\,
            I => data_in_1_1
        );

    \I__5483\ : InMux
    port map (
            O => \N__29250\,
            I => \c0.n16520\
        );

    \I__5482\ : InMux
    port map (
            O => \N__29247\,
            I => \c0.n16521\
        );

    \I__5481\ : InMux
    port map (
            O => \N__29244\,
            I => \c0.n16522\
        );

    \I__5480\ : InMux
    port map (
            O => \N__29241\,
            I => \c0.n16523\
        );

    \I__5479\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__29226\,
            I => \c0.n18254\
        );

    \I__5474\ : SRMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29217\
        );

    \I__5472\ : Sp12to4
    port map (
            O => \N__29217\,
            I => \N__29214\
        );

    \I__5471\ : Span12Mux_v
    port map (
            O => \N__29214\,
            I => \N__29211\
        );

    \I__5470\ : Odrv12
    port map (
            O => \N__29211\,
            I => \c0.n4_adj_2231\
        );

    \I__5469\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29205\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__29205\,
            I => \N__29201\
        );

    \I__5467\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29197\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__29201\,
            I => \N__29194\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29191\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29186\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__29194\,
            I => \N__29186\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__29191\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__29186\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__5460\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29178\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__29178\,
            I => \N__29174\
        );

    \I__5458\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29170\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__29174\,
            I => \N__29167\
        );

    \I__5456\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29164\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29159\
        );

    \I__5454\ : Span4Mux_v
    port map (
            O => \N__29167\,
            I => \N__29159\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__29164\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__29159\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__5451\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__29151\,
            I => \N__29147\
        );

    \I__5449\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__29147\,
            I => \N__29138\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__29144\,
            I => \N__29138\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29135\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__29138\,
            I => \N__29130\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__29135\,
            I => \N__29130\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__29130\,
            I => \c0.rx.n73\
        );

    \I__5442\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__29124\,
            I => \c0.n44\
        );

    \I__5440\ : IoInMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__5438\ : IoSpan4Mux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__5437\ : IoSpan4Mux
    port map (
            O => \N__29112\,
            I => \N__29109\
        );

    \I__5436\ : Span4Mux_s3_h
    port map (
            O => \N__29109\,
            I => \N__29106\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__29103\,
            I => tx_enable
        );

    \I__5433\ : InMux
    port map (
            O => \N__29100\,
            I => \c0.tx2.n16542\
        );

    \I__5432\ : InMux
    port map (
            O => \N__29097\,
            I => \c0.tx2.n16543\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29091\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29088\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__29088\,
            I => \N__29084\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29081\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__29084\,
            I => \N__29078\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__29081\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__29078\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__5424\ : InMux
    port map (
            O => \N__29073\,
            I => \c0.tx2.n16544\
        );

    \I__5423\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29067\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__29067\,
            I => \N__29064\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__29064\,
            I => \N__29060\
        );

    \I__5420\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29057\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__29060\,
            I => \N__29054\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__29057\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__29054\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__5416\ : InMux
    port map (
            O => \N__29049\,
            I => \c0.tx2.n16545\
        );

    \I__5415\ : InMux
    port map (
            O => \N__29046\,
            I => \bfn_9_7_0_\
        );

    \I__5414\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__29037\,
            I => \N__29033\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29030\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__29033\,
            I => \N__29027\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__29030\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__29027\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__5407\ : SRMux
    port map (
            O => \N__29022\,
            I => \N__29018\
        );

    \I__5406\ : SRMux
    port map (
            O => \N__29021\,
            I => \N__29015\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__29018\,
            I => \N__29012\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29015\,
            I => \N__29009\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__29012\,
            I => \N__29006\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__29009\,
            I => \N__29003\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__29006\,
            I => \c0.tx2.n11312\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__29003\,
            I => \c0.tx2.n11312\
        );

    \I__5399\ : InMux
    port map (
            O => \N__28998\,
            I => \c0.n16517\
        );

    \I__5398\ : InMux
    port map (
            O => \N__28995\,
            I => \c0.n16518\
        );

    \I__5397\ : InMux
    port map (
            O => \N__28992\,
            I => \c0.n16519\
        );

    \I__5396\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28977\
        );

    \I__5395\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28977\
        );

    \I__5394\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28974\
        );

    \I__5393\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28971\
        );

    \I__5392\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28968\
        );

    \I__5391\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28961\
        );

    \I__5390\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28961\
        );

    \I__5389\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28961\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28958\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28949\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28949\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28949\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28949\
        );

    \I__5383\ : Span4Mux_h
    port map (
            O => \N__28958\,
            I => \N__28946\
        );

    \I__5382\ : Span12Mux_s4_v
    port map (
            O => \N__28949\,
            I => \N__28943\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__28946\,
            I => \c0.n6033\
        );

    \I__5380\ : Odrv12
    port map (
            O => \N__28943\,
            I => \c0.n6033\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__28938\,
            I => \c0.n18085_cascade_\
        );

    \I__5378\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28930\
        );

    \I__5377\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28925\
        );

    \I__5376\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28925\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28921\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__28925\,
            I => \N__28916\
        );

    \I__5373\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28913\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__28921\,
            I => \N__28910\
        );

    \I__5371\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28905\
        );

    \I__5370\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28905\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__28916\,
            I => \N__28900\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28900\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__28910\,
            I => \c0.n4494\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__28905\,
            I => \c0.n4494\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__28900\,
            I => \c0.n4494\
        );

    \I__5364\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28887\
        );

    \I__5363\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28887\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__28884\,
            I => \N__28879\
        );

    \I__5360\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28874\
        );

    \I__5359\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28874\
        );

    \I__5358\ : Odrv4
    port map (
            O => \N__28879\,
            I => \c0.n28\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__28874\,
            I => \c0.n28\
        );

    \I__5356\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28863\
        );

    \I__5355\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28863\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28855\
        );

    \I__5353\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28850\
        );

    \I__5352\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28850\
        );

    \I__5351\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28843\
        );

    \I__5350\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28843\
        );

    \I__5349\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28843\
        );

    \I__5348\ : Odrv4
    port map (
            O => \N__28855\,
            I => \c0.n12704\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__28850\,
            I => \c0.n12704\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__28843\,
            I => \c0.n12704\
        );

    \I__5345\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28833\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28830\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__28830\,
            I => \N__28827\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__28827\,
            I => \c0.n18082\
        );

    \I__5341\ : InMux
    port map (
            O => \N__28824\,
            I => \N__28821\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__28821\,
            I => \c0.n18270\
        );

    \I__5339\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28805\
        );

    \I__5338\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28805\
        );

    \I__5337\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28805\
        );

    \I__5336\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28805\
        );

    \I__5335\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28800\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__28805\,
            I => \N__28797\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__28804\,
            I => \N__28794\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__28803\,
            I => \N__28788\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__28800\,
            I => \N__28784\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__28797\,
            I => \N__28781\
        );

    \I__5329\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28778\
        );

    \I__5328\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28767\
        );

    \I__5327\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28767\
        );

    \I__5326\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28767\
        );

    \I__5325\ : InMux
    port map (
            O => \N__28788\,
            I => \N__28767\
        );

    \I__5324\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28767\
        );

    \I__5323\ : Odrv12
    port map (
            O => \N__28784\,
            I => \c0.n6035\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__28781\,
            I => \c0.n6035\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__28778\,
            I => \c0.n6035\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__28767\,
            I => \c0.n6035\
        );

    \I__5319\ : InMux
    port map (
            O => \N__28758\,
            I => \bfn_9_6_0_\
        );

    \I__5318\ : InMux
    port map (
            O => \N__28755\,
            I => \c0.tx2.n16539\
        );

    \I__5317\ : InMux
    port map (
            O => \N__28752\,
            I => \c0.tx2.n16540\
        );

    \I__5316\ : InMux
    port map (
            O => \N__28749\,
            I => \c0.tx2.n16541\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__28746\,
            I => \c0.n18284_cascade_\
        );

    \I__5314\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__28737\,
            I => \c0.n27_adj_2405\
        );

    \I__5311\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28731\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__28728\,
            I => \N__28725\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__28725\,
            I => \c0.n29_adj_2408\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__28722\,
            I => \c0.n12704_cascade_\
        );

    \I__5306\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28716\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__28716\,
            I => \c0.n18287\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__28713\,
            I => \N__28709\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__28712\,
            I => \N__28706\
        );

    \I__5302\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28703\
        );

    \I__5301\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28700\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__28703\,
            I => \N__28693\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28690\
        );

    \I__5298\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28681\
        );

    \I__5297\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28681\
        );

    \I__5296\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28681\
        );

    \I__5295\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28681\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__28693\,
            I => \N__28678\
        );

    \I__5293\ : Span4Mux_v
    port map (
            O => \N__28690\,
            I => \N__28675\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__28681\,
            I => \N__28672\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__28678\,
            I => \N__28669\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__28675\,
            I => \N__28664\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__28672\,
            I => \N__28664\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__28669\,
            I => n612
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__28664\,
            I => n612
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__28659\,
            I => \c0.n18289_cascade_\
        );

    \I__5285\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28651\
        );

    \I__5284\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28646\
        );

    \I__5283\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28646\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__28651\,
            I => \c0.n18831\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__28646\,
            I => \c0.n18831\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__28641\,
            I => \c0.n18079_cascade_\
        );

    \I__5279\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28635\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__28635\,
            I => \N__28632\
        );

    \I__5277\ : Odrv12
    port map (
            O => \N__28632\,
            I => \c0.n17725\
        );

    \I__5276\ : InMux
    port map (
            O => \N__28629\,
            I => \N__28626\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__28626\,
            I => \N__28623\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__28623\,
            I => \N__28620\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__28620\,
            I => \c0.n16863\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__5271\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__28608\,
            I => \c0.n16982\
        );

    \I__5268\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__28596\,
            I => \c0.n17722\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__5263\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__28587\,
            I => \c0.n28_adj_2403\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__28584\,
            I => \n17689_cascade_\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__28578\,
            I => \c0.n18684\
        );

    \I__5258\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28569\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__28569\,
            I => \c0.n18072\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__28566\,
            I => \c0.tx2.n14_cascade_\
        );

    \I__5254\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__28560\,
            I => \c0.n18843\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__28557\,
            I => \c0.n18846_cascade_\
        );

    \I__5251\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__28551\,
            I => \c0.n22_adj_2239\
        );

    \I__5249\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28545\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__28533\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__28530\,
            I => \c0.n18675_cascade_\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__28527\,
            I => \c0.n18678_cascade_\
        );

    \I__5241\ : CascadeMux
    port map (
            O => \N__28524\,
            I => \c0.n18741_cascade_\
        );

    \I__5240\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__28518\,
            I => \c0.n22_adj_2242\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__28515\,
            I => \c0.n18744_cascade_\
        );

    \I__5237\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28509\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__5234\ : Span4Mux_h
    port map (
            O => \N__28503\,
            I => \N__28500\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__28500\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__5232\ : InMux
    port map (
            O => \N__28497\,
            I => \bfn_7_16_0_\
        );

    \I__5231\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28490\
        );

    \I__5230\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28487\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28484\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28487\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__28484\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__5226\ : SRMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__28476\,
            I => \N__28472\
        );

    \I__5224\ : SRMux
    port map (
            O => \N__28475\,
            I => \N__28469\
        );

    \I__5223\ : Sp12to4
    port map (
            O => \N__28472\,
            I => \N__28464\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28464\
        );

    \I__5221\ : Odrv12
    port map (
            O => \N__28464\,
            I => \c0.tx.n11297\
        );

    \I__5220\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28457\
        );

    \I__5219\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28454\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__28457\,
            I => \control.n8\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__28454\,
            I => \control.n8\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__28449\,
            I => \control.PHASES_5_N_2152_1_cascade_\
        );

    \I__5215\ : SRMux
    port map (
            O => \N__28446\,
            I => \N__28443\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__28443\,
            I => \control.n10356\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__28440\,
            I => \c0.n18801_cascade_\
        );

    \I__5212\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__28434\,
            I => \c0.n18804\
        );

    \I__5210\ : InMux
    port map (
            O => \N__28431\,
            I => \N__28428\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__28428\,
            I => \c0.tx.n54\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__28425\,
            I => \c0.tx.n47_cascade_\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__28422\,
            I => \N__28418\
        );

    \I__5206\ : InMux
    port map (
            O => \N__28421\,
            I => \N__28414\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28409\
        );

    \I__5204\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28409\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__28414\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__28409\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__5201\ : InMux
    port map (
            O => \N__28404\,
            I => \bfn_7_15_0_\
        );

    \I__5200\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28397\
        );

    \I__5199\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28394\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__28397\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__28394\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__5196\ : InMux
    port map (
            O => \N__28389\,
            I => \c0.tx.n16524\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28382\
        );

    \I__5194\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__5193\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__28379\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__28376\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__5190\ : InMux
    port map (
            O => \N__28371\,
            I => \c0.tx.n16525\
        );

    \I__5189\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28363\
        );

    \I__5188\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28358\
        );

    \I__5187\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28358\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__28363\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__28358\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__5184\ : InMux
    port map (
            O => \N__28353\,
            I => \c0.tx.n16526\
        );

    \I__5183\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28346\
        );

    \I__5182\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28343\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__28346\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__28343\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__5179\ : InMux
    port map (
            O => \N__28338\,
            I => \c0.tx.n16527\
        );

    \I__5178\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28331\
        );

    \I__5177\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__28331\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__28328\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__5174\ : InMux
    port map (
            O => \N__28323\,
            I => \c0.tx.n16528\
        );

    \I__5173\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28316\
        );

    \I__5172\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28313\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__28316\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__28313\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__5169\ : InMux
    port map (
            O => \N__28308\,
            I => \c0.tx.n16529\
        );

    \I__5168\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28301\
        );

    \I__5167\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28298\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__28301\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__28298\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__5164\ : InMux
    port map (
            O => \N__28293\,
            I => \c0.tx.n16530\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__28290\,
            I => \c0.rx.n18024_cascade_\
        );

    \I__5162\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28283\
        );

    \I__5161\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28280\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28277\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__28280\,
            I => \c0.rx.n12828\
        );

    \I__5158\ : Odrv12
    port map (
            O => \N__28277\,
            I => \c0.rx.n12828\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__28272\,
            I => \c0.rx.n12828_cascade_\
        );

    \I__5156\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__28263\,
            I => \c0.rx.n18303\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__5152\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__28254\,
            I => \N__28247\
        );

    \I__5150\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28244\
        );

    \I__5149\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28239\
        );

    \I__5148\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28239\
        );

    \I__5147\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28236\
        );

    \I__5146\ : Span4Mux_h
    port map (
            O => \N__28247\,
            I => \N__28233\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__28244\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__28239\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__28236\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__28233\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__5141\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28219\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28223\,
            I => \N__28216\
        );

    \I__5139\ : InMux
    port map (
            O => \N__28222\,
            I => \N__28213\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28210\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28207\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__28213\,
            I => \c0.rx.n15902\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__28210\,
            I => \c0.rx.n15902\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__28207\,
            I => \c0.rx.n15902\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28193\
        );

    \I__5132\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28190\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28185\
        );

    \I__5130\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28185\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__28196\,
            I => \N__28182\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28179\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28174\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28174\
        );

    \I__5125\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28171\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28168\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__28174\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__28171\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__28168\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__5120\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28158\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__28158\,
            I => \c0.rx.n18211\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__28155\,
            I => \N__28151\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__28154\,
            I => \N__28145\
        );

    \I__5116\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28140\
        );

    \I__5115\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28140\
        );

    \I__5114\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28132\
        );

    \I__5113\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28127\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28127\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__28140\,
            I => \N__28124\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__28139\,
            I => \N__28120\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__28138\,
            I => \N__28114\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__28137\,
            I => \N__28111\
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__28136\,
            I => \N__28108\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__28135\,
            I => \N__28103\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__28132\,
            I => \N__28095\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28095\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__28124\,
            I => \N__28095\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28090\
        );

    \I__5101\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28090\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28087\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__28118\,
            I => \N__28083\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28077\
        );

    \I__5097\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28077\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28070\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28070\
        );

    \I__5094\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28070\
        );

    \I__5093\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28063\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28063\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28063\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__28095\,
            I => \N__28056\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28056\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__28087\,
            I => \N__28056\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28053\
        );

    \I__5086\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28050\
        );

    \I__5085\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28047\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28042\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__28070\,
            I => \N__28042\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28037\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__28056\,
            I => \N__28037\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28034\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__28050\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__28047\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__5077\ : Odrv12
    port map (
            O => \N__28042\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__28037\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__28034\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__5074\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28015\
        );

    \I__5073\ : InMux
    port map (
            O => \N__28022\,
            I => \N__28015\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28021\,
            I => \N__28012\
        );

    \I__5071\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28007\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__28000\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__28012\,
            I => \N__28000\
        );

    \I__5068\ : InMux
    port map (
            O => \N__28011\,
            I => \N__27994\
        );

    \I__5067\ : InMux
    port map (
            O => \N__28010\,
            I => \N__27994\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__27990\
        );

    \I__5065\ : InMux
    port map (
            O => \N__28006\,
            I => \N__27985\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27985\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__28000\,
            I => \N__27982\
        );

    \I__5062\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27978\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27975\
        );

    \I__5060\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27972\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27965\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27965\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__27982\,
            I => \N__27965\
        );

    \I__5056\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27962\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__27978\,
            I => \N__27959\
        );

    \I__5054\ : Odrv12
    port map (
            O => \N__27975\,
            I => \r_Rx_Data\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__27972\,
            I => \r_Rx_Data\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__27965\,
            I => \r_Rx_Data\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__27962\,
            I => \r_Rx_Data\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__27959\,
            I => \r_Rx_Data\
        );

    \I__5049\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27935\
        );

    \I__5048\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27930\
        );

    \I__5047\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27930\
        );

    \I__5046\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27927\
        );

    \I__5045\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27921\
        );

    \I__5044\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27921\
        );

    \I__5043\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27911\
        );

    \I__5042\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27911\
        );

    \I__5041\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27911\
        );

    \I__5040\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27911\
        );

    \I__5039\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27908\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__27935\,
            I => \N__27901\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__27930\,
            I => \N__27901\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__27927\,
            I => \N__27901\
        );

    \I__5035\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27898\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__27921\,
            I => \N__27895\
        );

    \I__5033\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27892\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27889\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__27908\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5030\ : Odrv12
    port map (
            O => \N__27901\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__27898\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__27895\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__27892\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5026\ : Odrv12
    port map (
            O => \N__27889\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__5025\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27873\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__27873\,
            I => \c0.rx.n4\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__27870\,
            I => \c0.tx.n54_cascade_\
        );

    \I__5022\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27861\
        );

    \I__5021\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27861\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__27861\,
            I => \c0.tx.n10\
        );

    \I__5019\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27850\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \N__27847\
        );

    \I__5017\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27842\
        );

    \I__5016\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27837\
        );

    \I__5015\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27837\
        );

    \I__5014\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27834\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27831\
        );

    \I__5012\ : InMux
    port map (
            O => \N__27847\,
            I => \N__27828\
        );

    \I__5011\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27823\
        );

    \I__5010\ : InMux
    port map (
            O => \N__27845\,
            I => \N__27823\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__27842\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__27837\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__27834\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__27831\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__27828\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__27823\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__5003\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27804\
        );

    \I__5002\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27801\
        );

    \I__5001\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27798\
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__27807\,
            I => \N__27793\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__27804\,
            I => \N__27790\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__27801\,
            I => \N__27785\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__27798\,
            I => \N__27785\
        );

    \I__4996\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27782\
        );

    \I__4995\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27779\
        );

    \I__4994\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27776\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__27790\,
            I => \N__27773\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__27785\,
            I => \N__27770\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__27782\,
            I => \N__27763\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27763\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__27776\,
            I => \N__27763\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__27773\,
            I => \N__27758\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__27770\,
            I => \N__27758\
        );

    \I__4986\ : Odrv12
    port map (
            O => \N__27763\,
            I => \c0.rx.n167\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__27758\,
            I => \c0.rx.n167\
        );

    \I__4984\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27749\
        );

    \I__4983\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27745\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27742\
        );

    \I__4981\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27739\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27736\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__27742\,
            I => n12527
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__27739\,
            I => n12527
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__27736\,
            I => n12527
        );

    \I__4976\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27722\
        );

    \I__4975\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27722\
        );

    \I__4974\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27719\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__27722\,
            I => data_in_0_0
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__27719\,
            I => data_in_0_0
        );

    \I__4971\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27704\
        );

    \I__4970\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27704\
        );

    \I__4969\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27704\
        );

    \I__4968\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27701\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__27704\,
            I => data_in_3_7
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__27701\,
            I => data_in_3_7
        );

    \I__4965\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__27693\,
            I => \c0.n6_adj_2368\
        );

    \I__4963\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27685\
        );

    \I__4962\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27680\
        );

    \I__4961\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27680\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__27685\,
            I => data_in_1_3
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__27680\,
            I => data_in_1_3
        );

    \I__4958\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27670\
        );

    \I__4957\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27665\
        );

    \I__4956\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27665\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__27670\,
            I => data_in_0_3
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__27665\,
            I => data_in_0_3
        );

    \I__4953\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27655\
        );

    \I__4952\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27650\
        );

    \I__4951\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27650\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__27655\,
            I => data_in_0_1
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__27650\,
            I => data_in_0_1
        );

    \I__4948\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__27642\,
            I => \c0.rx.n18196\
        );

    \I__4946\ : InMux
    port map (
            O => \N__27639\,
            I => \N__27636\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27633\
        );

    \I__4944\ : Odrv12
    port map (
            O => \N__27633\,
            I => \c0.rx.n18194\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__27630\,
            I => \c0.rx.n12552_cascade_\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__27627\,
            I => \N__27624\
        );

    \I__4941\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27617\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27614\
        );

    \I__4939\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27611\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27608\
        );

    \I__4937\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27605\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27599\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27599\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__27611\,
            I => \N__27596\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27591\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27591\
        );

    \I__4931\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27588\
        );

    \I__4930\ : Span4Mux_v
    port map (
            O => \N__27599\,
            I => \N__27579\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__27596\,
            I => \N__27579\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__27591\,
            I => \N__27579\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27576\
        );

    \I__4926\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27573\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__27586\,
            I => \N__27569\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__27579\,
            I => \N__27566\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__27576\,
            I => \N__27561\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__27573\,
            I => \N__27561\
        );

    \I__4921\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27556\
        );

    \I__4920\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27556\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__27566\,
            I => rx_data_6
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__27561\,
            I => rx_data_6
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__27556\,
            I => rx_data_6
        );

    \I__4916\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27544\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__27548\,
            I => \N__27536\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__27547\,
            I => \N__27533\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27530\
        );

    \I__4912\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27523\
        );

    \I__4911\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27523\
        );

    \I__4910\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27520\
        );

    \I__4909\ : CascadeMux
    port map (
            O => \N__27540\,
            I => \N__27517\
        );

    \I__4908\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27514\
        );

    \I__4907\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27511\
        );

    \I__4906\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27507\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__27530\,
            I => \N__27504\
        );

    \I__4904\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27501\
        );

    \I__4903\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27498\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__27523\,
            I => \N__27493\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27493\
        );

    \I__4900\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27490\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27487\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27484\
        );

    \I__4897\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27481\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__27507\,
            I => \N__27474\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__27504\,
            I => \N__27474\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__27501\,
            I => \N__27474\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__27498\,
            I => \N__27469\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__27493\,
            I => \N__27469\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__27490\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4890\ : Odrv12
    port map (
            O => \N__27487\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__27484\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__27481\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__27474\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__27469\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__4885\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27452\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27444\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__27452\,
            I => \N__27441\
        );

    \I__4882\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27436\
        );

    \I__4881\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27436\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__27449\,
            I => \N__27431\
        );

    \I__4879\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27423\
        );

    \I__4878\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27423\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27416\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__27441\,
            I => \N__27416\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27416\
        );

    \I__4874\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27411\
        );

    \I__4873\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27411\
        );

    \I__4872\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27405\
        );

    \I__4871\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27405\
        );

    \I__4870\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27402\
        );

    \I__4869\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27399\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27396\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__27416\,
            I => \N__27391\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27391\
        );

    \I__4865\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27388\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__27405\,
            I => \N__27385\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__27402\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__27399\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4861\ : Odrv12
    port map (
            O => \N__27396\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__27391\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__27388\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4858\ : Odrv12
    port map (
            O => \N__27385\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__4857\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27366\
        );

    \I__4856\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27366\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__27357\,
            I => n164_adj_2464
        );

    \I__4851\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27349\
        );

    \I__4850\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27346\
        );

    \I__4849\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27343\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__27349\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__27346\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__27343\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__4845\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27331\
        );

    \I__4844\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27328\
        );

    \I__4843\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27325\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__27331\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__27328\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__27325\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__27318\,
            I => \N__27313\
        );

    \I__4838\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27310\
        );

    \I__4837\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27307\
        );

    \I__4836\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27304\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__27310\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__27307\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27304\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__27297\,
            I => \c0.rx.n17990_cascade_\
        );

    \I__4831\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27289\
        );

    \I__4830\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27286\
        );

    \I__4829\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27283\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__27289\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__27286\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__27283\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__4825\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27271\
        );

    \I__4824\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27268\
        );

    \I__4823\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27265\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__27271\,
            I => data_in_2_6
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__27268\,
            I => data_in_2_6
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__27265\,
            I => data_in_2_6
        );

    \I__4819\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__27255\,
            I => \N__27249\
        );

    \I__4817\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27246\
        );

    \I__4816\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27241\
        );

    \I__4815\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27241\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__27249\,
            I => data_in_1_6
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__27246\,
            I => data_in_1_6
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__27241\,
            I => data_in_1_6
        );

    \I__4811\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__4808\ : Span4Mux_h
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__27222\,
            I => \c0.rx.n18304\
        );

    \I__4806\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27213\
        );

    \I__4805\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27206\
        );

    \I__4804\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27206\
        );

    \I__4803\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27202\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27199\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27194\
        );

    \I__4800\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27194\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27191\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__27205\,
            I => \N__27188\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27202\,
            I => \N__27184\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__27199\,
            I => \N__27181\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__27194\,
            I => \N__27178\
        );

    \I__4794\ : Span4Mux_h
    port map (
            O => \N__27191\,
            I => \N__27175\
        );

    \I__4793\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27172\
        );

    \I__4792\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27169\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__27184\,
            I => rx_data_5
        );

    \I__4790\ : Odrv4
    port map (
            O => \N__27181\,
            I => rx_data_5
        );

    \I__4789\ : Odrv12
    port map (
            O => \N__27178\,
            I => rx_data_5
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__27175\,
            I => rx_data_5
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__27172\,
            I => rx_data_5
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27169\,
            I => rx_data_5
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__27156\,
            I => \N__27152\
        );

    \I__4784\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27145\
        );

    \I__4783\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27145\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27140\
        );

    \I__4781\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27140\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__27145\,
            I => data_in_3_5
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__27140\,
            I => data_in_3_5
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27131\
        );

    \I__4777\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27128\
        );

    \I__4776\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27125\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27128\,
            I => \N__27122\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__27125\,
            I => \N__27116\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__27122\,
            I => \N__27116\
        );

    \I__4772\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27113\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__27116\,
            I => \N__27107\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__27113\,
            I => \N__27103\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27100\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27097\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__27110\,
            I => \N__27093\
        );

    \I__4766\ : Span4Mux_h
    port map (
            O => \N__27107\,
            I => \N__27090\
        );

    \I__4765\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27087\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__27103\,
            I => \N__27080\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27080\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__27097\,
            I => \N__27080\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27075\
        );

    \I__4760\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27075\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__27090\,
            I => rx_data_1
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__27087\,
            I => rx_data_1
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__27080\,
            I => rx_data_1
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__27075\,
            I => rx_data_1
        );

    \I__4755\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27063\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__27063\,
            I => \N__27057\
        );

    \I__4753\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27054\
        );

    \I__4752\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27051\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27060\,
            I => \N__27048\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__27057\,
            I => data_in_3_0
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__27054\,
            I => data_in_3_0
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__27051\,
            I => data_in_3_0
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__27048\,
            I => data_in_3_0
        );

    \I__4746\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27036\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27032\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__27035\,
            I => \N__27027\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__27032\,
            I => \N__27024\
        );

    \I__4742\ : InMux
    port map (
            O => \N__27031\,
            I => \N__27021\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27016\
        );

    \I__4740\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27016\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__27024\,
            I => data_in_2_0
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__27021\,
            I => data_in_2_0
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__27016\,
            I => data_in_2_0
        );

    \I__4736\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27005\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__27008\,
            I => \N__27002\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__27005\,
            I => \N__26997\
        );

    \I__4733\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26992\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26992\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26989\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__26997\,
            I => data_in_1_7
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__26992\,
            I => data_in_1_7
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__26989\,
            I => data_in_1_7
        );

    \I__4727\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__26979\,
            I => \c0.n13693\
        );

    \I__4725\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26971\
        );

    \I__4724\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26968\
        );

    \I__4723\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26964\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__26971\,
            I => \N__26959\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__26968\,
            I => \N__26959\
        );

    \I__4720\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26951\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26946\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__26959\,
            I => \N__26946\
        );

    \I__4717\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26943\
        );

    \I__4716\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26938\
        );

    \I__4715\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26938\
        );

    \I__4714\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26933\
        );

    \I__4713\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26933\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__26951\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__26946\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__26943\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__26938\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__26933\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__26922\,
            I => \c0.rx.n11041_cascade_\
        );

    \I__4706\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__26913\,
            I => \c0.n8_adj_2385\
        );

    \I__4703\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__26907\,
            I => \c0.n15_adj_2372\
        );

    \I__4701\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26896\
        );

    \I__4700\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26896\
        );

    \I__4699\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26891\
        );

    \I__4698\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26891\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__26896\,
            I => data_in_1_2
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__26891\,
            I => data_in_1_2
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \N__26882\
        );

    \I__4694\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26879\
        );

    \I__4693\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26876\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__26879\,
            I => data_in_0_7
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__26876\,
            I => data_in_0_7
        );

    \I__4690\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26867\
        );

    \I__4689\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26860\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__26867\,
            I => \N__26857\
        );

    \I__4687\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26852\
        );

    \I__4686\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26852\
        );

    \I__4685\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26848\
        );

    \I__4684\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26845\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26842\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__26857\,
            I => \N__26837\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26837\
        );

    \I__4680\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26834\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__26848\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__26845\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__26842\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__26837\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__26834\,
            I => \c0.rx.r_Bit_Index_0\
        );

    \I__4674\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__4672\ : Span12Mux_s9_v
    port map (
            O => \N__26817\,
            I => \N__26814\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__26814\,
            I => n151
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__26811\,
            I => \n151_cascade_\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__26808\,
            I => \N__26804\
        );

    \I__4668\ : InMux
    port map (
            O => \N__26807\,
            I => \N__26799\
        );

    \I__4667\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26796\
        );

    \I__4666\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26793\
        );

    \I__4665\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26790\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26783\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26783\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__26793\,
            I => \N__26783\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__26790\,
            I => data_in_2_2
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__26783\,
            I => data_in_2_2
        );

    \I__4659\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__26775\,
            I => \c0.n18008\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__26772\,
            I => \c0.n8_adj_2369_cascade_\
        );

    \I__4656\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26765\
        );

    \I__4655\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26762\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__26765\,
            I => \c0.n10493\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__26762\,
            I => \c0.n10493\
        );

    \I__4652\ : InMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__26751\,
            I => \N__26746\
        );

    \I__4649\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26743\
        );

    \I__4648\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26740\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__26746\,
            I => data_in_1_0
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__26743\,
            I => data_in_1_0
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__26740\,
            I => data_in_1_0
        );

    \I__4644\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__26730\,
            I => \c0.rx.n110\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__26727\,
            I => \N__26722\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__26726\,
            I => \N__26719\
        );

    \I__4640\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26715\
        );

    \I__4639\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26712\
        );

    \I__4638\ : InMux
    port map (
            O => \N__26719\,
            I => \N__26709\
        );

    \I__4637\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26706\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__26715\,
            I => \N__26700\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26693\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26693\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__26706\,
            I => \N__26693\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26690\
        );

    \I__4631\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26684\
        );

    \I__4630\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26684\
        );

    \I__4629\ : Sp12to4
    port map (
            O => \N__26700\,
            I => \N__26681\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__26693\,
            I => \N__26676\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__26690\,
            I => \N__26676\
        );

    \I__4626\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26673\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__26684\,
            I => rx_data_2
        );

    \I__4624\ : Odrv12
    port map (
            O => \N__26681\,
            I => rx_data_2
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__26676\,
            I => rx_data_2
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__26673\,
            I => rx_data_2
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__26664\,
            I => \c0.rx.r_SM_Main_2_N_2088_2_cascade_\
        );

    \I__4620\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26656\
        );

    \I__4619\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26651\
        );

    \I__4618\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26651\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__26656\,
            I => \c0.rx.n161\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__26651\,
            I => \c0.rx.n161\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__4614\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26639\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__26642\,
            I => \N__26634\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26630\
        );

    \I__4611\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26625\
        );

    \I__4610\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26621\
        );

    \I__4609\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26616\
        );

    \I__4608\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26616\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__26630\,
            I => \N__26613\
        );

    \I__4606\ : InMux
    port map (
            O => \N__26629\,
            I => \N__26610\
        );

    \I__4605\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26607\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26604\
        );

    \I__4603\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26601\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__26621\,
            I => \N__26598\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__26616\,
            I => \N__26595\
        );

    \I__4600\ : Sp12to4
    port map (
            O => \N__26613\,
            I => \N__26592\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26585\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__26607\,
            I => \N__26585\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__26604\,
            I => \N__26585\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__26601\,
            I => rx_data_0
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__26598\,
            I => rx_data_0
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__26595\,
            I => rx_data_0
        );

    \I__4593\ : Odrv12
    port map (
            O => \N__26592\,
            I => rx_data_0
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__26585\,
            I => rx_data_0
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__26574\,
            I => \N__26568\
        );

    \I__4590\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26563\
        );

    \I__4589\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26563\
        );

    \I__4588\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26560\
        );

    \I__4587\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26557\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__26563\,
            I => data_in_3_2
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26560\,
            I => data_in_3_2
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__26557\,
            I => data_in_3_2
        );

    \I__4583\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26546\
        );

    \I__4582\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26542\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__26546\,
            I => \N__26539\
        );

    \I__4580\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26536\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__26542\,
            I => data_in_0_6
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__26539\,
            I => data_in_0_6
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__26536\,
            I => data_in_0_6
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__26529\,
            I => \N__26524\
        );

    \I__4575\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26520\
        );

    \I__4574\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26515\
        );

    \I__4573\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26515\
        );

    \I__4572\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26512\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__26520\,
            I => data_in_3_6
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__26515\,
            I => data_in_3_6
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__26512\,
            I => data_in_3_6
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__4567\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26497\
        );

    \I__4566\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26491\
        );

    \I__4565\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26488\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__26497\,
            I => \N__26485\
        );

    \I__4563\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26482\
        );

    \I__4562\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26479\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__26494\,
            I => \N__26476\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__26491\,
            I => \N__26471\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__26488\,
            I => \N__26468\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__26485\,
            I => \N__26465\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26460\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__26479\,
            I => \N__26460\
        );

    \I__4555\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26455\
        );

    \I__4554\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26455\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__26474\,
            I => \N__26452\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__26471\,
            I => \N__26449\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__26468\,
            I => \N__26446\
        );

    \I__4550\ : Sp12to4
    port map (
            O => \N__26465\,
            I => \N__26439\
        );

    \I__4549\ : Span12Mux_v
    port map (
            O => \N__26460\,
            I => \N__26439\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__26455\,
            I => \N__26439\
        );

    \I__4547\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26436\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__26449\,
            I => rx_data_4
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__26446\,
            I => rx_data_4
        );

    \I__4544\ : Odrv12
    port map (
            O => \N__26439\,
            I => rx_data_4
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__26436\,
            I => rx_data_4
        );

    \I__4542\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26416\
        );

    \I__4541\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26416\
        );

    \I__4540\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26413\
        );

    \I__4539\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26410\
        );

    \I__4538\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26403\
        );

    \I__4537\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26403\
        );

    \I__4536\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26403\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__26416\,
            I => n120
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__26413\,
            I => n120
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__26410\,
            I => n120
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__26403\,
            I => n120
        );

    \I__4531\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26390\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__26393\,
            I => \N__26386\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26383\
        );

    \I__4528\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26378\
        );

    \I__4527\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26378\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__26383\,
            I => data_in_frame_2_4
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__26378\,
            I => data_in_frame_2_4
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \c0.rx.n18729_cascade_\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \c0.rx.n18732_cascade_\
        );

    \I__4522\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26364\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26361\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__26361\,
            I => \c0.rx.n11\
        );

    \I__4519\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__26355\,
            I => \N__26351\
        );

    \I__4517\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26348\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__26351\,
            I => n12582
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__26348\,
            I => n12582
        );

    \I__4514\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26340\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26336\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26333\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__26336\,
            I => \N__26328\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__26333\,
            I => \N__26328\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__26328\,
            I => n135_adj_2463
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__26325\,
            I => \n4_adj_2471_cascade_\
        );

    \I__4507\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26318\
        );

    \I__4506\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26315\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__26318\,
            I => \N__26312\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__26315\,
            I => data_in_frame_5_5
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__26312\,
            I => data_in_frame_5_5
        );

    \I__4502\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26304\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__26304\,
            I => \N__26299\
        );

    \I__4500\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26294\
        );

    \I__4499\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26291\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__26299\,
            I => \N__26288\
        );

    \I__4497\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26285\
        );

    \I__4496\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26282\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__26294\,
            I => \c0.data_in_frame_1_3\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__26291\,
            I => \c0.data_in_frame_1_3\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__26288\,
            I => \c0.data_in_frame_1_3\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__26285\,
            I => \c0.data_in_frame_1_3\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__26282\,
            I => \c0.data_in_frame_1_3\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__26271\,
            I => \c0.n16981_cascade_\
        );

    \I__4489\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26265\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__26265\,
            I => \c0.n20_adj_2397\
        );

    \I__4487\ : InMux
    port map (
            O => \N__26262\,
            I => \N__26259\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__26259\,
            I => \N__26256\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__26256\,
            I => \N__26253\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__26250\,
            I => \c0.n20_adj_2350\
        );

    \I__4482\ : InMux
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__26244\,
            I => \c0.n2128\
        );

    \I__4480\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26237\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26234\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__26234\,
            I => data_in_frame_6_4
        );

    \I__4476\ : Odrv4
    port map (
            O => \N__26231\,
            I => data_in_frame_6_4
        );

    \I__4475\ : InMux
    port map (
            O => \N__26226\,
            I => \N__26223\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__26223\,
            I => \N__26219\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26216\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__26219\,
            I => \N__26213\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__26216\,
            I => data_in_frame_5_0
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__26213\,
            I => data_in_frame_5_0
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__26208\,
            I => \c0.n2128_cascade_\
        );

    \I__4468\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26202\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__26202\,
            I => \N__26199\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__26199\,
            I => \c0.n22_adj_2392\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__26193\,
            I => \N__26188\
        );

    \I__4463\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26185\
        );

    \I__4462\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26182\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__26188\,
            I => data_in_frame_0_2
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__26185\,
            I => data_in_frame_0_2
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__26182\,
            I => data_in_frame_0_2
        );

    \I__4458\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26171\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__26174\,
            I => \N__26167\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26164\
        );

    \I__4455\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26160\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26157\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__26164\,
            I => \N__26154\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26151\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__26160\,
            I => data_in_frame_0_3
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__26157\,
            I => data_in_frame_0_3
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__26154\,
            I => data_in_frame_0_3
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__26151\,
            I => data_in_frame_0_3
        );

    \I__4447\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26136\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26136\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__26136\,
            I => \c0.n2120\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26128\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26125\
        );

    \I__4442\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26122\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__26128\,
            I => \N__26119\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__26125\,
            I => \c0.n2124\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__26122\,
            I => \c0.n2124\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__26119\,
            I => \c0.n2124\
        );

    \I__4437\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26108\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26102\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__26105\,
            I => \c0.data_in_frame_3_4\
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__26102\,
            I => \c0.data_in_frame_3_4\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__26097\,
            I => \c0.n2120_cascade_\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26094\,
            I => \N__26090\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__26084\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__26087\,
            I => \c0.data_in_frame_3_6\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__26084\,
            I => \c0.data_in_frame_3_6\
        );

    \I__4426\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__26073\,
            I => \c0.n19_adj_2415\
        );

    \I__4423\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26063\
        );

    \I__4422\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26060\
        );

    \I__4421\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26057\
        );

    \I__4420\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26052\
        );

    \I__4419\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26052\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__26063\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__26060\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__26057\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__26052\,
            I => \c0.data_in_frame_1_0\
        );

    \I__4414\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26039\
        );

    \I__4413\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26033\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__26039\,
            I => \N__26030\
        );

    \I__4411\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26025\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26037\,
            I => \N__26025\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26022\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__26033\,
            I => \c0.data_in_frame_1_1\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__26030\,
            I => \c0.data_in_frame_1_1\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__26025\,
            I => \c0.data_in_frame_1_1\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__26022\,
            I => \c0.data_in_frame_1_1\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26009\
        );

    \I__4403\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26005\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__25999\
        );

    \I__4401\ : InMux
    port map (
            O => \N__26008\,
            I => \N__25995\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__26005\,
            I => \N__25991\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25986\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25986\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25983\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__25999\,
            I => \N__25980\
        );

    \I__4395\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25977\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__25995\,
            I => \N__25974\
        );

    \I__4393\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25971\
        );

    \I__4392\ : Span4Mux_v
    port map (
            O => \N__25991\,
            I => \N__25966\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__25986\,
            I => \N__25966\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__25983\,
            I => data_in_frame_0_7
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__25980\,
            I => data_in_frame_0_7
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__25977\,
            I => data_in_frame_0_7
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__25974\,
            I => data_in_frame_0_7
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__25971\,
            I => data_in_frame_0_7
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__25966\,
            I => data_in_frame_0_7
        );

    \I__4384\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25949\
        );

    \I__4383\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25946\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25941\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__25946\,
            I => \N__25937\
        );

    \I__4380\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25932\
        );

    \I__4379\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25932\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__25941\,
            I => \N__25929\
        );

    \I__4377\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25926\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__25937\,
            I => \c0.data_in_frame_1_4\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__25932\,
            I => \c0.data_in_frame_1_4\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__25929\,
            I => \c0.data_in_frame_1_4\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__25926\,
            I => \c0.data_in_frame_1_4\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__25917\,
            I => \c0.n17721_cascade_\
        );

    \I__4371\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25910\
        );

    \I__4370\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25906\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__25910\,
            I => \N__25903\
        );

    \I__4368\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25897\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__25906\,
            I => \N__25894\
        );

    \I__4366\ : Span4Mux_h
    port map (
            O => \N__25903\,
            I => \N__25891\
        );

    \I__4365\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25888\
        );

    \I__4364\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25883\
        );

    \I__4363\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25883\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__25897\,
            I => data_in_frame_0_6
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__25894\,
            I => data_in_frame_0_6
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__25891\,
            I => data_in_frame_0_6
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__25888\,
            I => data_in_frame_0_6
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__25883\,
            I => data_in_frame_0_6
        );

    \I__4357\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25869\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__25869\,
            I => \c0.n10_adj_2390\
        );

    \I__4355\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25855\
        );

    \I__4354\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25855\
        );

    \I__4353\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25852\
        );

    \I__4352\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25849\
        );

    \I__4351\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25846\
        );

    \I__4350\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25841\
        );

    \I__4349\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25841\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__25855\,
            I => n16797
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__25852\,
            I => n16797
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__25849\,
            I => n16797
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__25846\,
            I => n16797
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__25841\,
            I => n16797
        );

    \I__4343\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__25827\,
            I => \N__25823\
        );

    \I__4341\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25820\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__25823\,
            I => \N__25817\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__25820\,
            I => data_in_frame_5_4
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__25817\,
            I => data_in_frame_5_4
        );

    \I__4337\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__25809\,
            I => n158
        );

    \I__4335\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__25803\,
            I => \N__25799\
        );

    \I__4333\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25796\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__25799\,
            I => \N__25793\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25790\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__25793\,
            I => n12600
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__25790\,
            I => n12600
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__25785\,
            I => \N__25776\
        );

    \I__4327\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25773\
        );

    \I__4326\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25770\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25767\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__25781\,
            I => \N__25764\
        );

    \I__4323\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25758\
        );

    \I__4322\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25758\
        );

    \I__4321\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25755\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25752\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__25770\,
            I => \N__25749\
        );

    \I__4318\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25746\
        );

    \I__4317\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25743\
        );

    \I__4316\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25740\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25737\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__25755\,
            I => \N__25734\
        );

    \I__4313\ : Sp12to4
    port map (
            O => \N__25752\,
            I => \N__25729\
        );

    \I__4312\ : Sp12to4
    port map (
            O => \N__25749\,
            I => \N__25729\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__25746\,
            I => rx_data_3
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__25743\,
            I => rx_data_3
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__25740\,
            I => rx_data_3
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__25737\,
            I => rx_data_3
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__25734\,
            I => rx_data_3
        );

    \I__4306\ : Odrv12
    port map (
            O => \N__25729\,
            I => rx_data_3
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__25716\,
            I => \N__25707\
        );

    \I__4304\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25689\
        );

    \I__4303\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25689\
        );

    \I__4302\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25689\
        );

    \I__4301\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25689\
        );

    \I__4300\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25689\
        );

    \I__4299\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25686\
        );

    \I__4298\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25679\
        );

    \I__4297\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25679\
        );

    \I__4296\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25679\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \N__25674\
        );

    \I__4294\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25663\
        );

    \I__4293\ : InMux
    port map (
            O => \N__25702\,
            I => \N__25663\
        );

    \I__4292\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25663\
        );

    \I__4291\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25660\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25652\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25652\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__25679\,
            I => \N__25652\
        );

    \I__4287\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25649\
        );

    \I__4286\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25642\
        );

    \I__4285\ : InMux
    port map (
            O => \N__25674\,
            I => \N__25642\
        );

    \I__4284\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25635\
        );

    \I__4283\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25635\
        );

    \I__4282\ : InMux
    port map (
            O => \N__25671\,
            I => \N__25635\
        );

    \I__4281\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25632\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25627\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__25660\,
            I => \N__25627\
        );

    \I__4278\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25623\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__25652\,
            I => \N__25618\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25618\
        );

    \I__4275\ : InMux
    port map (
            O => \N__25648\,
            I => \N__25615\
        );

    \I__4274\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25612\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25607\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__25635\,
            I => \N__25607\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25602\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__25627\,
            I => \N__25602\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__25626\,
            I => \N__25599\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25587\
        );

    \I__4267\ : Span4Mux_v
    port map (
            O => \N__25618\,
            I => \N__25587\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__25615\,
            I => \N__25587\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25587\
        );

    \I__4264\ : Span12Mux_h
    port map (
            O => \N__25607\,
            I => \N__25584\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__25602\,
            I => \N__25581\
        );

    \I__4262\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25578\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25571\
        );

    \I__4260\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25571\
        );

    \I__4259\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25571\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__25587\,
            I => \N__25568\
        );

    \I__4257\ : Odrv12
    port map (
            O => \N__25584\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__25581\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__25578\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__25571\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__25568\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__4252\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25540\
        );

    \I__4251\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25533\
        );

    \I__4250\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25533\
        );

    \I__4249\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25533\
        );

    \I__4248\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25528\
        );

    \I__4247\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25528\
        );

    \I__4246\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25523\
        );

    \I__4245\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25523\
        );

    \I__4244\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25516\
        );

    \I__4243\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25516\
        );

    \I__4242\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25516\
        );

    \I__4241\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25507\
        );

    \I__4240\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25507\
        );

    \I__4239\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25507\
        );

    \I__4238\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25507\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__25540\,
            I => \c0.rx.n129\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__25533\,
            I => \c0.rx.n129\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__25528\,
            I => \c0.rx.n129\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__25523\,
            I => \c0.rx.n129\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__25516\,
            I => \c0.rx.n129\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__25507\,
            I => \c0.rx.n129\
        );

    \I__4231\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25490\
        );

    \I__4230\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__25490\,
            I => \N__25484\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__25487\,
            I => data_in_frame_5_3
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__25484\,
            I => data_in_frame_5_3
        );

    \I__4226\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25472\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__25478\,
            I => \N__25469\
        );

    \I__4224\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25466\
        );

    \I__4223\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25463\
        );

    \I__4222\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25460\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__25472\,
            I => \N__25457\
        );

    \I__4220\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25454\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__25466\,
            I => \c0.data_in_frame_1_2\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__25463\,
            I => \c0.data_in_frame_1_2\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__25460\,
            I => \c0.data_in_frame_1_2\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__25457\,
            I => \c0.data_in_frame_1_2\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__25454\,
            I => \c0.data_in_frame_1_2\
        );

    \I__4214\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25439\
        );

    \I__4213\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25436\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25432\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__25436\,
            I => \N__25429\
        );

    \I__4210\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25426\
        );

    \I__4209\ : Span4Mux_h
    port map (
            O => \N__25432\,
            I => \N__25423\
        );

    \I__4208\ : Odrv12
    port map (
            O => \N__25429\,
            I => \c0.n2122\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__25426\,
            I => \c0.n2122\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__25423\,
            I => \c0.n2122\
        );

    \I__4205\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25412\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__25415\,
            I => \N__25409\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25406\
        );

    \I__4202\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25403\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__25406\,
            I => data_in_frame_6_5
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__25403\,
            I => data_in_frame_6_5
        );

    \I__4199\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__25395\,
            I => \c0.n16994\
        );

    \I__4197\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25388\
        );

    \I__4196\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25382\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__25385\,
            I => \c0.data_in_frame_3_2\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__25382\,
            I => \c0.data_in_frame_3_2\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__4191\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__25371\,
            I => \N__25367\
        );

    \I__4189\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25364\
        );

    \I__4188\ : Span4Mux_h
    port map (
            O => \N__25367\,
            I => \N__25361\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__25364\,
            I => data_in_frame_6_6
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__25361\,
            I => data_in_frame_6_6
        );

    \I__4185\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__25350\,
            I => \N__25346\
        );

    \I__4182\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25343\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__25346\,
            I => \N__25340\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__25343\,
            I => data_in_frame_5_1
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__25340\,
            I => data_in_frame_5_1
        );

    \I__4178\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25332\,
            I => \N__25328\
        );

    \I__4176\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25325\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__25325\,
            I => data_in_frame_6_2
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__25322\,
            I => data_in_frame_6_2
        );

    \I__4172\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__25314\,
            I => \c0.n18315\
        );

    \I__4170\ : InMux
    port map (
            O => \N__25311\,
            I => \c0.n16481\
        );

    \I__4169\ : InMux
    port map (
            O => \N__25308\,
            I => \c0.n16482\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__4167\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25296\
        );

    \I__4166\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25293\
        );

    \I__4165\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25288\
        );

    \I__4164\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25288\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__25296\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__25293\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__25288\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__4160\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__25275\,
            I => \c0.n18316\
        );

    \I__4157\ : InMux
    port map (
            O => \N__25272\,
            I => \c0.n16483\
        );

    \I__4156\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25264\
        );

    \I__4155\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25261\
        );

    \I__4154\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25257\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__25264\,
            I => \N__25254\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__25261\,
            I => \N__25251\
        );

    \I__4151\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25248\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__25257\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__4149\ : Odrv12
    port map (
            O => \N__25254\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__25251\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__25248\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__4146\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__25233\,
            I => \c0.n18317\
        );

    \I__4143\ : InMux
    port map (
            O => \N__25230\,
            I => \c0.n16484\
        );

    \I__4142\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25222\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__25226\,
            I => \N__25219\
        );

    \I__4140\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25215\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25212\
        );

    \I__4138\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25207\
        );

    \I__4137\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25207\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__25215\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__25212\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__25207\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__4133\ : InMux
    port map (
            O => \N__25200\,
            I => \N__25185\
        );

    \I__4132\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25185\
        );

    \I__4131\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25185\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25185\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25185\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25179\
        );

    \I__4127\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25172\
        );

    \I__4126\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25172\
        );

    \I__4125\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25172\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__25179\,
            I => \c0.tx2_transmit_N_1996\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__25172\,
            I => \c0.tx2_transmit_N_1996\
        );

    \I__4122\ : InMux
    port map (
            O => \N__25167\,
            I => \c0.n16485\
        );

    \I__4121\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__25158\,
            I => \c0.n18318\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__25155\,
            I => \c0.n18100_cascade_\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__25152\,
            I => \c0.n18103_cascade_\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__25149\,
            I => \c0.n13808_cascade_\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__25146\,
            I => \c0.n14064_cascade_\
        );

    \I__4114\ : SRMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25137\
        );

    \I__4112\ : Span4Mux_s1_v
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__25134\,
            I => \c0.n4_adj_2203\
        );

    \I__4110\ : SRMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__25128\,
            I => \c0.n4_adj_2201\
        );

    \I__4108\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25116\
        );

    \I__4107\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25116\
        );

    \I__4106\ : InMux
    port map (
            O => \N__25123\,
            I => \N__25116\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25110\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__25115\,
            I => \N__25107\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__25114\,
            I => \N__25104\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__25113\,
            I => \N__25101\
        );

    \I__4101\ : Span4Mux_h
    port map (
            O => \N__25110\,
            I => \N__25095\
        );

    \I__4100\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25086\
        );

    \I__4099\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25086\
        );

    \I__4098\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25086\
        );

    \I__4097\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25086\
        );

    \I__4096\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25081\
        );

    \I__4095\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25081\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__25095\,
            I => n17694
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__25086\,
            I => n17694
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__25081\,
            I => n17694
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__25074\,
            I => \N__25070\
        );

    \I__4090\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25062\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25062\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25062\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__25059\,
            I => \N__25049\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25046\
        );

    \I__4084\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25033\
        );

    \I__4083\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25033\
        );

    \I__4082\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25033\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25033\
        );

    \I__4080\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25033\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25033\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__25049\,
            I => \c0.n43\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25046\,
            I => \c0.n43\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__25033\,
            I => \c0.n43\
        );

    \I__4075\ : SRMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__4073\ : Span4Mux_s0_v
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__25017\,
            I => \c0.n4_adj_2199\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25014\,
            I => \bfn_7_3_0_\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__4068\ : Span4Mux_h
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__24999\,
            I => \c0.n18253\
        );

    \I__4065\ : InMux
    port map (
            O => \N__24996\,
            I => \c0.n16479\
        );

    \I__4064\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__24990\,
            I => \c0.n18314\
        );

    \I__4062\ : InMux
    port map (
            O => \N__24987\,
            I => \c0.n16480\
        );

    \I__4061\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24977\
        );

    \I__4060\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24977\
        );

    \I__4059\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24974\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__24977\,
            I => blink_counter_22
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__24974\,
            I => blink_counter_22
        );

    \I__4056\ : InMux
    port map (
            O => \N__24969\,
            I => n16630
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__24966\,
            I => \N__24962\
        );

    \I__4054\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24956\
        );

    \I__4053\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__4052\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24953\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__24956\,
            I => blink_counter_23
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__24953\,
            I => blink_counter_23
        );

    \I__4049\ : InMux
    port map (
            O => \N__24948\,
            I => n16631
        );

    \I__4048\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24938\
        );

    \I__4047\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24938\
        );

    \I__4046\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24935\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__24938\,
            I => blink_counter_24
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__24935\,
            I => blink_counter_24
        );

    \I__4043\ : InMux
    port map (
            O => \N__24930\,
            I => \bfn_6_24_0_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__24927\,
            I => n16633
        );

    \I__4041\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24920\
        );

    \I__4040\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24917\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__24920\,
            I => blink_counter_25
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__24917\,
            I => blink_counter_25
        );

    \I__4037\ : CEMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__24906\,
            I => \control.n11\
        );

    \I__4034\ : IoInMux
    port map (
            O => \N__24903\,
            I => \N__24900\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__4032\ : Span4Mux_s3_v
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__24894\,
            I => \PIN_1_c_0\
        );

    \I__4030\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24888\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__24888\,
            I => n12
        );

    \I__4028\ : InMux
    port map (
            O => \N__24885\,
            I => n16622
        );

    \I__4027\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__24879\,
            I => n11
        );

    \I__4025\ : InMux
    port map (
            O => \N__24876\,
            I => n16623
        );

    \I__4024\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__24870\,
            I => n10_adj_2467
        );

    \I__4022\ : InMux
    port map (
            O => \N__24867\,
            I => \bfn_6_23_0_\
        );

    \I__4021\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__24861\,
            I => n9
        );

    \I__4019\ : InMux
    port map (
            O => \N__24858\,
            I => n16625
        );

    \I__4018\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__24852\,
            I => n8
        );

    \I__4016\ : InMux
    port map (
            O => \N__24849\,
            I => n16626
        );

    \I__4015\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__24843\,
            I => n7_adj_2476
        );

    \I__4013\ : InMux
    port map (
            O => \N__24840\,
            I => n16627
        );

    \I__4012\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__24834\,
            I => n6
        );

    \I__4010\ : InMux
    port map (
            O => \N__24831\,
            I => n16628
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__24828\,
            I => \N__24825\
        );

    \I__4008\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24818\
        );

    \I__4007\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24818\
        );

    \I__4006\ : InMux
    port map (
            O => \N__24823\,
            I => \N__24815\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__24818\,
            I => blink_counter_21
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__24815\,
            I => blink_counter_21
        );

    \I__4003\ : InMux
    port map (
            O => \N__24810\,
            I => n16629
        );

    \I__4002\ : InMux
    port map (
            O => \N__24807\,
            I => n16613
        );

    \I__4001\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__24801\,
            I => n20
        );

    \I__3999\ : InMux
    port map (
            O => \N__24798\,
            I => n16614
        );

    \I__3998\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__24792\,
            I => n19
        );

    \I__3996\ : InMux
    port map (
            O => \N__24789\,
            I => n16615
        );

    \I__3995\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__24783\,
            I => n18_adj_2480
        );

    \I__3993\ : InMux
    port map (
            O => \N__24780\,
            I => \bfn_6_22_0_\
        );

    \I__3992\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24774\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__24774\,
            I => n17
        );

    \I__3990\ : InMux
    port map (
            O => \N__24771\,
            I => n16617
        );

    \I__3989\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24765\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__24765\,
            I => n16
        );

    \I__3987\ : InMux
    port map (
            O => \N__24762\,
            I => n16618
        );

    \I__3986\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__24756\,
            I => n15_adj_2479
        );

    \I__3984\ : InMux
    port map (
            O => \N__24753\,
            I => n16619
        );

    \I__3983\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__24747\,
            I => n14_adj_2478
        );

    \I__3981\ : InMux
    port map (
            O => \N__24744\,
            I => n16620
        );

    \I__3980\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__24738\,
            I => n13
        );

    \I__3978\ : InMux
    port map (
            O => \N__24735\,
            I => n16621
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__24732\,
            I => \c0.rx.n12_cascade_\
        );

    \I__3976\ : CEMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__24720\,
            I => \c0.rx.n11082\
        );

    \I__3972\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__3970\ : Span4Mux_v
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__24708\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_18\
        );

    \I__3968\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24700\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__24704\,
            I => \N__24696\
        );

    \I__3966\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24693\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__24700\,
            I => \N__24690\
        );

    \I__3964\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24687\
        );

    \I__3963\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24684\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24681\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__24690\,
            I => \N__24678\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24673\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24673\
        );

    \I__3958\ : Span4Mux_h
    port map (
            O => \N__24681\,
            I => \N__24670\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__24678\,
            I => \N__24665\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__24673\,
            I => \N__24665\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__24670\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__24665\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__3953\ : SRMux
    port map (
            O => \N__24660\,
            I => \N__24657\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__24657\,
            I => \N__24654\
        );

    \I__3951\ : Span4Mux_h
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__24648\,
            I => \c0.n3_adj_2305\
        );

    \I__3948\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24640\
        );

    \I__3947\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24637\
        );

    \I__3946\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24634\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24617\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24612\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24612\
        );

    \I__3942\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24609\
        );

    \I__3941\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24606\
        );

    \I__3940\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24603\
        );

    \I__3939\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24600\
        );

    \I__3938\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24596\
        );

    \I__3937\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24593\
        );

    \I__3936\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24590\
        );

    \I__3935\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24587\
        );

    \I__3934\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24582\
        );

    \I__3933\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24579\
        );

    \I__3932\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24576\
        );

    \I__3931\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24573\
        );

    \I__3930\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24570\
        );

    \I__3929\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24562\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__24617\,
            I => \N__24549\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__24612\,
            I => \N__24549\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24549\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__24606\,
            I => \N__24549\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24549\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__24600\,
            I => \N__24549\
        );

    \I__3922\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24546\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24537\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__24593\,
            I => \N__24537\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__24590\,
            I => \N__24537\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__24587\,
            I => \N__24537\
        );

    \I__3917\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24534\
        );

    \I__3916\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24530\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__24582\,
            I => \N__24519\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__24579\,
            I => \N__24519\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__24576\,
            I => \N__24519\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24519\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24519\
        );

    \I__3910\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24516\
        );

    \I__3909\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24513\
        );

    \I__3908\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24510\
        );

    \I__3907\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24507\
        );

    \I__3906\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24504\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__24562\,
            I => \N__24495\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__24549\,
            I => \N__24490\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__24546\,
            I => \N__24490\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__24537\,
            I => \N__24485\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__24534\,
            I => \N__24485\
        );

    \I__3900\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24482\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24469\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__24519\,
            I => \N__24469\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24469\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__24513\,
            I => \N__24469\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__24510\,
            I => \N__24469\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__24507\,
            I => \N__24469\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__24504\,
            I => \N__24466\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24463\
        );

    \I__3891\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24460\
        );

    \I__3890\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24457\
        );

    \I__3889\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24454\
        );

    \I__3888\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24449\
        );

    \I__3887\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24449\
        );

    \I__3886\ : Span12Mux_v
    port map (
            O => \N__24495\,
            I => \N__24443\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__24490\,
            I => \N__24438\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__24485\,
            I => \N__24438\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__24482\,
            I => \N__24435\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__24469\,
            I => \N__24428\
        );

    \I__3881\ : Span4Mux_s2_h
    port map (
            O => \N__24466\,
            I => \N__24428\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24428\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24425\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__24457\,
            I => \N__24418\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__24454\,
            I => \N__24418\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24418\
        );

    \I__3875\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24415\
        );

    \I__3874\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24410\
        );

    \I__3873\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24410\
        );

    \I__3872\ : Odrv12
    port map (
            O => \N__24443\,
            I => n1166
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__24438\,
            I => n1166
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__24435\,
            I => n1166
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__24428\,
            I => n1166
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__24425\,
            I => n1166
        );

    \I__3867\ : Odrv12
    port map (
            O => \N__24418\,
            I => n1166
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__24415\,
            I => n1166
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__24410\,
            I => n1166
        );

    \I__3864\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__24384\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_13\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__24381\,
            I => \N__24375\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__24380\,
            I => \N__24372\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24369\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24366\
        );

    \I__3856\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24363\
        );

    \I__3855\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24360\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24351\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__24366\,
            I => \N__24351\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__24363\,
            I => \N__24351\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24351\
        );

    \I__3850\ : Span4Mux_h
    port map (
            O => \N__24351\,
            I => \N__24348\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__24348\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__3848\ : SRMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__24342\,
            I => \N__24339\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__24333\,
            I => \c0.n3_adj_2317\
        );

    \I__3843\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24327\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__24327\,
            I => n26
        );

    \I__3841\ : InMux
    port map (
            O => \N__24324\,
            I => \bfn_6_21_0_\
        );

    \I__3840\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__24318\,
            I => n25
        );

    \I__3838\ : InMux
    port map (
            O => \N__24315\,
            I => n16609
        );

    \I__3837\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24309\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__24309\,
            I => n24
        );

    \I__3835\ : InMux
    port map (
            O => \N__24306\,
            I => n16610
        );

    \I__3834\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24300\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__24300\,
            I => n23
        );

    \I__3832\ : InMux
    port map (
            O => \N__24297\,
            I => n16611
        );

    \I__3831\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__24291\,
            I => n22_adj_2481
        );

    \I__3829\ : InMux
    port map (
            O => \N__24288\,
            I => n16612
        );

    \I__3828\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__24282\,
            I => n21
        );

    \I__3826\ : InMux
    port map (
            O => \N__24279\,
            I => \c0.rx.n16536\
        );

    \I__3825\ : InMux
    port map (
            O => \N__24276\,
            I => \c0.rx.n16537\
        );

    \I__3824\ : InMux
    port map (
            O => \N__24273\,
            I => \c0.rx.n16538\
        );

    \I__3823\ : SRMux
    port map (
            O => \N__24270\,
            I => \N__24267\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24264\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__24264\,
            I => \c0.rx.n12819\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__24261\,
            I => \c0.n18225_cascade_\
        );

    \I__3819\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24255\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24252\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__24252\,
            I => \N__24249\
        );

    \I__3816\ : Span4Mux_h
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__24246\,
            I => \c0.rx.n5\
        );

    \I__3814\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24237\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__3811\ : Span4Mux_h
    port map (
            O => \N__24234\,
            I => \N__24231\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__24231\,
            I => \c0.rx.n57\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__24228\,
            I => \c0.rx.n15905_cascade_\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__24225\,
            I => \c0.rx.n6_cascade_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24219\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24219\,
            I => \c0.rx.n12\
        );

    \I__3805\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24208\
        );

    \I__3804\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24208\
        );

    \I__3803\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24203\
        );

    \I__3802\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24203\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__24208\,
            I => data_in_2_7
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__24203\,
            I => data_in_2_7
        );

    \I__3799\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24192\
        );

    \I__3798\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24185\
        );

    \I__3797\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24185\
        );

    \I__3796\ : InMux
    port map (
            O => \N__24195\,
            I => \N__24185\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24192\,
            I => data_in_2_5
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__24185\,
            I => data_in_2_5
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__24180\,
            I => \N__24174\
        );

    \I__3792\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24171\
        );

    \I__3791\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24166\
        );

    \I__3790\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24166\
        );

    \I__3789\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24162\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__24171\,
            I => \N__24159\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24156\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24150\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24147\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__24159\,
            I => \N__24142\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__24156\,
            I => \N__24142\
        );

    \I__3782\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24139\
        );

    \I__3781\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24136\
        );

    \I__3780\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24133\
        );

    \I__3779\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24130\
        );

    \I__3778\ : Odrv12
    port map (
            O => \N__24147\,
            I => rx_data_7
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__24142\,
            I => rx_data_7
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__24139\,
            I => rx_data_7
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__24136\,
            I => rx_data_7
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24133\,
            I => rx_data_7
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__24130\,
            I => rx_data_7
        );

    \I__3772\ : InMux
    port map (
            O => \N__24117\,
            I => \bfn_6_13_0_\
        );

    \I__3771\ : InMux
    port map (
            O => \N__24114\,
            I => \c0.rx.n16532\
        );

    \I__3770\ : InMux
    port map (
            O => \N__24111\,
            I => \c0.rx.n16533\
        );

    \I__3769\ : InMux
    port map (
            O => \N__24108\,
            I => \c0.rx.n16534\
        );

    \I__3768\ : InMux
    port map (
            O => \N__24105\,
            I => \c0.rx.n16535\
        );

    \I__3767\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24098\
        );

    \I__3766\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24094\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__24098\,
            I => \N__24091\
        );

    \I__3764\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24088\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__24094\,
            I => data_in_1_5
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__24091\,
            I => data_in_1_5
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__24088\,
            I => data_in_1_5
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__24081\,
            I => \N__24076\
        );

    \I__3759\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24073\
        );

    \I__3758\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24070\
        );

    \I__3757\ : InMux
    port map (
            O => \N__24076\,
            I => \N__24067\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__24073\,
            I => data_in_2_4
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__24070\,
            I => data_in_2_4
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__24067\,
            I => data_in_2_4
        );

    \I__3753\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24057\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__24057\,
            I => \c0.n18_adj_2370\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24051\
        );

    \I__3750\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24048\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__24048\,
            I => \c0.n13_adj_2380\
        );

    \I__3748\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24038\
        );

    \I__3746\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24035\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__24038\,
            I => \c0.rx.n10988\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__24035\,
            I => \c0.rx.n10988\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__24030\,
            I => \c0.n18006_cascade_\
        );

    \I__3742\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__24021\,
            I => \c0.n14_adj_2375\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__24018\,
            I => \c0.n20_adj_2371_cascade_\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24012\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__24012\,
            I => \c0.n10516\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__24009\,
            I => \c0.n10516_cascade_\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24006\,
            I => \N__24003\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__24003\,
            I => \c0.n10367\
        );

    \I__3733\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23995\
        );

    \I__3732\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23990\
        );

    \I__3731\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23990\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__23995\,
            I => data_in_0_5
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__23990\,
            I => data_in_0_5
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \c0.n10367_cascade_\
        );

    \I__3727\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23979\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__23979\,
            I => \c0.n15_adj_2389\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__23976\,
            I => \N__23973\
        );

    \I__3724\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23969\
        );

    \I__3723\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23964\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23961\
        );

    \I__3721\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23956\
        );

    \I__3720\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23956\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__23964\,
            I => data_in_1_4
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__23961\,
            I => data_in_1_4
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__23956\,
            I => data_in_1_4
        );

    \I__3716\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23943\
        );

    \I__3715\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23943\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__23943\,
            I => data_in_0_4
        );

    \I__3713\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23932\
        );

    \I__3712\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23932\
        );

    \I__3711\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23927\
        );

    \I__3710\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23927\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__23932\,
            I => data_in_3_4
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__23927\,
            I => data_in_3_4
        );

    \I__3707\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__23919\,
            I => \c0.n14_adj_2388\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__23916\,
            I => \N__23902\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__23915\,
            I => \N__23898\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__23914\,
            I => \N__23894\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__23913\,
            I => \N__23890\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__23912\,
            I => \N__23887\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__23911\,
            I => \N__23882\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__23910\,
            I => \N__23878\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__23909\,
            I => \N__23872\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__23908\,
            I => \N__23868\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__23907\,
            I => \N__23864\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__23906\,
            I => \N__23860\
        );

    \I__3694\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23846\
        );

    \I__3693\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23846\
        );

    \I__3692\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23846\
        );

    \I__3691\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23835\
        );

    \I__3690\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23835\
        );

    \I__3689\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23835\
        );

    \I__3688\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23835\
        );

    \I__3687\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23835\
        );

    \I__3686\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23824\
        );

    \I__3685\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23824\
        );

    \I__3684\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23824\
        );

    \I__3683\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23824\
        );

    \I__3682\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23824\
        );

    \I__3681\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23817\
        );

    \I__3680\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23817\
        );

    \I__3679\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23817\
        );

    \I__3678\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23800\
        );

    \I__3677\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23800\
        );

    \I__3676\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23800\
        );

    \I__3675\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23800\
        );

    \I__3674\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23800\
        );

    \I__3673\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23800\
        );

    \I__3672\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23800\
        );

    \I__3671\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23800\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__23859\,
            I => \N__23797\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__23858\,
            I => \N__23794\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__23857\,
            I => \N__23791\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__23856\,
            I => \N__23787\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__23855\,
            I => \N__23784\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__23854\,
            I => \N__23781\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__23853\,
            I => \N__23778\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__23846\,
            I => \N__23775\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__23835\,
            I => \N__23772\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23767\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__23817\,
            I => \N__23767\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23764\
        );

    \I__3658\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23753\
        );

    \I__3657\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23753\
        );

    \I__3656\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23753\
        );

    \I__3655\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23753\
        );

    \I__3654\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23753\
        );

    \I__3653\ : InMux
    port map (
            O => \N__23784\,
            I => \N__23746\
        );

    \I__3652\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23746\
        );

    \I__3651\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23746\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__23775\,
            I => \N__23743\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__23772\,
            I => \N__23740\
        );

    \I__3648\ : Span12Mux_s5_h
    port map (
            O => \N__23767\,
            I => \N__23737\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__23764\,
            I => \N__23734\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__23753\,
            I => \N__23729\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__23746\,
            I => \N__23729\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__23743\,
            I => \c0.n18631\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__23740\,
            I => \c0.n18631\
        );

    \I__3642\ : Odrv12
    port map (
            O => \N__23737\,
            I => \c0.n18631\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__23734\,
            I => \c0.n18631\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__23729\,
            I => \c0.n18631\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__23718\,
            I => \c0.n18002_cascade_\
        );

    \I__3638\ : InMux
    port map (
            O => \N__23715\,
            I => \N__23709\
        );

    \I__3637\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23709\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__23709\,
            I => \c0.n10498\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__23706\,
            I => \c0.rx.n10988_cascade_\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__23703\,
            I => \c0.rx.n12624_cascade_\
        );

    \I__3633\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23694\
        );

    \I__3632\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23694\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__23694\,
            I => data_in_0_2
        );

    \I__3630\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23687\
        );

    \I__3629\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23684\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__23687\,
            I => data_in_frame_5_7
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__23684\,
            I => data_in_frame_5_7
        );

    \I__3626\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23675\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__23678\,
            I => \N__23671\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__23675\,
            I => \N__23668\
        );

    \I__3623\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23665\
        );

    \I__3622\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23662\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__23668\,
            I => \N__23659\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__23665\,
            I => data_in_frame_2_7
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__23662\,
            I => data_in_frame_2_7
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__23659\,
            I => data_in_frame_2_7
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__23652\,
            I => \c0.rx.n17702_cascade_\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__3615\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__23643\,
            I => \c0.rx.n17702\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__23640\,
            I => \c0.rx.n17704_cascade_\
        );

    \I__3612\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23630\
        );

    \I__3611\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23627\
        );

    \I__3610\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23622\
        );

    \I__3609\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23617\
        );

    \I__3608\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23617\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23614\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23611\
        );

    \I__3605\ : InMux
    port map (
            O => \N__23626\,
            I => \N__23608\
        );

    \I__3604\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23605\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__23622\,
            I => n11058
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__23617\,
            I => n11058
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__23614\,
            I => n11058
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__23611\,
            I => n11058
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__23608\,
            I => n11058
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__23605\,
            I => n11058
        );

    \I__3597\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23583\
        );

    \I__3596\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23580\
        );

    \I__3595\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23575\
        );

    \I__3594\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23575\
        );

    \I__3593\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23570\
        );

    \I__3592\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23570\
        );

    \I__3591\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23567\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__23583\,
            I => n16802
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__23580\,
            I => n16802
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__23575\,
            I => n16802
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__23570\,
            I => n16802
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__23567\,
            I => n16802
        );

    \I__3585\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23551\
        );

    \I__3584\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23548\
        );

    \I__3583\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23545\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__23551\,
            I => \c0.n10569\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__23548\,
            I => \c0.n10569\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__23545\,
            I => \c0.n10569\
        );

    \I__3579\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23534\
        );

    \I__3578\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23531\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__23531\,
            I => data_in_frame_6_3
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__23528\,
            I => data_in_frame_6_3
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__23523\,
            I => \c0.n17734_cascade_\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__23520\,
            I => \N__23516\
        );

    \I__3572\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23511\
        );

    \I__3571\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23508\
        );

    \I__3570\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23503\
        );

    \I__3569\ : InMux
    port map (
            O => \N__23514\,
            I => \N__23503\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__23511\,
            I => \c0.data_in_frame_1_7\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__23508\,
            I => \c0.data_in_frame_1_7\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__23503\,
            I => \c0.data_in_frame_1_7\
        );

    \I__3565\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__23493\,
            I => \c0.n19_adj_2400\
        );

    \I__3563\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23487\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__23487\,
            I => \c0.n18_adj_2398\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \c0.n18000_cascade_\
        );

    \I__3560\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23477\
        );

    \I__3559\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23474\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__23477\,
            I => \N__23471\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__23474\,
            I => data_in_frame_5_2
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__23471\,
            I => data_in_frame_5_2
        );

    \I__3555\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23463\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23457\
        );

    \I__3553\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23454\
        );

    \I__3552\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23450\
        );

    \I__3551\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23447\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__23457\,
            I => \N__23440\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23440\
        );

    \I__3548\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23437\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23434\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__23447\,
            I => \N__23431\
        );

    \I__3545\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23428\
        );

    \I__3544\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23424\
        );

    \I__3543\ : Span4Mux_v
    port map (
            O => \N__23440\,
            I => \N__23421\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23414\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__23434\,
            I => \N__23414\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__23431\,
            I => \N__23414\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__23428\,
            I => \N__23411\
        );

    \I__3538\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23408\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__23424\,
            I => \N__23405\
        );

    \I__3536\ : Sp12to4
    port map (
            O => \N__23421\,
            I => \N__23398\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__23414\,
            I => \N__23393\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__23411\,
            I => \N__23393\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23388\
        );

    \I__3532\ : Span4Mux_s2_h
    port map (
            O => \N__23405\,
            I => \N__23388\
        );

    \I__3531\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23381\
        );

    \I__3530\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23381\
        );

    \I__3529\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23381\
        );

    \I__3528\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23378\
        );

    \I__3527\ : Odrv12
    port map (
            O => \N__23398\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__23393\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__23388\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__23381\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__23378\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__23367\,
            I => \N__23363\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__23366\,
            I => \N__23357\
        );

    \I__3520\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23353\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__23362\,
            I => \N__23350\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__23361\,
            I => \N__23346\
        );

    \I__3517\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23343\
        );

    \I__3516\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23339\
        );

    \I__3515\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23332\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23328\
        );

    \I__3513\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23325\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N__23322\
        );

    \I__3511\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23319\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__23343\,
            I => \N__23316\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__23342\,
            I => \N__23313\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23310\
        );

    \I__3507\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23305\
        );

    \I__3506\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23305\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__23336\,
            I => \N__23302\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__23335\,
            I => \N__23299\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23296\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__23331\,
            I => \N__23291\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__23328\,
            I => \N__23285\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__23325\,
            I => \N__23285\
        );

    \I__3499\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23282\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__23319\,
            I => \N__23277\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__23316\,
            I => \N__23277\
        );

    \I__3496\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23274\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__23310\,
            I => \N__23269\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23269\
        );

    \I__3493\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23266\
        );

    \I__3492\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23263\
        );

    \I__3491\ : Span4Mux_h
    port map (
            O => \N__23296\,
            I => \N__23260\
        );

    \I__3490\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23251\
        );

    \I__3489\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23251\
        );

    \I__3488\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23251\
        );

    \I__3487\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23251\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__23285\,
            I => \N__23240\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23240\
        );

    \I__3484\ : Span4Mux_h
    port map (
            O => \N__23277\,
            I => \N__23240\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__23274\,
            I => \N__23240\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__23269\,
            I => \N__23240\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__23266\,
            I => \N__23231\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__23263\,
            I => \N__23231\
        );

    \I__3479\ : Sp12to4
    port map (
            O => \N__23260\,
            I => \N__23231\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23231\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__23240\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__3476\ : Odrv12
    port map (
            O => \N__23231\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__3475\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23223\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__23223\,
            I => \N__23217\
        );

    \I__3473\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23214\
        );

    \I__3472\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23211\
        );

    \I__3471\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23207\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__23217\,
            I => \N__23200\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23200\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23200\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23197\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23194\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__23200\,
            I => \N__23187\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__23197\,
            I => \N__23187\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__23194\,
            I => \N__23187\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__23187\,
            I => \c0.rx.n12963\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__23184\,
            I => \n120_cascade_\
        );

    \I__3460\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23174\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23171\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23168\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__23171\,
            I => data_in_frame_2_3
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__23168\,
            I => data_in_frame_2_3
        );

    \I__3454\ : InMux
    port map (
            O => \N__23163\,
            I => \N__23160\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23154\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23151\
        );

    \I__3451\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23146\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23146\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__23154\,
            I => data_in_frame_0_4
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__23151\,
            I => data_in_frame_0_4
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__23146\,
            I => data_in_frame_0_4
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__23139\,
            I => \N__23136\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23133\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23127\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23124\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23121\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23118\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__23127\,
            I => data_in_frame_0_5
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__23124\,
            I => data_in_frame_0_5
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__23121\,
            I => data_in_frame_0_5
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__23118\,
            I => data_in_frame_0_5
        );

    \I__3436\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23104\
        );

    \I__3435\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23101\
        );

    \I__3434\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23098\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__23104\,
            I => data_in_frame_2_6
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__23101\,
            I => data_in_frame_2_6
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__23098\,
            I => data_in_frame_2_6
        );

    \I__3430\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23088\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__23088\,
            I => \c0.n15_adj_2416\
        );

    \I__3428\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23079\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23076\
        );

    \I__3426\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23073\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23070\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__23079\,
            I => \c0.n2138\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__23076\,
            I => \c0.n2138\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__23073\,
            I => \c0.n2138\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__23070\,
            I => \c0.n2138\
        );

    \I__3420\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__23055\,
            I => \c0.n22_adj_2419\
        );

    \I__3417\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23048\
        );

    \I__3416\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23045\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__23048\,
            I => data_in_frame_6_7
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__23045\,
            I => data_in_frame_6_7
        );

    \I__3413\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23036\
        );

    \I__3412\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23033\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__23036\,
            I => \c0.n17813\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__23033\,
            I => \c0.n17813\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__23025\,
            I => \c0.n10761\
        );

    \I__3407\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23013\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23013\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23013\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__23013\,
            I => \N__23007\
        );

    \I__3403\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23002\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23002\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23010\,
            I => \N__22999\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__23007\,
            I => data_in_frame_0_0
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23002\,
            I => data_in_frame_0_0
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__22999\,
            I => data_in_frame_0_0
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \c0.n10761_cascade_\
        );

    \I__3396\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22986\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__22986\,
            I => \N__22982\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__22985\,
            I => \N__22978\
        );

    \I__3393\ : Span4Mux_h
    port map (
            O => \N__22982\,
            I => \N__22973\
        );

    \I__3392\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22970\
        );

    \I__3391\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22965\
        );

    \I__3390\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22965\
        );

    \I__3389\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22962\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__22973\,
            I => \c0.data_in_frame_1_5\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__22970\,
            I => \c0.data_in_frame_1_5\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__22965\,
            I => \c0.data_in_frame_1_5\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__22962\,
            I => \c0.data_in_frame_1_5\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__22953\,
            I => \c0.n17733_cascade_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22946\
        );

    \I__3382\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22943\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__22946\,
            I => data_in_frame_6_0
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__22943\,
            I => data_in_frame_6_0
        );

    \I__3379\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__22935\,
            I => \c0.n17735\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__22932\,
            I => \N__22928\
        );

    \I__3376\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22923\
        );

    \I__3375\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22919\
        );

    \I__3374\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22914\
        );

    \I__3373\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22914\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22911\
        );

    \I__3371\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22908\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__22919\,
            I => \c0.data_in_frame_1_6\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__22914\,
            I => \c0.data_in_frame_1_6\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__22911\,
            I => \c0.data_in_frame_1_6\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__22908\,
            I => \c0.data_in_frame_1_6\
        );

    \I__3366\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__22896\,
            I => \c0.n17733\
        );

    \I__3364\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__22890\,
            I => \c0.n21_adj_2421\
        );

    \I__3362\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22881\
        );

    \I__3360\ : Span4Mux_h
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__22878\,
            I => \c0.n24_adj_2418\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \c0.n23_adj_2420_cascade_\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__22872\,
            I => \n16797_cascade_\
        );

    \I__3356\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22865\
        );

    \I__3355\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22859\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__22862\,
            I => \c0.data_in_frame_3_5\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__22859\,
            I => \c0.data_in_frame_3_5\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__22854\,
            I => \c0.rx.n129_cascade_\
        );

    \I__3350\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22847\
        );

    \I__3349\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22844\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22841\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__22844\,
            I => \c0.data_in_frame_3_7\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__22841\,
            I => \c0.data_in_frame_3_7\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__22836\,
            I => \N__22832\
        );

    \I__3344\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22829\
        );

    \I__3343\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22826\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__22829\,
            I => data_in_frame_6_1
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__22826\,
            I => data_in_frame_6_1
        );

    \I__3340\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__22818\,
            I => n18043
        );

    \I__3338\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__22812\,
            I => n18044
        );

    \I__3336\ : IoInMux
    port map (
            O => \N__22809\,
            I => \N__22806\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__3334\ : Span12Mux_s8_v
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__22800\,
            I => \LED_c\
        );

    \I__3332\ : IoInMux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__3330\ : Span4Mux_s3_h
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__22788\,
            I => \PIN_3_c_2\
        );

    \I__3328\ : SRMux
    port map (
            O => \N__22785\,
            I => \N__22782\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22779\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__3325\ : Span4Mux_s1_v
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__22773\,
            I => \c0.n4_adj_2225\
        );

    \I__3323\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22766\
        );

    \I__3322\ : IoInMux
    port map (
            O => \N__22769\,
            I => \N__22763\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__22766\,
            I => \N__22760\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22757\
        );

    \I__3319\ : Span4Mux_s2_v
    port map (
            O => \N__22760\,
            I => \N__22754\
        );

    \I__3318\ : Span4Mux_s2_v
    port map (
            O => \N__22757\,
            I => \N__22751\
        );

    \I__3317\ : Span4Mux_v
    port map (
            O => \N__22754\,
            I => \N__22748\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__22751\,
            I => \N__22742\
        );

    \I__3315\ : Span4Mux_v
    port map (
            O => \N__22748\,
            I => \N__22742\
        );

    \I__3314\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22739\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__22742\,
            I => tx2_o
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__22739\,
            I => tx2_o
        );

    \I__3311\ : IoInMux
    port map (
            O => \N__22734\,
            I => \N__22731\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__3309\ : Span4Mux_s1_v
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__22725\,
            I => tx2_enable
        );

    \I__3307\ : SRMux
    port map (
            O => \N__22722\,
            I => \N__22719\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__3304\ : Span4Mux_s2_h
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__22710\,
            I => \c0.n4_adj_2216\
        );

    \I__3302\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22703\
        );

    \I__3301\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22700\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__22703\,
            I => \N__22697\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__22700\,
            I => \c0.data_in_frame_3_3\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__22697\,
            I => \c0.data_in_frame_3_3\
        );

    \I__3297\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22688\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__22691\,
            I => \N__22685\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__22688\,
            I => \N__22681\
        );

    \I__3294\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22678\
        );

    \I__3293\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22675\
        );

    \I__3292\ : Span4Mux_v
    port map (
            O => \N__22681\,
            I => \N__22672\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22669\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__22675\,
            I => data_in_frame_2_2
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__22672\,
            I => data_in_frame_2_2
        );

    \I__3288\ : Odrv12
    port map (
            O => \N__22669\,
            I => data_in_frame_2_2
        );

    \I__3287\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22659\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__22659\,
            I => \c0.n18_adj_2417\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__3284\ : InMux
    port map (
            O => \N__22653\,
            I => \N__22649\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \N__22646\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__22649\,
            I => \N__22642\
        );

    \I__3281\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22639\
        );

    \I__3280\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22636\
        );

    \I__3279\ : Span4Mux_h
    port map (
            O => \N__22642\,
            I => \N__22631\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22631\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__22636\,
            I => data_in_frame_2_1
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__22631\,
            I => data_in_frame_2_1
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__22626\,
            I => \N__22623\
        );

    \I__3274\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22620\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22614\
        );

    \I__3272\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22611\
        );

    \I__3271\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22608\
        );

    \I__3270\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22605\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__22614\,
            I => \N__22602\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22595\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__22608\,
            I => \N__22595\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__22605\,
            I => \N__22595\
        );

    \I__3265\ : Span4Mux_s0_h
    port map (
            O => \N__22602\,
            I => \N__22592\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__22595\,
            I => \N__22589\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__22592\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__22589\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__3261\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__22581\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_12\
        );

    \I__3259\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__22575\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_27\
        );

    \I__3257\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22556\
        );

    \I__3256\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22556\
        );

    \I__3255\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22547\
        );

    \I__3254\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22547\
        );

    \I__3253\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22547\
        );

    \I__3252\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22547\
        );

    \I__3251\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22544\
        );

    \I__3250\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22533\
        );

    \I__3249\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22533\
        );

    \I__3248\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22533\
        );

    \I__3247\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22533\
        );

    \I__3246\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22533\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22525\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__22547\,
            I => \N__22522\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__22544\,
            I => \N__22519\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22516\
        );

    \I__3241\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22505\
        );

    \I__3240\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22505\
        );

    \I__3239\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22505\
        );

    \I__3238\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22505\
        );

    \I__3237\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22505\
        );

    \I__3236\ : Span4Mux_v
    port map (
            O => \N__22525\,
            I => \N__22488\
        );

    \I__3235\ : Span4Mux_v
    port map (
            O => \N__22522\,
            I => \N__22488\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__22519\,
            I => \N__22481\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__22516\,
            I => \N__22481\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N__22481\
        );

    \I__3231\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22472\
        );

    \I__3230\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22472\
        );

    \I__3229\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22472\
        );

    \I__3228\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22472\
        );

    \I__3227\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22463\
        );

    \I__3226\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22463\
        );

    \I__3225\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22463\
        );

    \I__3224\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22463\
        );

    \I__3223\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22460\
        );

    \I__3222\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22453\
        );

    \I__3221\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22453\
        );

    \I__3220\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22453\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__22488\,
            I => \c0.n13033\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__22481\,
            I => \c0.n13033\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__22472\,
            I => \c0.n13033\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__22463\,
            I => \c0.n13033\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__22460\,
            I => \c0.n13033\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__22453\,
            I => \c0.n13033\
        );

    \I__3213\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22435\
        );

    \I__3212\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22431\
        );

    \I__3211\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22428\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__22435\,
            I => \N__22425\
        );

    \I__3209\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22422\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22419\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__22428\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__22425\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__22422\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__22419\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__3203\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__22407\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_26\
        );

    \I__3201\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__22401\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_27\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__22398\,
            I => \N__22394\
        );

    \I__3198\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22391\
        );

    \I__3197\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22388\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__22391\,
            I => \N__22385\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22378\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__22385\,
            I => \N__22378\
        );

    \I__3193\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22373\
        );

    \I__3192\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22373\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__22378\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__22373\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__3189\ : SRMux
    port map (
            O => \N__22368\,
            I => \N__22365\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22362\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__22359\,
            I => \c0.n3_adj_2287\
        );

    \I__3185\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22353\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__3183\ : Span4Mux_v
    port map (
            O => \N__22350\,
            I => \N__22347\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__22347\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_3\
        );

    \I__3181\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22340\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22337\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22332\
        );

    \I__3178\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22329\
        );

    \I__3177\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22326\
        );

    \I__3176\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22323\
        );

    \I__3175\ : Span4Mux_h
    port map (
            O => \N__22332\,
            I => \N__22320\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22313\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22313\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22313\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__22320\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__3170\ : Odrv12
    port map (
            O => \N__22313\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__3169\ : SRMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__3167\ : Span4Mux_v
    port map (
            O => \N__22302\,
            I => \N__22299\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__22299\,
            I => \c0.n3_adj_2340\
        );

    \I__3165\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__22290\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_28\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__3161\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22279\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \N__22276\
        );

    \I__3159\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22272\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22269\
        );

    \I__3157\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22266\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22263\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22260\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__22269\,
            I => \N__22253\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22253\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22253\
        );

    \I__3151\ : Odrv12
    port map (
            O => \N__22260\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__22253\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__3149\ : SRMux
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__22236\,
            I => \c0.n3_adj_2285\
        );

    \I__3144\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22227\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__22227\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_13\
        );

    \I__3141\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22218\
        );

    \I__3140\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22215\
        );

    \I__3139\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22212\
        );

    \I__3138\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22209\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22204\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__22215\,
            I => \N__22204\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22201\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__22209\,
            I => \N__22196\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__22204\,
            I => \N__22196\
        );

    \I__3132\ : Span4Mux_s2_h
    port map (
            O => \N__22201\,
            I => \N__22193\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__22196\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__22193\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__3129\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22185\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__22182\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_10\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__22179\,
            I => \N__22175\
        );

    \I__3125\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22172\
        );

    \I__3124\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22169\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__22172\,
            I => \N__22165\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22162\
        );

    \I__3121\ : InMux
    port map (
            O => \N__22168\,
            I => \N__22159\
        );

    \I__3120\ : Span4Mux_h
    port map (
            O => \N__22165\,
            I => \N__22153\
        );

    \I__3119\ : Span4Mux_v
    port map (
            O => \N__22162\,
            I => \N__22153\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__22150\
        );

    \I__3117\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22147\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__22153\,
            I => \N__22144\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__22150\,
            I => \N__22141\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22138\
        );

    \I__3113\ : Span4Mux_s1_h
    port map (
            O => \N__22144\,
            I => \N__22135\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__22141\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3111\ : Odrv12
    port map (
            O => \N__22138\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__22135\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__3109\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__3107\ : Span4Mux_h
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__22119\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_6\
        );

    \I__3105\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__3103\ : Span4Mux_h
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__22107\,
            I => \c0.n109\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__22101\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_11\
        );

    \I__3099\ : SRMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22095\,
            I => \N__22092\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__22089\,
            I => \c0.n3_adj_2324\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__22086\,
            I => \c0.n26_adj_2379_cascade_\
        );

    \I__3094\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__3092\ : Span12Mux_s4_h
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__3091\ : Odrv12
    port map (
            O => \N__22074\,
            I => \c0.n44_adj_2382\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__22071\,
            I => \N__22067\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__22070\,
            I => \N__22064\
        );

    \I__3088\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22061\
        );

    \I__3087\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22058\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22053\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22050\
        );

    \I__3084\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22045\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22045\
        );

    \I__3082\ : Odrv12
    port map (
            O => \N__22053\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__22050\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__22045\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__3079\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__22035\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_11\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__22032\,
            I => \N__22029\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22023\
        );

    \I__3075\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22018\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22018\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__22026\,
            I => \N__22015\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22010\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__22010\
        );

    \I__3070\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22007\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__22004\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__22007\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__22004\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__3066\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21996\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__21996\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_20\
        );

    \I__3064\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__21990\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_5\
        );

    \I__3062\ : SRMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21981\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__21981\,
            I => \c0.n3_adj_2336\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__3058\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21966\
        );

    \I__3056\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21963\
        );

    \I__3055\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21958\
        );

    \I__3054\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21958\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__21966\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__21963\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__21958\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__3050\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21944\
        );

    \I__3048\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21941\
        );

    \I__3047\ : Span4Mux_h
    port map (
            O => \N__21944\,
            I => \N__21938\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__21941\,
            I => \N__21935\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__21938\,
            I => \c0.n10_adj_2378\
        );

    \I__3044\ : Odrv12
    port map (
            O => \N__21935\,
            I => \c0.n10_adj_2378\
        );

    \I__3043\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__21927\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_4\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__21924\,
            I => \N__21908\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \N__21905\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__21922\,
            I => \N__21899\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__21921\,
            I => \N__21894\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__21920\,
            I => \N__21891\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__21919\,
            I => \N__21888\
        );

    \I__3035\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21876\
        );

    \I__3034\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21876\
        );

    \I__3033\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21871\
        );

    \I__3032\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21871\
        );

    \I__3031\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21863\
        );

    \I__3030\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21863\
        );

    \I__3029\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21863\
        );

    \I__3028\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21860\
        );

    \I__3027\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21847\
        );

    \I__3026\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21847\
        );

    \I__3025\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21847\
        );

    \I__3024\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21847\
        );

    \I__3023\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21847\
        );

    \I__3022\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21847\
        );

    \I__3021\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21834\
        );

    \I__3020\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21834\
        );

    \I__3019\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21834\
        );

    \I__3018\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21834\
        );

    \I__3017\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21834\
        );

    \I__3016\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21834\
        );

    \I__3015\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21821\
        );

    \I__3014\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21821\
        );

    \I__3013\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21821\
        );

    \I__3012\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21821\
        );

    \I__3011\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21821\
        );

    \I__3010\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21821\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21818\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__21871\,
            I => \N__21815\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__21870\,
            I => \N__21807\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21802\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__21860\,
            I => \N__21802\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21797\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__21834\,
            I => \N__21797\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21794\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__21818\,
            I => \N__21789\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__21815\,
            I => \N__21789\
        );

    \I__2999\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21781\
        );

    \I__2998\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21781\
        );

    \I__2997\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21781\
        );

    \I__2996\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21774\
        );

    \I__2995\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21774\
        );

    \I__2994\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21774\
        );

    \I__2993\ : Span12Mux_v
    port map (
            O => \N__21802\,
            I => \N__21771\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__21797\,
            I => \N__21768\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__21794\,
            I => \N__21763\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__21789\,
            I => \N__21763\
        );

    \I__2989\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21760\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__21781\,
            I => \c0.n7199\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__21774\,
            I => \c0.n7199\
        );

    \I__2986\ : Odrv12
    port map (
            O => \N__21771\,
            I => \c0.n7199\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__21768\,
            I => \c0.n7199\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__21763\,
            I => \c0.n7199\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__21760\,
            I => \c0.n7199\
        );

    \I__2982\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21742\
        );

    \I__2981\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21739\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__21745\,
            I => \N__21736\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__21742\,
            I => \N__21730\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__21739\,
            I => \N__21730\
        );

    \I__2977\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21725\
        );

    \I__2976\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21725\
        );

    \I__2975\ : Sp12to4
    port map (
            O => \N__21730\,
            I => \N__21720\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21720\
        );

    \I__2973\ : Odrv12
    port map (
            O => \N__21720\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__21717\,
            I => \N__21705\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__21716\,
            I => \N__21702\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__21715\,
            I => \N__21692\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__21714\,
            I => \N__21689\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__21713\,
            I => \N__21686\
        );

    \I__2967\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21679\
        );

    \I__2966\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21679\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__21710\,
            I => \N__21675\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__21709\,
            I => \N__21672\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__21708\,
            I => \N__21666\
        );

    \I__2962\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21656\
        );

    \I__2961\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21656\
        );

    \I__2960\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21656\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__21700\,
            I => \N__21653\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__21699\,
            I => \N__21650\
        );

    \I__2957\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21643\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__21697\,
            I => \N__21640\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__21696\,
            I => \N__21636\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21623\
        );

    \I__2953\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21623\
        );

    \I__2952\ : InMux
    port map (
            O => \N__21689\,
            I => \N__21623\
        );

    \I__2951\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21623\
        );

    \I__2950\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21623\
        );

    \I__2949\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21623\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21620\
        );

    \I__2947\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21611\
        );

    \I__2946\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21611\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21611\
        );

    \I__2944\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21611\
        );

    \I__2943\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21598\
        );

    \I__2942\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21598\
        );

    \I__2941\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21598\
        );

    \I__2940\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21598\
        );

    \I__2939\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21598\
        );

    \I__2938\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21598\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__21656\,
            I => \N__21595\
        );

    \I__2936\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21582\
        );

    \I__2935\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21582\
        );

    \I__2934\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21582\
        );

    \I__2933\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21582\
        );

    \I__2932\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21582\
        );

    \I__2931\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21582\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21579\
        );

    \I__2929\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21572\
        );

    \I__2928\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21572\
        );

    \I__2927\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21572\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__21623\,
            I => \N__21567\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__21620\,
            I => \N__21567\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__21611\,
            I => \c0.n10353\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__21598\,
            I => \c0.n10353\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__21595\,
            I => \c0.n10353\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__21582\,
            I => \c0.n10353\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__21579\,
            I => \c0.n10353\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21572\,
            I => \c0.n10353\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__21567\,
            I => \c0.n10353\
        );

    \I__2917\ : SRMux
    port map (
            O => \N__21552\,
            I => \N__21549\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__2915\ : Odrv12
    port map (
            O => \N__21546\,
            I => \c0.n3_adj_2338\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__21543\,
            I => \N__21539\
        );

    \I__2913\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21536\
        );

    \I__2912\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21532\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21512\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21500\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__21532\,
            I => \N__21497\
        );

    \I__2908\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21486\
        );

    \I__2907\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21486\
        );

    \I__2906\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21486\
        );

    \I__2905\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21486\
        );

    \I__2904\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21486\
        );

    \I__2903\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21473\
        );

    \I__2902\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21473\
        );

    \I__2901\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21473\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21473\
        );

    \I__2899\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21473\
        );

    \I__2898\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21473\
        );

    \I__2897\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21460\
        );

    \I__2896\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21460\
        );

    \I__2895\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21460\
        );

    \I__2894\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21460\
        );

    \I__2893\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21460\
        );

    \I__2892\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21460\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__21512\,
            I => \N__21457\
        );

    \I__2890\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21439\
        );

    \I__2889\ : InMux
    port map (
            O => \N__21510\,
            I => \N__21439\
        );

    \I__2888\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21439\
        );

    \I__2887\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21439\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21436\
        );

    \I__2885\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21427\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21427\
        );

    \I__2883\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21427\
        );

    \I__2882\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21427\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__21500\,
            I => \N__21424\
        );

    \I__2880\ : Span4Mux_s2_h
    port map (
            O => \N__21497\,
            I => \N__21412\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21412\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__21473\,
            I => \N__21412\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21412\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__21457\,
            I => \N__21409\
        );

    \I__2875\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21402\
        );

    \I__2874\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21402\
        );

    \I__2873\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21402\
        );

    \I__2872\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21399\
        );

    \I__2871\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21385\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21385\
        );

    \I__2869\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21385\
        );

    \I__2868\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21385\
        );

    \I__2867\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21385\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__21439\,
            I => \N__21382\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__21436\,
            I => \N__21379\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21376\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__21424\,
            I => \N__21367\
        );

    \I__2862\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21360\
        );

    \I__2861\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21360\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21360\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__21412\,
            I => \N__21357\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__21409\,
            I => \N__21354\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21349\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21349\
        );

    \I__2855\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21342\
        );

    \I__2854\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21342\
        );

    \I__2853\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21342\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21335\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__21382\,
            I => \N__21335\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__21379\,
            I => \N__21335\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__21376\,
            I => \N__21332\
        );

    \I__2848\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21323\
        );

    \I__2847\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21323\
        );

    \I__2846\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21323\
        );

    \I__2845\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21323\
        );

    \I__2844\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21318\
        );

    \I__2843\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21318\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__21367\,
            I => n63
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__21360\,
            I => n63
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__21357\,
            I => n63
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__21354\,
            I => n63
        );

    \I__2838\ : Odrv12
    port map (
            O => \N__21349\,
            I => n63
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__21342\,
            I => n63
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__21335\,
            I => n63
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__21332\,
            I => n63
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__21323\,
            I => n63
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__21318\,
            I => n63
        );

    \I__2832\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21292\
        );

    \I__2831\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21286\
        );

    \I__2830\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21283\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21280\
        );

    \I__2828\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21277\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21273\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__21289\,
            I => \N__21268\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__21286\,
            I => \N__21265\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21262\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__21280\,
            I => \N__21259\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__21277\,
            I => \N__21256\
        );

    \I__2821\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21247\
        );

    \I__2820\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21247\
        );

    \I__2819\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21244\
        );

    \I__2818\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21239\
        );

    \I__2817\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21239\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__21265\,
            I => \N__21234\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__21262\,
            I => \N__21234\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__21259\,
            I => \N__21229\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__21256\,
            I => \N__21229\
        );

    \I__2812\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21224\
        );

    \I__2811\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21224\
        );

    \I__2810\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21219\
        );

    \I__2809\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21219\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__21247\,
            I => \c0.n63_adj_2262\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__21244\,
            I => \c0.n63_adj_2262\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__21239\,
            I => \c0.n63_adj_2262\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__21234\,
            I => \c0.n63_adj_2262\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__21229\,
            I => \c0.n63_adj_2262\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__21224\,
            I => \c0.n63_adj_2262\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__21219\,
            I => \c0.n63_adj_2262\
        );

    \I__2801\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21198\
        );

    \I__2800\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21198\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__21198\,
            I => \N__21192\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21189\
        );

    \I__2797\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21186\
        );

    \I__2796\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21183\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21178\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__21189\,
            I => \N__21178\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21175\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21170\
        );

    \I__2791\ : Span4Mux_h
    port map (
            O => \N__21178\,
            I => \N__21158\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__21175\,
            I => \N__21158\
        );

    \I__2789\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21153\
        );

    \I__2788\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21153\
        );

    \I__2787\ : Span4Mux_h
    port map (
            O => \N__21170\,
            I => \N__21150\
        );

    \I__2786\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21147\
        );

    \I__2785\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21140\
        );

    \I__2784\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21140\
        );

    \I__2783\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21140\
        );

    \I__2782\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21137\
        );

    \I__2781\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21132\
        );

    \I__2780\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21132\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__21158\,
            I => n63_adj_2534
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__21153\,
            I => n63_adj_2534
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__21150\,
            I => n63_adj_2534
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__21147\,
            I => n63_adj_2534
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__21140\,
            I => n63_adj_2534
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__21137\,
            I => n63_adj_2534
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__21132\,
            I => n63_adj_2534
        );

    \I__2772\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__21111\,
            I => \c0.n113\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__2768\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21100\
        );

    \I__2767\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21097\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21094\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21090\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__21097\,
            I => \N__21085\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21085\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21082\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__21090\,
            I => \N__21077\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__21085\,
            I => \N__21077\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21074\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__21077\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__2757\ : Odrv12
    port map (
            O => \N__21074\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__2756\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__21063\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_14\
        );

    \I__2753\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__2751\ : Span4Mux_v
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__21051\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_28\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__21048\,
            I => \N__21043\
        );

    \I__2748\ : InMux
    port map (
            O => \N__21047\,
            I => \N__21040\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__21046\,
            I => \N__21037\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21033\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__21030\
        );

    \I__2744\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21027\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21024\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__21033\,
            I => \N__21021\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__21030\,
            I => \N__21018\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21027\,
            I => \N__21015\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21012\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__21021\,
            I => \N__21009\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__21018\,
            I => \N__21004\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__21015\,
            I => \N__21004\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__21012\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__21009\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__21004\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__2732\ : InMux
    port map (
            O => \N__20997\,
            I => \N__20994\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20991\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__20988\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_19\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__20985\,
            I => \N__20978\
        );

    \I__2727\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20972\
        );

    \I__2726\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20965\
        );

    \I__2725\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20965\
        );

    \I__2724\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20965\
        );

    \I__2723\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20962\
        );

    \I__2722\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20959\
        );

    \I__2721\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20956\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \N__20953\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__20972\,
            I => \N__20946\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20943\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__20962\,
            I => \N__20936\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__20959\,
            I => \N__20936\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20936\
        );

    \I__2714\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20927\
        );

    \I__2713\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20927\
        );

    \I__2712\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20927\
        );

    \I__2711\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20927\
        );

    \I__2710\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20924\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__20946\,
            I => \N__20921\
        );

    \I__2708\ : Span4Mux_s2_h
    port map (
            O => \N__20943\,
            I => \N__20914\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__20936\,
            I => \N__20914\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20914\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20911\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__20921\,
            I => \N__20908\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__20914\,
            I => \N__20905\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__20911\,
            I => \FRAME_MATCHER_i_31\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__20908\,
            I => \FRAME_MATCHER_i_31\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__20905\,
            I => \FRAME_MATCHER_i_31\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2698\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__20889\,
            I => \N__20886\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__20886\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_31\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__20883\,
            I => \n63_adj_2534_cascade_\
        );

    \I__2693\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20877\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20874\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__20874\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_18\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__20871\,
            I => \c0.n63_adj_2262_cascade_\
        );

    \I__2689\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__20865\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_5\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__20862\,
            I => \n11058_cascade_\
        );

    \I__2686\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__20850\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_3\
        );

    \I__2682\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__20844\,
            I => \N__20840\
        );

    \I__2680\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20837\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__20840\,
            I => \N__20833\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__20837\,
            I => \N__20830\
        );

    \I__2677\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20827\
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__20833\,
            I => \c0.n1502\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__20830\,
            I => \c0.n1502\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__20827\,
            I => \c0.n1502\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__20820\,
            I => \c0.n1502_cascade_\
        );

    \I__2672\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20811\
        );

    \I__2671\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20808\
        );

    \I__2670\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20803\
        );

    \I__2669\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20803\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__20811\,
            I => \N__20798\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__20808\,
            I => \N__20798\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20792\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__20798\,
            I => \N__20789\
        );

    \I__2664\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20782\
        );

    \I__2663\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20782\
        );

    \I__2662\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20782\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__20792\,
            I => \c0.n10522\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__20789\,
            I => \c0.n10522\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__20782\,
            I => \c0.n10522\
        );

    \I__2658\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__20772\,
            I => \c0.n4_adj_2266\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__20769\,
            I => \c0.n13033_cascade_\
        );

    \I__2655\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20762\
        );

    \I__2654\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20759\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20756\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__20756\,
            I => \N__20748\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__20753\,
            I => \N__20745\
        );

    \I__2649\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20740\
        );

    \I__2648\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20740\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__20748\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__20745\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__20740\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__2644\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__20724\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_30\
        );

    \I__2640\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20718\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__20718\,
            I => \N__20713\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__20717\,
            I => \N__20709\
        );

    \I__2637\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20706\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__20713\,
            I => \N__20703\
        );

    \I__2635\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20698\
        );

    \I__2634\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20698\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__20706\,
            I => \N__20695\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__20703\,
            I => \N__20692\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20689\
        );

    \I__2630\ : Odrv12
    port map (
            O => \N__20695\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__20692\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__20689\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__2627\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__20673\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_29\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__20670\,
            I => \n16802_cascade_\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__20667\,
            I => \c0.n10569_cascade_\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20655\
        );

    \I__2620\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20655\
        );

    \I__2619\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20655\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20650\
        );

    \I__2617\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20645\
        );

    \I__2616\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20645\
        );

    \I__2615\ : Odrv12
    port map (
            O => \N__20650\,
            I => data_in_frame_0_1
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__20645\,
            I => data_in_frame_0_1
        );

    \I__2613\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__2611\ : Span4Mux_h
    port map (
            O => \N__20634\,
            I => \N__20631\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__20631\,
            I => \N__20628\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__20628\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__20625\,
            I => \N__20621\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__20624\,
            I => \N__20618\
        );

    \I__2606\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20615\
        );

    \I__2605\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20612\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__20615\,
            I => \c0.data_in_frame_3_1\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__20612\,
            I => \c0.data_in_frame_3_1\
        );

    \I__2602\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20603\
        );

    \I__2601\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20600\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__20603\,
            I => \c0.n2137_adj_2237\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__20600\,
            I => \c0.n2137_adj_2237\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__20595\,
            I => \c0.n2137_adj_2237_cascade_\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__20592\,
            I => \N__20587\
        );

    \I__2596\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20584\
        );

    \I__2595\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20579\
        );

    \I__2594\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20579\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__20584\,
            I => data_in_frame_2_0
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__20579\,
            I => data_in_frame_2_0
        );

    \I__2591\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20569\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__20573\,
            I => \N__20566\
        );

    \I__2589\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20563\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__20569\,
            I => \N__20560\
        );

    \I__2587\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20557\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__20563\,
            I => data_in_frame_2_5
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__20560\,
            I => data_in_frame_2_5
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__20557\,
            I => data_in_frame_2_5
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__20550\,
            I => \N__20547\
        );

    \I__2582\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20543\
        );

    \I__2581\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20540\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__20543\,
            I => \N__20537\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__20540\,
            I => data_in_frame_5_6
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__20537\,
            I => data_in_frame_5_6
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__20532\,
            I => \N__20528\
        );

    \I__2576\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20523\
        );

    \I__2575\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20523\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__20523\,
            I => \c0.data_in_frame_3_0\
        );

    \I__2573\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20516\
        );

    \I__2572\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20513\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__20516\,
            I => \c0.n2126\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__20513\,
            I => \c0.n2126\
        );

    \I__2569\ : SRMux
    port map (
            O => \N__20508\,
            I => \N__20505\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20502\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__20502\,
            I => \c0.n8_adj_2249\
        );

    \I__2566\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20492\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__20498\,
            I => \N__20488\
        );

    \I__2564\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20485\
        );

    \I__2563\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20482\
        );

    \I__2562\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20479\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20476\
        );

    \I__2560\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20473\
        );

    \I__2559\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20470\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__20485\,
            I => \N__20465\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__20482\,
            I => \N__20465\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20462\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__20476\,
            I => \N__20457\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20457\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20454\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__20465\,
            I => \N__20449\
        );

    \I__2551\ : Span4Mux_s0_v
    port map (
            O => \N__20462\,
            I => \N__20449\
        );

    \I__2550\ : Span4Mux_h
    port map (
            O => \N__20457\,
            I => \N__20446\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__20454\,
            I => \N__20443\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__20449\,
            I => \c0.n4_adj_2349\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__20446\,
            I => \c0.n4_adj_2349\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__20443\,
            I => \c0.n4_adj_2349\
        );

    \I__2545\ : SRMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20430\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__20427\,
            I => \c0.n8_adj_2244\
        );

    \I__2541\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20419\
        );

    \I__2540\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20416\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20413\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__20419\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__20416\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__20413\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2534\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N__20397\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__20397\,
            I => \N__20392\
        );

    \I__2531\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20387\
        );

    \I__2530\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20387\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__20392\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__20387\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__2526\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20375\
        );

    \I__2525\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20372\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__20375\,
            I => \N__20368\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__20372\,
            I => \N__20365\
        );

    \I__2522\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20362\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__20368\,
            I => \N__20359\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__20365\,
            I => \N__20356\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__20362\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__20359\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__20356\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__2516\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__20343\,
            I => \N__20338\
        );

    \I__2513\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20335\
        );

    \I__2512\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20332\
        );

    \I__2511\ : Sp12to4
    port map (
            O => \N__20338\,
            I => \N__20327\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20327\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__20332\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__2508\ : Odrv12
    port map (
            O => \N__20327\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__20322\,
            I => \c0.n30_adj_2355_cascade_\
        );

    \I__2506\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20315\
        );

    \I__2505\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20312\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20309\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20305\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__20309\,
            I => \N__20302\
        );

    \I__2501\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20299\
        );

    \I__2500\ : Span4Mux_v
    port map (
            O => \N__20305\,
            I => \N__20296\
        );

    \I__2499\ : Span4Mux_s0_v
    port map (
            O => \N__20302\,
            I => \N__20293\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__20299\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__20296\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__20293\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__20283\,
            I => \c0.n51\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__20280\,
            I => \c0.n10613_cascade_\
        );

    \I__2492\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20274\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__20274\,
            I => \c0.n22_adj_2346\
        );

    \I__2490\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20268\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__2488\ : Span4Mux_s3_h
    port map (
            O => \N__20265\,
            I => \N__20262\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__20262\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_30\
        );

    \I__2486\ : InMux
    port map (
            O => \N__20259\,
            I => \c0.n16515\
        );

    \I__2485\ : InMux
    port map (
            O => \N__20256\,
            I => \c0.n16516\
        );

    \I__2484\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__20247\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_31\
        );

    \I__2481\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20241\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__20238\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_9\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__20235\,
            I => \N__20230\
        );

    \I__2477\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20224\
        );

    \I__2476\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20224\
        );

    \I__2475\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20221\
        );

    \I__2474\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20218\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20213\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__20221\,
            I => \N__20213\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__20218\,
            I => \N__20210\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__20213\,
            I => \N__20207\
        );

    \I__2469\ : Span4Mux_s3_h
    port map (
            O => \N__20210\,
            I => \N__20204\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__20207\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__20204\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__2466\ : SRMux
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__20187\,
            I => \c0.n3_adj_2328\
        );

    \I__2461\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__2459\ : Odrv12
    port map (
            O => \N__20178\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_6\
        );

    \I__2458\ : SRMux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__2456\ : Span4Mux_v
    port map (
            O => \N__20169\,
            I => \N__20166\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__20166\,
            I => \c0.n3_adj_2334\
        );

    \I__2454\ : CEMux
    port map (
            O => \N__20163\,
            I => \N__20160\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__20154\,
            I => \control.n18909\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__2448\ : Span4Mux_s1_v
    port map (
            O => \N__20145\,
            I => \N__20142\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__20139\,
            I => \c0.n8_adj_2254\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20133\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20129\
        );

    \I__2443\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20126\
        );

    \I__2442\ : Span4Mux_s3_v
    port map (
            O => \N__20129\,
            I => \N__20120\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__20126\,
            I => \N__20120\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20117\
        );

    \I__2439\ : Span4Mux_h
    port map (
            O => \N__20120\,
            I => \N__20114\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20117\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__20114\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__2436\ : SRMux
    port map (
            O => \N__20109\,
            I => \N__20106\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__20106\,
            I => \c0.n8_adj_2250\
        );

    \I__2434\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20093\
        );

    \I__2433\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20084\
        );

    \I__2432\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20081\
        );

    \I__2431\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20078\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20075\
        );

    \I__2429\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20072\
        );

    \I__2428\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20069\
        );

    \I__2427\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20066\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20062\
        );

    \I__2425\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20059\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20056\
        );

    \I__2423\ : InMux
    port map (
            O => \N__20090\,
            I => \N__20052\
        );

    \I__2422\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20049\
        );

    \I__2421\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20046\
        );

    \I__2420\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20043\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__20084\,
            I => \N__20038\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20035\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20024\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20024\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20024\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__20069\,
            I => \N__20024\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20024\
        );

    \I__2412\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20021\
        );

    \I__2411\ : Span4Mux_s2_v
    port map (
            O => \N__20062\,
            I => \N__20015\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__20059\,
            I => \N__20015\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20012\
        );

    \I__2408\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20009\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20002\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20002\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20002\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__19999\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20042\,
            I => \N__19996\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20041\,
            I => \N__19993\
        );

    \I__2401\ : Span4Mux_v
    port map (
            O => \N__20038\,
            I => \N__19983\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__20035\,
            I => \N__19983\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__20024\,
            I => \N__19983\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__19980\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20020\,
            I => \N__19977\
        );

    \I__2396\ : Span4Mux_h
    port map (
            O => \N__20015\,
            I => \N__19970\
        );

    \I__2395\ : Span4Mux_s2_v
    port map (
            O => \N__20012\,
            I => \N__19970\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__20009\,
            I => \N__19970\
        );

    \I__2393\ : Span4Mux_v
    port map (
            O => \N__20002\,
            I => \N__19963\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__19999\,
            I => \N__19963\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__19996\,
            I => \N__19963\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__19993\,
            I => \N__19960\
        );

    \I__2389\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19957\
        );

    \I__2388\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19954\
        );

    \I__2387\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19951\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__19983\,
            I => \c0.n4_adj_2271\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__19980\,
            I => \c0.n4_adj_2271\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__19977\,
            I => \c0.n4_adj_2271\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__19970\,
            I => \c0.n4_adj_2271\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__19963\,
            I => \c0.n4_adj_2271\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__19960\,
            I => \c0.n4_adj_2271\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__19957\,
            I => \c0.n4_adj_2271\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__19954\,
            I => \c0.n4_adj_2271\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__19951\,
            I => \c0.n4_adj_2271\
        );

    \I__2377\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19926\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__19923\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_22\
        );

    \I__2373\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19916\
        );

    \I__2372\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19912\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19909\
        );

    \I__2370\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19906\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19902\
        );

    \I__2368\ : Span4Mux_v
    port map (
            O => \N__19909\,
            I => \N__19897\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__19906\,
            I => \N__19897\
        );

    \I__2366\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19894\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__19902\,
            I => \N__19891\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__19897\,
            I => \N__19888\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19885\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__19891\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__19888\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__19885\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__2359\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__2357\ : Span4Mux_s3_h
    port map (
            O => \N__19872\,
            I => \N__19869\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__19869\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_22\
        );

    \I__2355\ : InMux
    port map (
            O => \N__19866\,
            I => \c0.n16507\
        );

    \I__2354\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19860\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__19857\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_23\
        );

    \I__2351\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19848\
        );

    \I__2350\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19845\
        );

    \I__2349\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19842\
        );

    \I__2348\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19839\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__19848\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__19845\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__19842\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__19839\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__2343\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__19827\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_23\
        );

    \I__2341\ : InMux
    port map (
            O => \N__19824\,
            I => \c0.n16508\
        );

    \I__2340\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__2338\ : Span4Mux_v
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__19812\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_24\
        );

    \I__2336\ : InMux
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19801\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19798\
        );

    \I__2333\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19794\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__19801\,
            I => \N__19791\
        );

    \I__2331\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19786\
        );

    \I__2330\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19786\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19783\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__19791\,
            I => \N__19780\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19777\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__19783\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__19780\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__19777\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__2323\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__19764\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_24\
        );

    \I__2320\ : InMux
    port map (
            O => \N__19761\,
            I => \bfn_4_14_0_\
        );

    \I__2319\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__19752\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_25\
        );

    \I__2316\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19743\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__19748\,
            I => \N__19740\
        );

    \I__2314\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19737\
        );

    \I__2313\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19734\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19731\
        );

    \I__2311\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19728\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__19737\,
            I => \N__19725\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__19734\,
            I => \N__19722\
        );

    \I__2308\ : Span4Mux_h
    port map (
            O => \N__19731\,
            I => \N__19719\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19716\
        );

    \I__2306\ : Span4Mux_h
    port map (
            O => \N__19725\,
            I => \N__19713\
        );

    \I__2305\ : Span4Mux_h
    port map (
            O => \N__19722\,
            I => \N__19710\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__19719\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__2303\ : Odrv12
    port map (
            O => \N__19716\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__19713\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__19710\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__2300\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__19695\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_25\
        );

    \I__2297\ : InMux
    port map (
            O => \N__19692\,
            I => \c0.n16510\
        );

    \I__2296\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__19686\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_26\
        );

    \I__2294\ : InMux
    port map (
            O => \N__19683\,
            I => \c0.n16511\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19680\,
            I => \c0.n16512\
        );

    \I__2292\ : InMux
    port map (
            O => \N__19677\,
            I => \c0.n16513\
        );

    \I__2291\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__19671\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_29\
        );

    \I__2289\ : InMux
    port map (
            O => \N__19668\,
            I => \c0.n16514\
        );

    \I__2288\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19659\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__19656\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_14\
        );

    \I__2284\ : InMux
    port map (
            O => \N__19653\,
            I => \c0.n16499\
        );

    \I__2283\ : InMux
    port map (
            O => \N__19650\,
            I => \N__19647\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__19644\,
            I => \N__19641\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__19641\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_15\
        );

    \I__2279\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19634\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19631\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19627\
        );

    \I__2276\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19624\
        );

    \I__2275\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19620\
        );

    \I__2274\ : Span4Mux_h
    port map (
            O => \N__19627\,
            I => \N__19617\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19614\
        );

    \I__2272\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19611\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__19620\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__19617\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__19614\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__19611\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__2267\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19599\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__19596\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_15\
        );

    \I__2264\ : InMux
    port map (
            O => \N__19593\,
            I => \c0.n16500\
        );

    \I__2263\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__19584\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_16\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__19581\,
            I => \N__19578\
        );

    \I__2259\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19574\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__19577\,
            I => \N__19570\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19567\
        );

    \I__2256\ : InMux
    port map (
            O => \N__19573\,
            I => \N__19561\
        );

    \I__2255\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19561\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__19567\,
            I => \N__19558\
        );

    \I__2253\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19555\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__19561\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__19558\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__19555\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__2249\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__19545\,
            I => \N__19542\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__19542\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_16\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19539\,
            I => \bfn_4_13_0_\
        );

    \I__2245\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__19527\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_17\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__2240\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19517\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19514\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__19517\,
            I => \N__19509\
        );

    \I__2237\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19506\
        );

    \I__2236\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19503\
        );

    \I__2235\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19500\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__19509\,
            I => \N__19497\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__19506\,
            I => \N__19494\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19491\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__19500\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__19497\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__19494\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__19491\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2227\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__19476\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_17\
        );

    \I__2224\ : InMux
    port map (
            O => \N__19473\,
            I => \c0.n16502\
        );

    \I__2223\ : InMux
    port map (
            O => \N__19470\,
            I => \c0.n16503\
        );

    \I__2222\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__19458\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_19\
        );

    \I__2218\ : InMux
    port map (
            O => \N__19455\,
            I => \c0.n16504\
        );

    \I__2217\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19449\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__19446\,
            I => \N__19443\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__19443\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_20\
        );

    \I__2213\ : InMux
    port map (
            O => \N__19440\,
            I => \c0.n16505\
        );

    \I__2212\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19434\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__19428\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_21\
        );

    \I__2208\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19418\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__19418\,
            I => \N__19412\
        );

    \I__2204\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19409\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__19412\,
            I => \N__19402\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19402\
        );

    \I__2201\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19397\
        );

    \I__2200\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19397\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__19402\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__19397\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__2197\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19389\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__19389\,
            I => \N__19386\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__19386\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_21\
        );

    \I__2194\ : InMux
    port map (
            O => \N__19383\,
            I => \c0.n16506\
        );

    \I__2193\ : InMux
    port map (
            O => \N__19380\,
            I => \c0.n16491\
        );

    \I__2192\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__19374\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_7\
        );

    \I__2190\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19368\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__19368\,
            I => \N__19362\
        );

    \I__2188\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19359\
        );

    \I__2187\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19356\
        );

    \I__2186\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19353\
        );

    \I__2185\ : Span4Mux_s3_h
    port map (
            O => \N__19362\,
            I => \N__19350\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__19359\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__19356\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__19353\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__19350\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__2180\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__19338\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_7\
        );

    \I__2178\ : InMux
    port map (
            O => \N__19335\,
            I => \c0.n16492\
        );

    \I__2177\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__19326\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_8\
        );

    \I__2174\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19319\
        );

    \I__2173\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19314\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19311\
        );

    \I__2171\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19308\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19305\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__19314\,
            I => \N__19302\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__19311\,
            I => \N__19297\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19297\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__19305\,
            I => \N__19294\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__19302\,
            I => \N__19291\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__19297\,
            I => \N__19288\
        );

    \I__2163\ : Span4Mux_s2_h
    port map (
            O => \N__19294\,
            I => \N__19285\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__19291\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__19288\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__19285\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__2159\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__19269\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_8\
        );

    \I__2155\ : InMux
    port map (
            O => \N__19266\,
            I => \bfn_4_12_0_\
        );

    \I__2154\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__19257\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_9\
        );

    \I__2151\ : InMux
    port map (
            O => \N__19254\,
            I => \c0.n16494\
        );

    \I__2150\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__2148\ : Span4Mux_s3_h
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__19242\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_10\
        );

    \I__2146\ : InMux
    port map (
            O => \N__19239\,
            I => \c0.n16495\
        );

    \I__2145\ : InMux
    port map (
            O => \N__19236\,
            I => \c0.n16496\
        );

    \I__2144\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__2142\ : Span4Mux_s3_h
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__19224\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_12\
        );

    \I__2140\ : InMux
    port map (
            O => \N__19221\,
            I => \c0.n16497\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19218\,
            I => \c0.n16498\
        );

    \I__2138\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__19212\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_0\
        );

    \I__2136\ : InMux
    port map (
            O => \N__19209\,
            I => \bfn_4_11_0_\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__2133\ : Span4Mux_s3_h
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__19197\,
            I => \c0.n27_adj_2426\
        );

    \I__2131\ : InMux
    port map (
            O => \N__19194\,
            I => \c0.n16486\
        );

    \I__2130\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__2128\ : Span4Mux_v
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__19182\,
            I => \c0.n115\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__2124\ : Span4Mux_s3_h
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__19170\,
            I => \c0.n29\
        );

    \I__2122\ : InMux
    port map (
            O => \N__19167\,
            I => \c0.n16487\
        );

    \I__2121\ : InMux
    port map (
            O => \N__19164\,
            I => \c0.n16488\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__19155\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_4\
        );

    \I__2117\ : InMux
    port map (
            O => \N__19152\,
            I => \c0.n16489\
        );

    \I__2116\ : InMux
    port map (
            O => \N__19149\,
            I => \c0.n16490\
        );

    \I__2115\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19120\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19120\
        );

    \I__2113\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19120\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19120\
        );

    \I__2111\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19104\
        );

    \I__2110\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19104\
        );

    \I__2109\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19104\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19104\
        );

    \I__2107\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19104\
        );

    \I__2106\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19104\
        );

    \I__2105\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19104\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19089\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19089\
        );

    \I__2102\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19089\
        );

    \I__2101\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19089\
        );

    \I__2100\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19089\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19089\
        );

    \I__2098\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19089\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19083\
        );

    \I__2096\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19080\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19075\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__19089\,
            I => \N__19075\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19072\
        );

    \I__2092\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19067\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19086\,
            I => \N__19067\
        );

    \I__2090\ : Span4Mux_s3_h
    port map (
            O => \N__19083\,
            I => \N__19063\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__19080\,
            I => \N__19060\
        );

    \I__2088\ : Span4Mux_s3_h
    port map (
            O => \N__19075\,
            I => \N__19053\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19053\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__19067\,
            I => \N__19053\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19050\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__19063\,
            I => \c0.n9575\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__19060\,
            I => \c0.n9575\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__19053\,
            I => \c0.n9575\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__19050\,
            I => \c0.n9575\
        );

    \I__2080\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19036\
        );

    \I__2079\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19033\
        );

    \I__2078\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19030\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__19036\,
            I => n12966
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19033\,
            I => n12966
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19030\,
            I => n12966
        );

    \I__2074\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19020\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__19020\,
            I => \N__19017\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__19017\,
            I => \N__19013\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19010\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__19013\,
            I => n15118
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__19010\,
            I => n15118
        );

    \I__2068\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18997\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18994\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19003\,
            I => \N__18991\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18986\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18986\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18983\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__18997\,
            I => \N__18980\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18977\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__18991\,
            I => \N__18974\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18969\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18969\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__18980\,
            I => \N__18966\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__18977\,
            I => \N__18963\
        );

    \I__2055\ : Span4Mux_s2_h
    port map (
            O => \N__18974\,
            I => \N__18958\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__18969\,
            I => \N__18958\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__18966\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__18963\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__18958\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__18951\,
            I => \c0.n16685_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__18945\,
            I => \c0.n6_adj_2267\
        );

    \I__2047\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18937\
        );

    \I__2046\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18932\
        );

    \I__2045\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18932\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18929\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18926\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__18929\,
            I => \N__18921\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__18926\,
            I => \N__18918\
        );

    \I__2040\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18913\
        );

    \I__2039\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18913\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__18921\,
            I => \FRAME_MATCHER_i_31__N_1270\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__18918\,
            I => \FRAME_MATCHER_i_31__N_1270\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__18913\,
            I => \FRAME_MATCHER_i_31__N_1270\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__18906\,
            I => \N__18902\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__18905\,
            I => \N__18899\
        );

    \I__2033\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18894\
        );

    \I__2032\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18894\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__18894\,
            I => \N__18891\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__18891\,
            I => \c0.n7528\
        );

    \I__2029\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18884\
        );

    \I__2028\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18881\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__18884\,
            I => \N__18878\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__18881\,
            I => \N__18875\
        );

    \I__2025\ : Span4Mux_s3_h
    port map (
            O => \N__18878\,
            I => \N__18872\
        );

    \I__2024\ : Span12Mux_s3_v
    port map (
            O => \N__18875\,
            I => \N__18869\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__18872\,
            I => \c0.n46\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__18869\,
            I => \c0.n46\
        );

    \I__2021\ : SRMux
    port map (
            O => \N__18864\,
            I => \N__18861\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__18861\,
            I => \N__18858\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__18858\,
            I => \N__18855\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__18855\,
            I => \c0.n3_adj_2332\
        );

    \I__2017\ : SRMux
    port map (
            O => \N__18852\,
            I => \N__18849\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__18849\,
            I => \N__18846\
        );

    \I__2015\ : Span4Mux_s3_h
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__18840\,
            I => \c0.n3_adj_2330\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__18837\,
            I => \c0.n9575_cascade_\
        );

    \I__2011\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18830\
        );

    \I__2010\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18827\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__18830\,
            I => n12999
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__18827\,
            I => n12999
        );

    \I__2007\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__18819\,
            I => \N__18815\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18812\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__18815\,
            I => \N__18809\
        );

    \I__2003\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18806\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__18809\,
            I => \c0.n232\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__18806\,
            I => \c0.n232\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__18801\,
            I => \n12999_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18795\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__18792\,
            I => n18
        );

    \I__1996\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18786\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__18780\,
            I => \c0.n10346\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \c0.n17_cascade_\
        );

    \I__1991\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18771\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__18771\,
            I => \c0.n25_adj_2352\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__18768\,
            I => \c0.n17962_cascade_\
        );

    \I__1988\ : SRMux
    port map (
            O => \N__18765\,
            I => \N__18762\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__18762\,
            I => \N__18759\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__18759\,
            I => \N__18756\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__18756\,
            I => \c0.n4_adj_2226\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__18753\,
            I => \c0.n2126_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__18747\,
            I => \c0.n27\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__18744\,
            I => \c0.n23_cascade_\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__18741\,
            I => \c0.n30_cascade_\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__18738\,
            I => \c0.n50_cascade_\
        );

    \I__1978\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18732\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18727\
        );

    \I__1976\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18722\
        );

    \I__1975\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18722\
        );

    \I__1974\ : Span4Mux_s3_h
    port map (
            O => \N__18727\,
            I => \N__18717\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__18722\,
            I => \N__18717\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__18717\,
            I => n13849
        );

    \I__1971\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__18711\,
            I => \c0.n19_adj_2351\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__18708\,
            I => \c0.n8_adj_2273_cascade_\
        );

    \I__1968\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18698\
        );

    \I__1967\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18689\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18689\
        );

    \I__1965\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18689\
        );

    \I__1964\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18689\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__18698\,
            I => \c0.n8_adj_2273\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__18689\,
            I => \c0.n8_adj_2273\
        );

    \I__1961\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18680\
        );

    \I__1960\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18676\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__18680\,
            I => \N__18673\
        );

    \I__1958\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18670\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__18676\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__18673\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__18670\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__1954\ : SRMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__1952\ : Odrv12
    port map (
            O => \N__18657\,
            I => \c0.n17273\
        );

    \I__1951\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18649\
        );

    \I__1950\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18646\
        );

    \I__1949\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18643\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__18649\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__18646\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18643\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__1945\ : SRMux
    port map (
            O => \N__18636\,
            I => \N__18633\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__18633\,
            I => \c0.n17299\
        );

    \I__1943\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18627\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18624\
        );

    \I__1941\ : Odrv12
    port map (
            O => \N__18624\,
            I => \c0.n45\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__18621\,
            I => \N__18618\
        );

    \I__1939\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18615\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__18612\,
            I => \c0.n46_adj_2356\
        );

    \I__1936\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18606\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__18606\,
            I => \c0.n56\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__18603\,
            I => \c0.n10513_cascade_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18591\
        );

    \I__1932\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18591\
        );

    \I__1931\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18587\
        );

    \I__1930\ : InMux
    port map (
            O => \N__18597\,
            I => \N__18582\
        );

    \I__1929\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18582\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__18591\,
            I => \N__18579\
        );

    \I__1927\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18576\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18571\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__18582\,
            I => \N__18571\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__18579\,
            I => \N__18566\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__18576\,
            I => \N__18566\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__18571\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__18566\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__18561\,
            I => \c0.n6033_cascade_\
        );

    \I__1919\ : IoInMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__1917\ : Span4Mux_s3_v
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__18549\,
            I => \PIN_2_c_1\
        );

    \I__1915\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18541\
        );

    \I__1914\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18538\
        );

    \I__1913\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18535\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18530\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__18538\,
            I => \N__18530\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__18535\,
            I => \N__18525\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__18530\,
            I => \N__18525\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__18525\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__1907\ : SRMux
    port map (
            O => \N__18522\,
            I => \N__18519\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__1905\ : Span4Mux_s1_v
    port map (
            O => \N__18516\,
            I => \N__18513\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__18513\,
            I => \c0.n8_adj_2245\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__1902\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18503\
        );

    \I__1901\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18499\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__18503\,
            I => \N__18496\
        );

    \I__1899\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18493\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18499\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__18496\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__18493\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__1895\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18477\
        );

    \I__1894\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18477\
        );

    \I__1893\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18477\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__18477\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__1891\ : SRMux
    port map (
            O => \N__18474\,
            I => \N__18471\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__18471\,
            I => \N__18468\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__18468\,
            I => \c0.n17293\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__18465\,
            I => \N__18460\
        );

    \I__1887\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18457\
        );

    \I__1886\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18452\
        );

    \I__1885\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18452\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__18457\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__18452\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__1882\ : SRMux
    port map (
            O => \N__18447\,
            I => \N__18444\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__1880\ : Span4Mux_s1_v
    port map (
            O => \N__18441\,
            I => \N__18438\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__18438\,
            I => \c0.n8_adj_2247\
        );

    \I__1878\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18406\
        );

    \I__1877\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18406\
        );

    \I__1876\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18406\
        );

    \I__1875\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18406\
        );

    \I__1874\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18406\
        );

    \I__1873\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18406\
        );

    \I__1872\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18406\
        );

    \I__1871\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18391\
        );

    \I__1870\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18391\
        );

    \I__1869\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18391\
        );

    \I__1868\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18391\
        );

    \I__1867\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18391\
        );

    \I__1866\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18391\
        );

    \I__1865\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18391\
        );

    \I__1864\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18388\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__18406\,
            I => \N__18385\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__18391\,
            I => \N__18374\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__18388\,
            I => \N__18371\
        );

    \I__1860\ : Span4Mux_s2_h
    port map (
            O => \N__18385\,
            I => \N__18368\
        );

    \I__1859\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18353\
        );

    \I__1858\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18353\
        );

    \I__1857\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18353\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18353\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18353\
        );

    \I__1854\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18353\
        );

    \I__1853\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18353\
        );

    \I__1852\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18350\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__18374\,
            I => \N__18345\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__18371\,
            I => \N__18345\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__18368\,
            I => \c0.n10497\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__18353\,
            I => \c0.n10497\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__18350\,
            I => \c0.n10497\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__18345\,
            I => \c0.n10497\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__1844\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18327\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__18324\,
            I => \c0.n2_adj_2315\
        );

    \I__1840\ : SRMux
    port map (
            O => \N__18321\,
            I => \N__18318\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__18318\,
            I => \c0.n3_adj_2289\
        );

    \I__1838\ : SRMux
    port map (
            O => \N__18315\,
            I => \N__18312\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__18312\,
            I => \c0.n3_adj_2283\
        );

    \I__1836\ : SRMux
    port map (
            O => \N__18309\,
            I => \N__18306\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__1834\ : Span12Mux_v
    port map (
            O => \N__18303\,
            I => \N__18300\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__18300\,
            I => \c0.n3_adj_2279\
        );

    \I__1832\ : SRMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__18294\,
            I => \N__18291\
        );

    \I__1830\ : Span4Mux_s3_h
    port map (
            O => \N__18291\,
            I => \N__18288\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__18288\,
            I => \c0.n3_adj_2303\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__18285\,
            I => \c0.n10353_cascade_\
        );

    \I__1827\ : SRMux
    port map (
            O => \N__18282\,
            I => \N__18279\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__18279\,
            I => \N__18276\
        );

    \I__1825\ : Span4Mux_s2_h
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__18273\,
            I => \c0.n3_adj_2345\
        );

    \I__1823\ : SRMux
    port map (
            O => \N__18270\,
            I => \N__18267\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__18264\,
            I => \N__18261\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__18261\,
            I => \c0.n3_adj_2343\
        );

    \I__1819\ : SRMux
    port map (
            O => \N__18258\,
            I => \N__18255\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__18252\,
            I => \N__18249\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__18249\,
            I => \c0.n3\
        );

    \I__1815\ : SRMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__1813\ : Span4Mux_s3_h
    port map (
            O => \N__18240\,
            I => \N__18237\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__18237\,
            I => \c0.n3_adj_2295\
        );

    \I__1811\ : SRMux
    port map (
            O => \N__18234\,
            I => \N__18231\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__18231\,
            I => \N__18228\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__1808\ : Span4Mux_s2_h
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__18222\,
            I => \c0.n3_adj_2291\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__18219\,
            I => \c0.n232_cascade_\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__18216\,
            I => \N__18213\
        );

    \I__1804\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__18210\,
            I => \N__18207\
        );

    \I__1802\ : Span4Mux_s2_h
    port map (
            O => \N__18207\,
            I => \N__18204\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__18204\,
            I => \c0.n6_adj_2364\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__18201\,
            I => \N__18198\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18195\,
            I => n237
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__18192\,
            I => \n237_cascade_\
        );

    \I__1796\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18186\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__18186\,
            I => n22_adj_2465
        );

    \I__1794\ : SRMux
    port map (
            O => \N__18183\,
            I => \N__18180\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__18180\,
            I => \N__18177\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__18177\,
            I => \c0.n3_adj_2309\
        );

    \I__1791\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18168\
        );

    \I__1790\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18168\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__18168\,
            I => \N__18165\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__18165\,
            I => n1437
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__18162\,
            I => \N__18157\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18153\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18146\
        );

    \I__1784\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18146\
        );

    \I__1783\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18146\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__18153\,
            I => \N__18143\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18140\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__18143\,
            I => n8_adj_2498
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__18140\,
            I => n8_adj_2498
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__18135\,
            I => \c0.n6_adj_2265_cascade_\
        );

    \I__1777\ : SRMux
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__1775\ : Span4Mux_s3_h
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__18123\,
            I => \c0.n18907\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__18120\,
            I => \n13_adj_2469_cascade_\
        );

    \I__1772\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__18111\,
            I => n7
        );

    \I__1769\ : SRMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__1767\ : Span4Mux_s2_h
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__18099\,
            I => \c0.n3_adj_2301\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__18096\,
            I => \n1166_cascade_\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18086\
        );

    \I__1762\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18083\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__18086\,
            I => \N__18077\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__18083\,
            I => \N__18077\
        );

    \I__1759\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18074\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__18077\,
            I => \N__18071\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__18074\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__18071\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__18066\,
            I => \c0.n10497_cascade_\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__18063\,
            I => \N__18052\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__18062\,
            I => \N__18048\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__18061\,
            I => \N__18044\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__18060\,
            I => \N__18037\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__18059\,
            I => \N__18033\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18029\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__18057\,
            I => \N__18024\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__18056\,
            I => \N__18021\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__18055\,
            I => \N__18018\
        );

    \I__1745\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18000\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18000\
        );

    \I__1743\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18000\
        );

    \I__1742\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18000\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18000\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18043\,
            I => \N__18000\
        );

    \I__1739\ : InMux
    port map (
            O => \N__18042\,
            I => \N__18000\
        );

    \I__1738\ : InMux
    port map (
            O => \N__18041\,
            I => \N__17997\
        );

    \I__1737\ : InMux
    port map (
            O => \N__18040\,
            I => \N__17994\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18037\,
            I => \N__17979\
        );

    \I__1735\ : InMux
    port map (
            O => \N__18036\,
            I => \N__17979\
        );

    \I__1734\ : InMux
    port map (
            O => \N__18033\,
            I => \N__17979\
        );

    \I__1733\ : InMux
    port map (
            O => \N__18032\,
            I => \N__17979\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18029\,
            I => \N__17979\
        );

    \I__1731\ : InMux
    port map (
            O => \N__18028\,
            I => \N__17979\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17979\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18024\,
            I => \N__17966\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18021\,
            I => \N__17966\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18018\,
            I => \N__17966\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18017\,
            I => \N__17966\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18016\,
            I => \N__17966\
        );

    \I__1724\ : InMux
    port map (
            O => \N__18015\,
            I => \N__17966\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__18000\,
            I => \c0.n17713\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__17997\,
            I => \c0.n17713\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__17994\,
            I => \c0.n17713\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__17979\,
            I => \c0.n17713\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__17966\,
            I => \c0.n17713\
        );

    \I__1718\ : SRMux
    port map (
            O => \N__17955\,
            I => \N__17952\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__17952\,
            I => \N__17949\
        );

    \I__1716\ : Span4Mux_s2_h
    port map (
            O => \N__17949\,
            I => \N__17946\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__17946\,
            I => \c0.n17239\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__17943\,
            I => \N__17940\
        );

    \I__1713\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17937\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17933\
        );

    \I__1711\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17929\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__17933\,
            I => \N__17926\
        );

    \I__1709\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17923\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__17929\,
            I => n15
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__17926\,
            I => n15
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__17923\,
            I => n15
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__17916\,
            I => \n17694_cascade_\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__17913\,
            I => \N__17908\
        );

    \I__1703\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17905\
        );

    \I__1702\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17900\
        );

    \I__1701\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17900\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17897\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__17900\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__17897\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__1697\ : SRMux
    port map (
            O => \N__17892\,
            I => \N__17889\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17886\
        );

    \I__1695\ : Span4Mux_s3_h
    port map (
            O => \N__17886\,
            I => \N__17883\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__17883\,
            I => \c0.n17279\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__17880\,
            I => \FRAME_MATCHER_state_31_N_1406_0_cascade_\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__17877\,
            I => \N__17873\
        );

    \I__1691\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17867\
        );

    \I__1690\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17867\
        );

    \I__1689\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17864\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__17867\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__17864\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__1686\ : SRMux
    port map (
            O => \N__17859\,
            I => \N__17856\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17853\
        );

    \I__1684\ : Span4Mux_s3_h
    port map (
            O => \N__17853\,
            I => \N__17850\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__17850\,
            I => \c0.n8_adj_2252\
        );

    \I__1682\ : SRMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__1680\ : Span4Mux_s1_v
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__17838\,
            I => \c0.n8_adj_2246\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__17835\,
            I => \N__17831\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__17834\,
            I => \N__17828\
        );

    \I__1676\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17825\
        );

    \I__1675\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17822\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17816\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17816\
        );

    \I__1672\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17813\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__17816\,
            I => \N__17810\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__17813\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__17810\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__1668\ : SRMux
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__17802\,
            I => \N__17799\
        );

    \I__1666\ : Span4Mux_s2_h
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__17796\,
            I => \c0.n17277\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \N__17789\
        );

    \I__1663\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17786\
        );

    \I__1662\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17783\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__17786\,
            I => \N__17779\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17776\
        );

    \I__1659\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17773\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__17779\,
            I => \N__17770\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__17776\,
            I => \N__17767\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__17773\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__17770\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__17767\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__1653\ : SRMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__17757\,
            I => \N__17754\
        );

    \I__1651\ : Span4Mux_s3_v
    port map (
            O => \N__17754\,
            I => \N__17751\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__17751\,
            I => \c0.n17283\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__17748\,
            I => \N__17744\
        );

    \I__1648\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__1647\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17737\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17734\
        );

    \I__1645\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17731\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__17737\,
            I => \N__17726\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__17734\,
            I => \N__17726\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__17731\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__17726\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__1640\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17718\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__17718\,
            I => \N__17713\
        );

    \I__1638\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17710\
        );

    \I__1637\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17707\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__17713\,
            I => \N__17704\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__17710\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__17707\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__17704\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__17697\,
            I => \N__17694\
        );

    \I__1631\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17691\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17686\
        );

    \I__1629\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17683\
        );

    \I__1628\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17680\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__17686\,
            I => \N__17677\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__17683\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__17680\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__17677\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__17670\,
            I => \c0.n49_cascade_\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__17667\,
            I => \N__17662\
        );

    \I__1621\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17659\
        );

    \I__1620\ : InMux
    port map (
            O => \N__17665\,
            I => \N__17656\
        );

    \I__1619\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17653\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17650\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17656\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__17653\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__17650\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__17643\,
            I => \N__17640\
        );

    \I__1613\ : InMux
    port map (
            O => \N__17640\,
            I => \N__17637\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__17637\,
            I => \N__17633\
        );

    \I__1611\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17629\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__17633\,
            I => \N__17626\
        );

    \I__1609\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17623\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__17629\,
            I => \N__17620\
        );

    \I__1607\ : Span4Mux_s1_h
    port map (
            O => \N__17626\,
            I => \N__17617\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__17623\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__17620\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__17617\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__1603\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17607\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__17607\,
            I => \c0.n50_adj_2353\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__17604\,
            I => \N__17600\
        );

    \I__1600\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17594\
        );

    \I__1599\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17594\
        );

    \I__1598\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17591\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__17594\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__17591\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__1595\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17583\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__17583\,
            I => \c0.n47\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__1592\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17572\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \N__17569\
        );

    \I__1590\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17566\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17563\
        );

    \I__1588\ : InMux
    port map (
            O => \N__17569\,
            I => \N__17560\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__17566\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__17563\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__17560\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__17553\,
            I => \N__17550\
        );

    \I__1583\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17546\
        );

    \I__1582\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17542\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17539\
        );

    \I__1580\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17536\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__17542\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__17539\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17536\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__1576\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17526\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__17526\,
            I => \c0.n48\
        );

    \I__1574\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17514\
        );

    \I__1573\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17514\
        );

    \I__1572\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17514\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__17514\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__1570\ : SRMux
    port map (
            O => \N__17511\,
            I => \N__17508\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__17508\,
            I => \N__17505\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__17505\,
            I => \c0.n17275\
        );

    \I__1567\ : SRMux
    port map (
            O => \N__17502\,
            I => \N__17499\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__17499\,
            I => \N__17496\
        );

    \I__1565\ : Sp12to4
    port map (
            O => \N__17496\,
            I => \N__17493\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__17493\,
            I => \c0.n3_adj_2293\
        );

    \I__1563\ : SRMux
    port map (
            O => \N__17490\,
            I => \N__17487\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__17487\,
            I => \N__17484\
        );

    \I__1561\ : Span4Mux_s1_h
    port map (
            O => \N__17484\,
            I => \N__17481\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__17481\,
            I => \c0.n3_adj_2297\
        );

    \I__1559\ : SRMux
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17472\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__17472\,
            I => \c0.n3_adj_2326\
        );

    \I__1556\ : SRMux
    port map (
            O => \N__17469\,
            I => \N__17466\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__17466\,
            I => \N__17463\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__17463\,
            I => \N__17460\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__17460\,
            I => \c0.n3_adj_2313\
        );

    \I__1552\ : SRMux
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17451\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__17451\,
            I => \c0.n3_adj_2281\
        );

    \I__1549\ : SRMux
    port map (
            O => \N__17448\,
            I => \N__17445\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__17445\,
            I => \N__17442\
        );

    \I__1547\ : Span4Mux_s1_h
    port map (
            O => \N__17442\,
            I => \N__17439\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__17439\,
            I => \c0.n3_adj_2322\
        );

    \I__1545\ : SRMux
    port map (
            O => \N__17436\,
            I => \N__17433\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__17430\,
            I => \c0.n3_adj_2311\
        );

    \I__1542\ : SRMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17421\
        );

    \I__1540\ : Span4Mux_s1_h
    port map (
            O => \N__17421\,
            I => \N__17418\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__17418\,
            I => \c0.n3_adj_2307\
        );

    \I__1538\ : InMux
    port map (
            O => \N__17415\,
            I => \N__17412\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__17412\,
            I => \N__17409\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__17409\,
            I => \c0.n42\
        );

    \I__1535\ : SRMux
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17400\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__17400\,
            I => \c0.n3_adj_2299\
        );

    \I__1532\ : SRMux
    port map (
            O => \N__17397\,
            I => \N__17394\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__17394\,
            I => \N__17391\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__17391\,
            I => \c0.n8_adj_2258\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__17388\,
            I => \c0.n39_cascade_\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__17385\,
            I => \c0.n48_adj_2383_cascade_\
        );

    \I__1527\ : InMux
    port map (
            O => \N__17382\,
            I => \N__17379\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__17379\,
            I => \c0.n40\
        );

    \I__1525\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17373\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__17373\,
            I => \c0.n41\
        );

    \I__1523\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17367\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__17367\,
            I => \c0.n43_adj_2384\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__17364\,
            I => \c0.n17713_cascade_\
        );

    \I__1520\ : SRMux
    port map (
            O => \N__17361\,
            I => \N__17358\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__17358\,
            I => \N__17355\
        );

    \I__1518\ : Span4Mux_s3_v
    port map (
            O => \N__17355\,
            I => \N__17352\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__17352\,
            I => \c0.n8_adj_2234\
        );

    \I__1516\ : SRMux
    port map (
            O => \N__17349\,
            I => \N__17346\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__17343\,
            I => \c0.n17281\
        );

    \I__1513\ : SRMux
    port map (
            O => \N__17340\,
            I => \N__17337\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__17337\,
            I => \N__17334\
        );

    \I__1511\ : Span4Mux_s1_h
    port map (
            O => \N__17334\,
            I => \N__17331\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__17331\,
            I => \c0.n17259\
        );

    \I__1509\ : SRMux
    port map (
            O => \N__17328\,
            I => \N__17325\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__17325\,
            I => \c0.n17261\
        );

    \I__1507\ : SRMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17316\
        );

    \I__1505\ : Span4Mux_s2_h
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__17313\,
            I => \c0.n13900\
        );

    \I__1503\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17305\
        );

    \I__1502\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17300\
        );

    \I__1501\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17300\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__17305\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__17300\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__1498\ : SRMux
    port map (
            O => \N__17295\,
            I => \N__17292\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__17292\,
            I => \N__17289\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__17286\,
            I => \c0.n8_adj_2257\
        );

    \I__1494\ : SRMux
    port map (
            O => \N__17283\,
            I => \N__17280\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__17280\,
            I => \N__17277\
        );

    \I__1492\ : Span4Mux_s2_h
    port map (
            O => \N__17277\,
            I => \N__17274\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__17274\,
            I => \c0.n17263\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__17271\,
            I => \N__17268\
        );

    \I__1489\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17265\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__17265\,
            I => \N__17260\
        );

    \I__1487\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17257\
        );

    \I__1486\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17254\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__17260\,
            I => \N__17251\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__17257\,
            I => \N__17248\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__17254\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__17251\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__1481\ : Odrv12
    port map (
            O => \N__17248\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__1480\ : SRMux
    port map (
            O => \N__17241\,
            I => \N__17238\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__17238\,
            I => \N__17235\
        );

    \I__1478\ : Span4Mux_s1_h
    port map (
            O => \N__17235\,
            I => \N__17232\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__17232\,
            I => \c0.n17265\
        );

    \I__1476\ : InMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__17226\,
            I => \N__17221\
        );

    \I__1474\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17218\
        );

    \I__1473\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17215\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__17221\,
            I => \N__17210\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17210\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__17215\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__17210\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__1468\ : SRMux
    port map (
            O => \N__17205\,
            I => \N__17202\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__17202\,
            I => \N__17199\
        );

    \I__1466\ : Sp12to4
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__1465\ : Odrv12
    port map (
            O => \N__17196\,
            I => \c0.n17267\
        );

    \I__1464\ : SRMux
    port map (
            O => \N__17193\,
            I => \N__17190\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__17190\,
            I => \c0.n17269\
        );

    \I__1462\ : SRMux
    port map (
            O => \N__17187\,
            I => \N__17184\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__17184\,
            I => \N__17181\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__17181\,
            I => \N__17178\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__17178\,
            I => \c0.n17303\
        );

    \I__1458\ : SRMux
    port map (
            O => \N__17175\,
            I => \N__17172\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17169\
        );

    \I__1456\ : Span4Mux_s1_h
    port map (
            O => \N__17169\,
            I => \N__17166\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__17166\,
            I => \c0.n17271\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__17163\,
            I => \n10429_cascade_\
        );

    \I__1453\ : InMux
    port map (
            O => \N__17160\,
            I => \N__17157\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__17157\,
            I => n12965
        );

    \I__1451\ : InMux
    port map (
            O => \N__17154\,
            I => \N__17151\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__17151\,
            I => n242
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__17148\,
            I => \n12965_cascade_\
        );

    \I__1448\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17142\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__17142\,
            I => n10429
        );

    \I__1446\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17136\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__17133\,
            I => n8_adj_2541
        );

    \I__1443\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17127\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__17127\,
            I => n18_adj_2539
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__17124\,
            I => \n21_adj_2538_cascade_\
        );

    \I__1440\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17118\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__17118\,
            I => n15_adj_2540
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__17115\,
            I => \c0.n4_adj_2271_cascade_\
        );

    \I__1437\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17109\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__17109\,
            I => \c0.n2_adj_2341\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__17106\,
            I => \c0.n2_adj_2341_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17100\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__17100\,
            I => \c0.n10425\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__17097\,
            I => \N__17094\
        );

    \I__1431\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17091\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__17091\,
            I => \c0.n10465\
        );

    \I__1429\ : IoInMux
    port map (
            O => \N__17088\,
            I => \N__17085\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__17085\,
            I => \N__17082\
        );

    \I__1427\ : IoSpan4Mux
    port map (
            O => \N__17082\,
            I => \N__17079\
        );

    \I__1426\ : IoSpan4Mux
    port map (
            O => \N__17079\,
            I => \N__17076\
        );

    \I__1425\ : IoSpan4Mux
    port map (
            O => \N__17076\,
            I => \N__17073\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__17073\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16585,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16593,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16601,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16554,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16562,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16570,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \control.n16654\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n16546\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n16531\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16641\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16493\,
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16501\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16509\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16616,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16624,
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16632,
            carryinitout => \bfn_6_24_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17088\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i4_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20308\,
            in2 => \_gnd_net_\,
            in3 => \N__20091\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49785\,
            ce => 'H',
            sr => \N__17361\
        );

    \c0.FRAME_MATCHER_state_i11_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17263\,
            in2 => \_gnd_net_\,
            in3 => \N__20065\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49769\,
            ce => 'H',
            sr => \N__17241\
        );

    \c0.FRAME_MATCHER_state_i12_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17224\,
            in2 => \_gnd_net_\,
            in3 => \N__20041\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49756\,
            ce => 'H',
            sr => \N__17205\
        );

    \c0.FRAME_MATCHER_state_i15_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17665\,
            in2 => \_gnd_net_\,
            in3 => \N__19991\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49743\,
            ce => 'H',
            sr => \N__17175\
        );

    \c0.i1_4_lut_adj_507_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__18596\,
            in1 => \N__17112\,
            in2 => \N__17097\,
            in3 => \N__21297\,
            lcout => \c0.n4_adj_2271\,
            ltout => \c0.n4_adj_2271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i8_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__17309\,
            in1 => \_gnd_net_\,
            in2 => \N__17115\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49731\,
            ce => 'H',
            sr => \N__17295\
        );

    \c0.i16_4_lut_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17225\,
            in1 => \N__17264\,
            in2 => \N__17793\,
            in3 => \N__17308\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_620_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30517\,
            in1 => \N__21915\,
            in2 => \N__28712\,
            in3 => \N__21505\,
            lcout => \c0.n2_adj_2341\,
            ltout => \c0.n2_adj_2341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_553_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__21916\,
            in1 => \N__18598\,
            in2 => \N__17106\,
            in3 => \N__17103\,
            lcout => \c0.n4_adj_2349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_550_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21504\,
            lcout => \c0.n10425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_708_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21503\,
            in1 => \N__18160\,
            in2 => \_gnd_net_\,
            in3 => \N__21203\,
            lcout => \c0.n10465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21204\,
            in1 => \N__18597\,
            in2 => \N__18162\,
            in3 => \N__21506\,
            lcout => n8_adj_2541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i3_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17740\,
            in2 => \_gnd_net_\,
            in3 => \N__19992\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49720\,
            ce => 'H',
            sr => \N__17349\
        );

    \c0.FRAME_MATCHER_state_i6_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17717\,
            in2 => \_gnd_net_\,
            in3 => \N__20055\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49707\,
            ce => 'H',
            sr => \N__17328\
        );

    \c0.FRAME_MATCHER_state_i5_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20371\,
            in2 => \_gnd_net_\,
            in3 => \N__20087\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \N__17340\
        );

    \c0.i1_2_lut_3_lut_adj_686_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__23338\,
            in1 => \_gnd_net_\,
            in2 => \N__25626\,
            in3 => \N__23445\,
            lcout => n242,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__19023\,
            in1 => \N__19005\,
            in2 => \_gnd_net_\,
            in3 => \N__17160\,
            lcout => n18_adj_2539,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_597_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21195\,
            in2 => \_gnd_net_\,
            in3 => \N__21453\,
            lcout => n10429,
            ltout => \n10429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_450_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__20982\,
            in1 => \N__18173\,
            in2 => \N__17163\,
            in3 => \N__20815\,
            lcout => n12965,
            ltout => \n12965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_827_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__18942\,
            in1 => \N__17154\,
            in2 => \N__17148\,
            in3 => \N__20983\,
            lcout => n15_adj_2540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__18174\,
            in2 => \N__17943\,
            in3 => \N__17139\,
            lcout => OPEN,
            ltout => \n21_adj_2538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__17130\,
            in1 => \N__18735\,
            in2 => \N__17124\,
            in3 => \N__17121\,
            lcout => \c0.FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_779_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__20981\,
            in1 => \N__23337\,
            in2 => \_gnd_net_\,
            in3 => \N__20814\,
            lcout => n8_adj_2498,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24565\,
            in2 => \_gnd_net_\,
            in3 => \N__19233\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49685\,
            ce => 'H',
            sr => \N__17448\
        );

    \c0.FRAME_MATCHER_i_i4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24586\,
            in2 => \_gnd_net_\,
            in3 => \N__19161\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49680\,
            ce => 'H',
            sr => \N__21552\
        );

    \c0.FRAME_MATCHER_i_i15_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24626\,
            in2 => \_gnd_net_\,
            in3 => \N__19602\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49675\,
            ce => 'H',
            sr => \N__17436\
        );

    \c0.FRAME_MATCHER_i_i17_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24627\,
            in2 => \_gnd_net_\,
            in3 => \N__19482\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49671\,
            ce => 'H',
            sr => \N__17427\
        );

    \c0.FRAME_MATCHER_i_i24_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24628\,
            in2 => \_gnd_net_\,
            in3 => \N__19770\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49668\,
            ce => 'H',
            sr => \N__17502\
        );

    \c0.FRAME_MATCHER_i_i22_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24629\,
            in2 => \_gnd_net_\,
            in3 => \N__19878\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \N__17490\
        );

    \c0.FRAME_MATCHER_state_i27_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17821\,
            in2 => \_gnd_net_\,
            in3 => \N__20495\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49798\,
            ce => 'H',
            sr => \N__17805\
        );

    \c0.FRAME_MATCHER_state_i14_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17632\,
            in2 => \_gnd_net_\,
            in3 => \N__20098\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49786\,
            ce => 'H',
            sr => \N__17187\
        );

    \c0.FRAME_MATCHER_state_i25_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17549\,
            in2 => \_gnd_net_\,
            in3 => \N__20097\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49770\,
            ce => 'H',
            sr => \N__17322\
        );

    \c0.FRAME_MATCHER_state_i13_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17575\,
            in2 => \_gnd_net_\,
            in3 => \N__20020\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49757\,
            ce => 'H',
            sr => \N__17193\
        );

    \c0.i1_2_lut_4_lut_adj_647_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18429\,
            in1 => \N__18027\,
            in2 => \N__17604\,
            in3 => \N__19136\,
            lcout => \c0.n17263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i10_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19990\,
            in2 => \_gnd_net_\,
            in3 => \N__17603\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49744\,
            ce => 'H',
            sr => \N__17283\
        );

    \c0.i1_2_lut_4_lut_adj_650_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18430\,
            in1 => \N__18028\,
            in2 => \N__17271\,
            in3 => \N__19137\,
            lcout => \c0.n17265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_657_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19138\,
            in1 => \N__17229\,
            in2 => \N__18058\,
            in3 => \N__18431\,
            lcout => \c0.n17267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_659_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18432\,
            in1 => \N__18032\,
            in2 => \N__17580\,
            in3 => \N__19139\,
            lcout => \c0.n17269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_663_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19140\,
            in1 => \N__17636\,
            in2 => \N__18059\,
            in3 => \N__18433\,
            lcout => \c0.n17303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_669_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18434\,
            in1 => \N__18036\,
            in2 => \N__17667\,
            in3 => \N__19141\,
            lcout => \c0.n17271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_673_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19142\,
            in1 => \N__20349\,
            in2 => \N__18060\,
            in3 => \N__18435\,
            lcout => \c0.n8_adj_2254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_548_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__19003\,
            in1 => \N__18888\,
            in2 => \N__18216\,
            in3 => \N__22567\,
            lcout => \c0.n17713\,
            ltout => \c0.n17713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_442_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__22569\,
            in1 => \N__20318\,
            in2 => \N__17364\,
            in3 => \N__18380\,
            lcout => \c0.n8_adj_2234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18379\,
            in1 => \N__18016\,
            in2 => \N__17748\,
            in3 => \N__22568\,
            lcout => \c0.n17281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_639_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19145\,
            in1 => \N__17689\,
            in2 => \N__18056\,
            in3 => \N__18383\,
            lcout => \c0.n8_adj_2258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_446_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18381\,
            in1 => \N__18017\,
            in2 => \N__20382\,
            in3 => \N__22570\,
            lcout => \c0.n17259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_638_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19144\,
            in1 => \N__17716\,
            in2 => \N__18055\,
            in3 => \N__18382\,
            lcout => \c0.n17261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11136_2_lut_4_lut_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18378\,
            in1 => \N__18015\,
            in2 => \N__17553\,
            in3 => \N__19143\,
            lcout => \c0.n13900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_640_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19146\,
            in1 => \N__17310\,
            in2 => \N__18057\,
            in3 => \N__18384\,
            lcout => \c0.n8_adj_2257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i7_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17690\,
            in2 => \_gnd_net_\,
            in3 => \N__20101\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49721\,
            ce => 'H',
            sr => \N__17397\
        );

    \c0.FRAME_MATCHER_state_i9_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18082\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49708\,
            ce => 'H',
            sr => \N__17955\
        );

    \c0.FRAME_MATCHER_i_i1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24502\,
            in2 => \_gnd_net_\,
            in3 => \N__19206\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \N__18282\
        );

    \c0.FRAME_MATCHER_i_i20_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19452\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49692\,
            ce => 'H',
            sr => \N__18108\
        );

    \c0.i14_4_lut_adj_607_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20229\,
            in1 => \N__22222\,
            in2 => \N__21046\,
            in3 => \N__19371\,
            lcout => OPEN,
            ltout => \c0.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17415\,
            in1 => \N__17382\,
            in2 => \N__17388\,
            in3 => \N__17376\,
            lcout => OPEN,
            ltout => \c0.n48_adj_2383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_612_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21947\,
            in1 => \N__17370\,
            in2 => \N__17385\,
            in3 => \N__22083\,
            lcout => \c0.n10522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_605_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19746\,
            in1 => \N__22439\,
            in2 => \N__22179\,
            in3 => \N__19851\,
            lcout => \c0.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_606_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19623\,
            in1 => \N__19513\,
            in2 => \N__24704\,
            in3 => \N__19317\,
            lcout => \c0.n41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_611_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21093\,
            in1 => \N__19566\,
            in2 => \N__24380\,
            in3 => \N__20751\,
            lcout => \c0.n43_adj_2384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i30_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24567\,
            in2 => \_gnd_net_\,
            in3 => \N__20271\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49681\,
            ce => 'H',
            sr => \N__17457\
        );

    \c0.select_284_Select_30_i3_2_lut_3_lut_4_lut_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__20752\,
            in2 => \N__21924\,
            in3 => \N__21670\,
            lcout => \c0.n3_adj_2281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_14_i3_2_lut_3_lut_4_lut_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21664\,
            in1 => \N__21902\,
            in2 => \N__21108\,
            in3 => \N__21516\,
            lcout => \c0.n3_adj_2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_13_i3_2_lut_3_lut_4_lut_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21515\,
            in1 => \N__24379\,
            in2 => \N__21922\,
            in3 => \N__21663\,
            lcout => \c0.n3_adj_2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_12_i3_2_lut_3_lut_4_lut_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__21903\,
            in2 => \N__22626\,
            in3 => \N__21517\,
            lcout => \c0.n3_adj_2322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_15_i3_2_lut_3_lut_4_lut_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21519\,
            in1 => \N__21669\,
            in2 => \N__21923\,
            in3 => \N__19630\,
            lcout => \c0.n3_adj_2311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_17_i3_2_lut_3_lut_4_lut_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19512\,
            in1 => \N__21904\,
            in2 => \N__21708\,
            in3 => \N__21518\,
            lcout => \c0.n3_adj_2307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_602_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19905\,
            in1 => \N__19797\,
            in2 => \N__20717\,
            in3 => \N__19407\,
            lcout => \c0.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i21_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19392\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49676\,
            ce => 'H',
            sr => \N__17406\
        );

    \c0.select_284_Select_21_i3_2_lut_3_lut_4_lut_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21531\,
            in1 => \N__19408\,
            in2 => \N__21715\,
            in3 => \N__21885\,
            lcout => \c0.n3_adj_2299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_24_i3_2_lut_3_lut_4_lut_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21881\,
            in1 => \N__21684\,
            in2 => \N__19805\,
            in3 => \N__21527\,
            lcout => \c0.n3_adj_2293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_22_i3_2_lut_3_lut_4_lut_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21528\,
            in1 => \N__19919\,
            in2 => \N__21713\,
            in3 => \N__21883\,
            lcout => \c0.n3_adj_2297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_29_i3_2_lut_3_lut_4_lut_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21886\,
            in1 => \N__20712\,
            in2 => \N__21543\,
            in3 => \N__21695\,
            lcout => \c0.n3_adj_2283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_10_i3_2_lut_3_lut_4_lut_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21530\,
            in1 => \N__22221\,
            in2 => \N__21714\,
            in3 => \N__21884\,
            lcout => \c0.n3_adj_2326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_11_i3_2_lut_3_lut_4_lut_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__21685\,
            in2 => \N__22071\,
            in3 => \N__21529\,
            lcout => \c0.n3_adj_2324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19701\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \N__18234\
        );

    \c0.FRAME_MATCHER_i_i10_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19251\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49669\,
            ce => 'H',
            sr => \N__17478\
        );

    \c0.FRAME_MATCHER_i_i14_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24625\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49667\,
            ce => 'H',
            sr => \N__17469\
        );

    \c0.FRAME_MATCHER_state_i30_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17782\,
            in2 => \_gnd_net_\,
            in3 => \N__20496\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49810\,
            ce => 'H',
            sr => \N__17760\
        );

    \c0.FRAME_MATCHER_state_i24_LC_3_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18506\,
            in2 => \_gnd_net_\,
            in3 => \N__20100\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49799\,
            ce => 'H',
            sr => \N__17847\
        );

    \c0.FRAME_MATCHER_state_i22_LC_3_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18683\,
            in2 => \_gnd_net_\,
            in3 => \N__20099\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49787\,
            ce => 'H',
            sr => \N__18663\
        );

    \c0.i20_4_lut_LC_3_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17747\,
            in1 => \N__17721\,
            in2 => \N__17697\,
            in3 => \N__20132\,
            lcout => OPEN,
            ltout => \c0.n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17610\,
            in1 => \N__17529\,
            in2 => \N__17670\,
            in3 => \N__17586\,
            lcout => \c0.n56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17666\,
            in1 => \N__18089\,
            in2 => \N__17643\,
            in3 => \N__18545\,
            lcout => \c0.n50_adj_2353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_3_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17912\,
            in1 => \N__17599\,
            in2 => \N__17834\,
            in3 => \N__17521\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_3_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17872\,
            in1 => \N__18679\,
            in2 => \N__17576\,
            in3 => \N__17545\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i23_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17523\,
            in2 => \_gnd_net_\,
            in3 => \N__20096\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49771\,
            ce => 'H',
            sr => \N__17511\
        );

    \c0.i1_2_lut_adj_497_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18705\,
            lcout => \c0.n17275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_697_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18422\,
            in1 => \N__18042\,
            in2 => \N__17877\,
            in3 => \N__19129\,
            lcout => \c0.n8_adj_2252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i17_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17876\,
            in2 => \_gnd_net_\,
            in3 => \N__20042\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49759\,
            ce => 'H',
            sr => \N__17859\
        );

    \c0.i1_2_lut_4_lut_adj_698_LC_3_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18423\,
            in1 => \N__18043\,
            in2 => \N__18510\,
            in3 => \N__19130\,
            lcout => \c0.n8_adj_2246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_720_LC_3_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19131\,
            in1 => \N__18546\,
            in2 => \N__18061\,
            in3 => \N__18424\,
            lcout => \c0.n8_adj_2245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_732_LC_3_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18425\,
            in1 => \N__18047\,
            in2 => \N__17835\,
            in3 => \N__19132\,
            lcout => \c0.n17277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_736_LC_3_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19133\,
            in1 => \N__18653\,
            in2 => \N__18062\,
            in3 => \N__18426\,
            lcout => \c0.n17299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_742_LC_3_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__18051\,
            in2 => \N__20406\,
            in3 => \N__19134\,
            lcout => \c0.n8_adj_2244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_745_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__19135\,
            in1 => \N__17792\,
            in2 => \N__18063\,
            in3 => \N__18428\,
            lcout => \c0.n17283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_749_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__18377\,
            in1 => \N__18040\,
            in2 => \N__17913\,
            in3 => \N__19088\,
            lcout => \c0.n17279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_451_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__30492\,
            in1 => \N__25052\,
            in2 => \N__29943\,
            in3 => \N__30114\,
            lcout => n17694,
            ltout => \n17694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_755_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__25053\,
            in1 => \N__46151\,
            in2 => \N__17916\,
            in3 => \N__33057\,
            lcout => \c0.n4_adj_2231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_765_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__33060\,
            in1 => \N__25056\,
            in2 => \N__25114\,
            in3 => \N__49107\,
            lcout => \c0.n4_adj_2216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_760_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__25054\,
            in1 => \N__25100\,
            in2 => \N__48570\,
            in3 => \N__33058\,
            lcout => \c0.n4_adj_2226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_761_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__33059\,
            in1 => \N__25055\,
            in2 => \N__25113\,
            in3 => \N__48017\,
            lcout => \c0.n4_adj_2225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i31_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__17911\,
            in1 => \_gnd_net_\,
            in2 => \N__20498\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49745\,
            ce => 'H',
            sr => \N__17892\
        );

    \c0.i1_2_lut_4_lut_adj_768_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__25057\,
            in2 => \N__25115\,
            in3 => \N__48928\,
            lcout => \c0.n4_adj_2204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10973_2_lut_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30011\,
            in2 => \_gnd_net_\,
            in3 => \N__19086\,
            lcout => OPEN,
            ltout => \FRAME_MATCHER_state_31_N_1406_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_829_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__17932\,
            in1 => \N__18925\,
            in2 => \N__17880\,
            in3 => \N__18798\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__24446\,
            in1 => \N__25099\,
            in2 => \N__28713\,
            in3 => \N__30518\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24447\,
            in2 => \_gnd_net_\,
            in3 => \N__19179\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49732\,
            ce => 'H',
            sr => \N__18270\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_625_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21197\,
            in1 => \N__21295\,
            in2 => \N__23342\,
            in3 => \N__21507\,
            lcout => \c0.n115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_718_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__19000\,
            in1 => \N__18924\,
            in2 => \_gnd_net_\,
            in3 => \N__18590\,
            lcout => n1166,
            ltout => \n1166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_588_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25098\,
            in2 => \N__18096\,
            in3 => \_gnd_net_\,
            lcout => \c0.n10497\,
            ltout => \c0.n10497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_644_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__19087\,
            in1 => \N__18093\,
            in2 => \N__18066\,
            in3 => \N__18041\,
            lcout => \c0.n17239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17936\,
            in1 => \N__20847\,
            in2 => \_gnd_net_\,
            in3 => \N__21535\,
            lcout => \c0.FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49722\,
            ce => 'H',
            sr => \N__18132\
        );

    \c0.rx.i1_2_lut_adj_398_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27999\,
            in2 => \_gnd_net_\,
            in3 => \N__27939\,
            lcout => \c0.rx.n57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15583_2_lut_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26975\,
            lcout => \c0.rx.n18304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_397_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27430\,
            in2 => \_gnd_net_\,
            in3 => \N__27940\,
            lcout => \c0.rx.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_421_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27941\,
            in1 => \_gnd_net_\,
            in2 => \N__27449\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.n167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_adj_413_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__34220\,
            in1 => \N__21951\,
            in2 => \_gnd_net_\,
            in3 => \N__24448\,
            lcout => \c0.rx.n12963\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_510_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__33237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21291\,
            lcout => n1437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_452_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__20843\,
            in1 => \N__18161\,
            in2 => \_gnd_net_\,
            in3 => \N__21454\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_455_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011101"
        )
    port map (
            in0 => \N__18730\,
            in1 => \N__18599\,
            in2 => \N__18135\,
            in3 => \N__18948\,
            lcout => \c0.n18907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_593_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__18600\,
            in1 => \N__18834\,
            in2 => \N__23336\,
            in3 => \N__19041\,
            lcout => OPEN,
            ltout => \n13_adj_2469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__18731\,
            in1 => \N__18189\,
            in2 => \N__18120\,
            in3 => \N__18117\,
            lcout => \c0.FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_31_i3_2_lut_3_lut_4_lut_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21711\,
            in1 => \N__21917\,
            in2 => \N__20985\,
            in3 => \N__21455\,
            lcout => \c0.n3_adj_2279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_20_i3_2_lut_3_lut_4_lut_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21712\,
            in1 => \N__21918\,
            in2 => \N__22026\,
            in3 => \N__21456\,
            lcout => \c0.n3_adj_2301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_716_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__20797\,
            in1 => \N__20952\,
            in2 => \N__18201\,
            in3 => \N__19001\,
            lcout => \c0.n2_adj_2315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_746_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23404\,
            in1 => \N__23295\,
            in2 => \N__20975\,
            in3 => \N__25598\,
            lcout => n15118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_614_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23402\,
            lcout => \c0.n232\,
            ltout => \c0.n232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_777_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__20950\,
            in1 => \N__23290\,
            in2 => \N__18219\,
            in3 => \N__20795\,
            lcout => \c0.n7528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i0_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24500\,
            in2 => \_gnd_net_\,
            in3 => \N__19215\,
            lcout => \c0.FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \N__18258\
        );

    \c0.i1_3_lut_4_lut_adj_634_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111111"
        )
    port map (
            in0 => \N__20951\,
            in1 => \N__23294\,
            in2 => \N__18818\,
            in3 => \N__20796\,
            lcout => \c0.n6_adj_2364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_578_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__25597\,
            in1 => \_gnd_net_\,
            in2 => \N__23331\,
            in3 => \N__23403\,
            lcout => n237,
            ltout => \n237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_828_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__19002\,
            in1 => \N__18833\,
            in2 => \N__18192\,
            in3 => \N__19040\,
            lcout => n22_adj_2465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10991_2_lut_3_lut_4_lut_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21196\,
            in1 => \N__21296\,
            in2 => \N__19577\,
            in3 => \N__21508\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19548\,
            in2 => \_gnd_net_\,
            in3 => \N__24499\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49693\,
            ce => 'H',
            sr => \N__18183\
        );

    \c0.select_284_Select_16_i3_2_lut_3_lut_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19573\,
            in1 => \N__21678\,
            in2 => \_gnd_net_\,
            in3 => \N__22571\,
            lcout => \c0.n3_adj_2309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_556_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__33142\,
            in1 => \N__18789\,
            in2 => \N__30043\,
            in3 => \N__24498\,
            lcout => \c0.n10353\,
            ltout => \c0.n10353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_18_i3_2_lut_3_lut_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__24699\,
            in1 => \_gnd_net_\,
            in2 => \N__18285\,
            in3 => \N__22572\,
            lcout => \c0.n3_adj_2305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_596_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21511\,
            in1 => \N__25659\,
            in2 => \N__21710\,
            in3 => \N__21914\,
            lcout => \c0.n3_adj_2345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_598_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21912\,
            in1 => \N__21671\,
            in2 => \N__23335\,
            in3 => \N__21510\,
            lcout => \c0.n3_adj_2343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_627_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21509\,
            in1 => \N__23427\,
            in2 => \N__21709\,
            in3 => \N__21913\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_23_i3_2_lut_3_lut_4_lut_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19854\,
            in1 => \N__21897\,
            in2 => \N__21699\,
            in3 => \N__21525\,
            lcout => \c0.n3_adj_2295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i23_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24501\,
            in2 => \_gnd_net_\,
            in3 => \N__19830\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \N__18246\
        );

    \c0.i10982_2_lut_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19853\,
            in2 => \_gnd_net_\,
            in3 => \N__22566\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_25_i3_2_lut_3_lut_4_lut_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21521\,
            in1 => \N__21647\,
            in2 => \N__21919\,
            in3 => \N__19749\,
            lcout => \c0.n3_adj_2291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_26_i3_2_lut_3_lut_4_lut_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22438\,
            in1 => \N__21898\,
            in2 => \N__21700\,
            in3 => \N__21526\,
            lcout => \c0.n3_adj_2289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_27_i3_2_lut_3_lut_4_lut_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21524\,
            in1 => \N__22397\,
            in2 => \N__21921\,
            in3 => \N__21649\,
            lcout => \c0.n3_adj_2287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_28_i3_2_lut_3_lut_4_lut_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21646\,
            in1 => \N__21887\,
            in2 => \N__22287\,
            in3 => \N__21522\,
            lcout => \c0.n3_adj_2285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_6_i3_2_lut_3_lut_4_lut_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21523\,
            in1 => \N__22178\,
            in2 => \N__21920\,
            in3 => \N__21648\,
            lcout => \c0.n3_adj_2334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i26_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24566\,
            in2 => \_gnd_net_\,
            in3 => \N__19689\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49682\,
            ce => 'H',
            sr => \N__18321\
        );

    \c0.FRAME_MATCHER_i_i29_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24568\,
            in2 => \_gnd_net_\,
            in3 => \N__19674\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49677\,
            ce => 'H',
            sr => \N__18315\
        );

    \c0.FRAME_MATCHER_i_i8_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24621\,
            in2 => \_gnd_net_\,
            in3 => \N__19278\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \N__18852\
        );

    \c0.FRAME_MATCHER_i_i31_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24622\,
            in2 => \_gnd_net_\,
            in3 => \N__20253\,
            lcout => \FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49670\,
            ce => 'H',
            sr => \N__18309\
        );

    \c0.FRAME_MATCHER_i_i19_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24624\,
            in2 => \_gnd_net_\,
            in3 => \N__19467\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \N__18297\
        );

    \c0.select_284_Select_19_i3_2_lut_3_lut_4_lut_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21698\,
            in1 => \N__21911\,
            in2 => \N__21036\,
            in3 => \N__21542\,
            lcout => \c0.n3_adj_2303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.PHASES_i2_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__35639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35411\,
            lcout => \PIN_2_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49758\,
            ce => \N__20163\,
            sr => \N__35352\
        );

    \c0.FRAME_MATCHER_state_i26_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18544\,
            in2 => \_gnd_net_\,
            in3 => \N__20497\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49823\,
            ce => 'H',
            sr => \N__18522\
        );

    \c0.FRAME_MATCHER_state_i21_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18464\,
            in2 => \_gnd_net_\,
            in3 => \N__20089\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49811\,
            ce => 'H',
            sr => \N__18447\
        );

    \c0.i17_4_lut_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18502\,
            in1 => \N__18652\,
            in2 => \N__18465\,
            in3 => \N__18484\,
            lcout => \c0.n46_adj_2356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i18_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20092\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49800\,
            ce => 'H',
            sr => \N__18474\
        );

    \c0.i1_2_lut_adj_473_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18485\,
            in2 => \_gnd_net_\,
            in3 => \N__18703\,
            lcout => \c0.n17293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_480_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18702\,
            in1 => \N__18463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n8_adj_2247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_475_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20136\,
            in2 => \_gnd_net_\,
            in3 => \N__18701\,
            lcout => \c0.n8_adj_2250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_491_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111001100"
        )
    port map (
            in0 => \N__18421\,
            in1 => \N__18887\,
            in2 => \N__18336\,
            in3 => \N__19119\,
            lcout => \c0.n8_adj_2273\,
            ltout => \c0.n8_adj_2273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_477_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18708\,
            in3 => \N__20423\,
            lcout => \c0.n8_adj_2249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_488_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18684\,
            lcout => \c0.n17273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i28_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18654\,
            in2 => \_gnd_net_\,
            in3 => \N__20491\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49788\,
            ce => 'H',
            sr => \N__18636\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_791_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__33180\,
            in1 => \N__33263\,
            in2 => \N__30044\,
            in3 => \N__30108\,
            lcout => \c0.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18630\,
            in1 => \N__20286\,
            in2 => \N__18621\,
            in3 => \N__18609\,
            lcout => \c0.n10513\,
            ltout => \c0.n10513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_804_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33179\,
            in1 => \N__30034\,
            in2 => \N__18603\,
            in3 => \N__33264\,
            lcout => \FRAME_MATCHER_i_31__N_1275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_547_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__30110\,
            in1 => \N__30022\,
            in2 => \N__33282\,
            in3 => \N__33182\,
            lcout => \c0.n6033\,
            ltout => \c0.n6033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i7_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__28814\,
            in1 => \N__28935\,
            in2 => \N__18561\,
            in3 => \N__28836\,
            lcout => \c0.data_out_frame2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_799_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30109\,
            in1 => \N__30021\,
            in2 => \N__33281\,
            in3 => \N__33181\,
            lcout => \FRAME_MATCHER_i_31__N_1272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1014_2_lut_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23132\,
            in2 => \_gnd_net_\,
            in3 => \N__25914\,
            lcout => \c0.n2126\,
            ltout => \c0.n2126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_509_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111011"
        )
    port map (
            in0 => \N__23679\,
            in1 => \N__22931\,
            in2 => \N__18753\,
            in3 => \N__20277\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30112\,
            in1 => \N__33170\,
            in2 => \N__33277\,
            in3 => \N__30007\,
            lcout => \FRAME_MATCHER_i_31__N_1273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_616_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33169\,
            in1 => \N__33255\,
            in2 => \N__30035\,
            in3 => \N__30111\,
            lcout => \FRAME_MATCHER_i_31__N_1270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_469_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__26008\,
            in1 => \N__23083\,
            in2 => \N__23520\,
            in3 => \N__26043\,
            lcout => OPEN,
            ltout => \c0.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__18750\,
            in1 => \N__26307\,
            in2 => \N__18744\,
            in3 => \N__25952\,
            lcout => OPEN,
            ltout => \c0.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26262\,
            in1 => \N__18714\,
            in2 => \N__18741\,
            in3 => \N__18774\,
            lcout => \c0.n50\,
            ltout => \c0.n50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11086_2_lut_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25058\,
            in2 => \N__18738\,
            in3 => \_gnd_net_\,
            lcout => n13849,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_519_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__20574\,
            in1 => \N__25443\,
            in2 => \N__22652\,
            in3 => \N__20607\,
            lcout => \c0.n19_adj_2351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_714_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33259\,
            in2 => \_gnd_net_\,
            in3 => \N__30113\,
            lcout => \c0.n10346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22747\,
            in1 => \N__30724\,
            in2 => \_gnd_net_\,
            in3 => \N__30306\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26002\,
            in1 => \N__23591\,
            in2 => \_gnd_net_\,
            in3 => \N__24155\,
            lcout => data_in_frame_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27621\,
            in1 => \N__20546\,
            in2 => \_gnd_net_\,
            in3 => \N__23635\,
            lcout => data_in_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_514_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__26133\,
            in1 => \N__23107\,
            in2 => \N__20592\,
            in3 => \N__23082\,
            lcout => OPEN,
            ltout => \c0.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_521_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111111"
        )
    port map (
            in0 => \N__23556\,
            in1 => \N__23180\,
            in2 => \N__18777\,
            in3 => \N__22989\,
            lcout => \c0.n25_adj_2352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15103_3_lut_4_lut_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__20590\,
            in1 => \N__25998\,
            in2 => \N__20573\,
            in3 => \N__25913\,
            lcout => OPEN,
            ltout => \c0.n17962_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_695_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__26394\,
            in1 => \N__23181\,
            in2 => \N__18768\,
            in3 => \N__26079\,
            lcout => \c0.n24_adj_2418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i1_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25011\,
            in1 => \N__48286\,
            in2 => \N__30663\,
            in3 => \N__30519\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49733\,
            ce => 'H',
            sr => \N__18765\
        );

    \c0.tx2.i15302_3_lut_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33941\,
            in1 => \N__28512\,
            in2 => \_gnd_net_\,
            in3 => \N__48840\,
            lcout => \c0.tx2.n18163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15303_3_lut_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28548\,
            in1 => \N__33942\,
            in2 => \_gnd_net_\,
            in3 => \N__42993\,
            lcout => \c0.tx2.n18164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__29094\,
            in1 => \N__29070\,
            in2 => \_gnd_net_\,
            in3 => \N__29043\,
            lcout => \c0.tx2.n12769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10981_2_lut_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19809\,
            in2 => \_gnd_net_\,
            in3 => \N__22501\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10983_2_lut_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22502\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19920\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10984_2_lut_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22503\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10992_2_lut_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19638\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_576_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21163\,
            in1 => \N__21254\,
            in2 => \_gnd_net_\,
            in3 => \N__21373\,
            lcout => \c0.n9575\,
            ltout => \c0.n9575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_575_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29982\,
            in2 => \N__18837\,
            in3 => \N__20816\,
            lcout => n12999,
            ltout => \n12999_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_591_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__18822\,
            in1 => \N__23356\,
            in2 => \N__18801\,
            in3 => \N__19039\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_571_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__20976\,
            in1 => \N__29983\,
            in2 => \_gnd_net_\,
            in3 => \N__19066\,
            lcout => n12966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10989_2_lut_3_lut_4_lut_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21164\,
            in1 => \N__21255\,
            in2 => \N__19524\,
            in3 => \N__21374\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_449_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21375\,
            in1 => \N__18941\,
            in2 => \N__18906\,
            in3 => \N__20836\,
            lcout => OPEN,
            ltout => \c0.n16685_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_453_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__19016\,
            in1 => \N__19004\,
            in2 => \N__18951\,
            in3 => \N__20775\,
            lcout => \c0.n6_adj_2267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i57_3_lut_4_lut_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21372\,
            in1 => \N__18940\,
            in2 => \N__18905\,
            in3 => \N__21788\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_7_i3_2_lut_3_lut_4_lut_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__21811\,
            in2 => \N__21697\,
            in3 => \N__21423\,
            lcout => \c0.n3_adj_2332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i7_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24533\,
            in2 => \_gnd_net_\,
            in3 => \N__19341\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \N__18864\
        );

    \c0.i11000_2_lut_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19366\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_8_i3_2_lut_3_lut_4_lut_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__21639\,
            in2 => \N__21870\,
            in3 => \N__19322\,
            lcout => \c0.n3_adj_2330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_9_i3_2_lut_3_lut_4_lut_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20234\,
            in1 => \N__21810\,
            in2 => \N__21696\,
            in3 => \N__21422\,
            lcout => \c0.n3_adj_2328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10998_2_lut_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20233\,
            in2 => \_gnd_net_\,
            in3 => \N__22498\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10999_2_lut_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19323\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10980_2_lut_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19747\,
            in2 => \_gnd_net_\,
            in3 => \N__22497\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_2_lut_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22116\,
            in1 => \N__23401\,
            in2 => \N__23853\,
            in3 => \N__19209\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_0\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \c0.n16486\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_3_lut_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__21117\,
            in1 => \N__25647\,
            in2 => \N__23856\,
            in3 => \N__19194\,
            lcout => \c0.n27_adj_2426\,
            ltout => OPEN,
            carryin => \c0.n16486\,
            carryout => \c0.n16487\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_4_lut_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19191\,
            in1 => \N__23790\,
            in2 => \N__23366\,
            in3 => \N__19167\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \c0.n16487\,
            carryout => \c0.n16488\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_5_lut_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20859\,
            in1 => \N__22344\,
            in2 => \N__23857\,
            in3 => \N__19164\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_3\,
            ltout => OPEN,
            carryin => \c0.n16488\,
            carryout => \c0.n16489\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_6_lut_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__21930\,
            in1 => \N__21746\,
            in2 => \N__23854\,
            in3 => \N__19152\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_4\,
            ltout => OPEN,
            carryin => \c0.n16489\,
            carryout => \c0.n16490\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_7_lut_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20868\,
            in1 => \N__21971\,
            in2 => \N__23858\,
            in3 => \N__19149\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_5\,
            ltout => OPEN,
            carryin => \c0.n16490\,
            carryout => \c0.n16491\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_8_lut_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22128\,
            in1 => \N__22158\,
            in2 => \N__23855\,
            in3 => \N__19380\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_6\,
            ltout => OPEN,
            carryin => \c0.n16491\,
            carryout => \c0.n16492\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_9_lut_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19377\,
            in1 => \N__19365\,
            in2 => \N__23859\,
            in3 => \N__19335\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_7\,
            ltout => OPEN,
            carryin => \c0.n16492\,
            carryout => \c0.n16493\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_10_lut_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__19318\,
            in2 => \N__23906\,
            in3 => \N__19266\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_8\,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \c0.n16494\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_11_lut_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19263\,
            in1 => \N__23863\,
            in2 => \N__20235\,
            in3 => \N__19254\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_9\,
            ltout => OPEN,
            carryin => \c0.n16494\,
            carryout => \c0.n16495\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_12_lut_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22188\,
            in1 => \N__22223\,
            in2 => \N__23907\,
            in3 => \N__19239\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_10\,
            ltout => OPEN,
            carryin => \c0.n16495\,
            carryout => \c0.n16496\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_13_lut_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__22038\,
            in1 => \N__23867\,
            in2 => \N__22070\,
            in3 => \N__19236\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_11\,
            ltout => OPEN,
            carryin => \c0.n16496\,
            carryout => \c0.n16497\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_14_lut_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22584\,
            in1 => \N__22618\,
            in2 => \N__23908\,
            in3 => \N__19221\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_12\,
            ltout => OPEN,
            carryin => \c0.n16497\,
            carryout => \c0.n16498\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_15_lut_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__22233\,
            in1 => \N__23871\,
            in2 => \N__24381\,
            in3 => \N__19218\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_13\,
            ltout => OPEN,
            carryin => \c0.n16498\,
            carryout => \c0.n16499\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_16_lut_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__21103\,
            in2 => \N__23909\,
            in3 => \N__19653\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_14\,
            ltout => OPEN,
            carryin => \c0.n16499\,
            carryout => \c0.n16500\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_17_lut_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19650\,
            in1 => \N__23875\,
            in2 => \N__19637\,
            in3 => \N__19593\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_15\,
            ltout => OPEN,
            carryin => \c0.n16500\,
            carryout => \c0.n16501\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_18_lut_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19590\,
            in1 => \N__23877\,
            in2 => \N__19581\,
            in3 => \N__19539\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_16\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \c0.n16502\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_19_lut_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19536\,
            in1 => \N__23881\,
            in2 => \N__19520\,
            in3 => \N__19473\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_17\,
            ltout => OPEN,
            carryin => \c0.n16502\,
            carryout => \c0.n16503\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_20_lut_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20880\,
            in1 => \N__24703\,
            in2 => \N__23911\,
            in3 => \N__19470\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_18\,
            ltout => OPEN,
            carryin => \c0.n16503\,
            carryout => \c0.n16504\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_21_lut_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20997\,
            in1 => \N__23885\,
            in2 => \N__21048\,
            in3 => \N__19455\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_19\,
            ltout => OPEN,
            carryin => \c0.n16504\,
            carryout => \c0.n16505\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_22_lut_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__21999\,
            in1 => \N__23876\,
            in2 => \N__22032\,
            in3 => \N__19440\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_20\,
            ltout => OPEN,
            carryin => \c0.n16505\,
            carryout => \c0.n16506\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_23_lut_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19437\,
            in1 => \N__23886\,
            in2 => \N__19421\,
            in3 => \N__19383\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_21\,
            ltout => OPEN,
            carryin => \c0.n16506\,
            carryout => \c0.n16507\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_24_lut_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19932\,
            in1 => \N__19915\,
            in2 => \N__23912\,
            in3 => \N__19866\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_22\,
            ltout => OPEN,
            carryin => \c0.n16507\,
            carryout => \c0.n16508\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_25_lut_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19863\,
            in1 => \N__19852\,
            in2 => \N__23910\,
            in3 => \N__19824\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_23\,
            ltout => OPEN,
            carryin => \c0.n16508\,
            carryout => \c0.n16509\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_26_lut_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19821\,
            in1 => \N__19804\,
            in2 => \N__23913\,
            in3 => \N__19761\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_24\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \c0.n16510\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_27_lut_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19758\,
            in1 => \N__23893\,
            in2 => \N__19748\,
            in3 => \N__19692\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_25\,
            ltout => OPEN,
            carryin => \c0.n16510\,
            carryout => \c0.n16511\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_28_lut_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22410\,
            in1 => \N__22434\,
            in2 => \N__23914\,
            in3 => \N__19683\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_26\,
            ltout => OPEN,
            carryin => \c0.n16511\,
            carryout => \c0.n16512\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_29_lut_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__22578\,
            in1 => \N__23897\,
            in2 => \N__22398\,
            in3 => \N__19680\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_27\,
            ltout => OPEN,
            carryin => \c0.n16512\,
            carryout => \c0.n16513\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_30_lut_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__21060\,
            in1 => \N__23901\,
            in2 => \N__22283\,
            in3 => \N__19677\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_28\,
            ltout => OPEN,
            carryin => \c0.n16513\,
            carryout => \c0.n16514\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_31_lut_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20682\,
            in1 => \N__20716\,
            in2 => \N__23916\,
            in3 => \N__19668\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_29\,
            ltout => OPEN,
            carryin => \c0.n16514\,
            carryout => \c0.n16515\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_32_lut_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20733\,
            in1 => \N__20766\,
            in2 => \N__23915\,
            in3 => \N__20259\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_30\,
            ltout => OPEN,
            carryin => \c0.n16515\,
            carryout => \c0.n16516\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_33_lut_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__23905\,
            in1 => \N__20949\,
            in2 => \N__20898\,
            in3 => \N__20256\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i9_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20244\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49678\,
            ce => 'H',
            sr => \N__20199\
        );

    \c0.FRAME_MATCHER_i_i6_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20184\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \N__20175\
        );

    \control.i3_4_lut_4_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111110"
        )
    port map (
            in0 => \N__35675\,
            in1 => \N__35546\,
            in2 => \N__35454\,
            in3 => \N__35351\,
            lcout => \control.n18909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i16_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20341\,
            in2 => \_gnd_net_\,
            in3 => \N__20103\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__20151\
        );

    \c0.FRAME_MATCHER_state_i19_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20125\,
            in2 => \_gnd_net_\,
            in3 => \N__20090\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => 'H',
            sr => \N__20109\
        );

    \c0.FRAME_MATCHER_state_i20_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20424\,
            in2 => \_gnd_net_\,
            in3 => \N__20088\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49812\,
            ce => 'H',
            sr => \N__20508\
        );

    \c0.FRAME_MATCHER_state_i29_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20499\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => 'H',
            sr => \N__20436\
        );

    \c0.i1_2_lut_adj_525_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20422\,
            in2 => \_gnd_net_\,
            in3 => \N__20395\,
            lcout => OPEN,
            ltout => \c0.n30_adj_2355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20378\,
            in1 => \N__20342\,
            in2 => \N__20322\,
            in3 => \N__20319\,
            lcout => \c0.n51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_554_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__25335\,
            in2 => \N__22932\,
            in3 => \N__23022\,
            lcout => \c0.n16863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_447_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23021\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20663\,
            lcout => OPEN,
            ltout => \c0.n10613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_701_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__25392\,
            in1 => \N__22869\,
            in2 => \N__20280\,
            in3 => \N__25435\,
            lcout => \c0.n21_adj_2421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011101111011"
        )
    port map (
            in0 => \N__23020\,
            in1 => \N__25479\,
            in2 => \N__22691\,
            in3 => \N__20662\,
            lcout => \c0.n22_adj_2346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1010_2_lut_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23163\,
            in2 => \_gnd_net_\,
            in3 => \N__26175\,
            lcout => \c0.n2122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__25671\,
            in1 => \N__20531\,
            in2 => \N__26642\,
            in3 => \N__25548\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_655_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011111111"
        )
    port map (
            in0 => \N__22981\,
            in1 => \N__25953\,
            in2 => \N__20550\,
            in3 => \N__22938\,
            lcout => \c0.n19_adj_2400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26633\,
            in1 => \N__22950\,
            in2 => \_gnd_net_\,
            in3 => \N__25864\,
            lcout => data_in_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__25549\,
            in1 => \N__25673\,
            in2 => \N__20625\,
            in3 => \N__27096\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__28011\,
            in1 => \N__27372\,
            in2 => \N__26474\,
            in3 => \N__26823\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__25547\,
            in1 => \N__25672\,
            in2 => \N__24180\,
            in3 => \N__23519\,
            lcout => \c0.data_in_frame_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__28010\,
            in1 => \N__27371\,
            in2 => \N__27110\,
            in3 => \N__25802\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_692_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__22851\,
            in2 => \N__20532\,
            in3 => \N__23084\,
            lcout => \c0.n18_adj_2417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27217\,
            in1 => \N__26321\,
            in2 => \_gnd_net_\,
            in3 => \N__23637\,
            lcout => data_in_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_653_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__20520\,
            in1 => \N__23051\,
            in2 => \N__25377\,
            in3 => \N__26132\,
            lcout => \c0.n18_adj_2398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26638\,
            in1 => \N__23012\,
            in2 => \_gnd_net_\,
            in3 => \N__23587\,
            lcout => data_in_frame_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__23588\,
            in1 => \N__27218\,
            in2 => \N__23139\,
            in3 => \_gnd_net_\,
            lcout => data_in_frame_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_691_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__23555\,
            in2 => \N__20624\,
            in3 => \N__20606\,
            lcout => \c0.n15_adj_2416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_748_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25994\,
            in1 => \N__25902\,
            in2 => \_gnd_net_\,
            in3 => \N__23040\,
            lcout => \c0.n2137_adj_2237\,
            ltout => \c0.n2137_adj_2237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1026_2_lut_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20595\,
            in3 => \N__23011\,
            lcout => \c0.n2138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31910\,
            in1 => \N__46065\,
            in2 => \_gnd_net_\,
            in3 => \N__44057\,
            lcout => \c0.n5_adj_2197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26624\,
            in1 => \N__20591\,
            in2 => \_gnd_net_\,
            in3 => \N__26421\,
            lcout => data_in_frame_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26422\,
            in1 => \_gnd_net_\,
            in2 => \N__27205\,
            in3 => \N__20572\,
            lcout => data_in_frame_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27620\,
            in1 => \N__23109\,
            in2 => \_gnd_net_\,
            in3 => \N__26423\,
            lcout => data_in_frame_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_adj_405_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23221\,
            in1 => \N__25670\,
            in2 => \N__23349\,
            in3 => \N__23462\,
            lcout => n16802,
            ltout => \n16802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23158\,
            in1 => \_gnd_net_\,
            in2 => \N__20670\,
            in3 => \N__26495\,
            lcout => data_in_frame_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_444_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26191\,
            in2 => \_gnd_net_\,
            in3 => \N__20653\,
            lcout => \c0.n10569\,
            ltout => \c0.n10569_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_445_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23157\,
            in1 => \N__26163\,
            in2 => \N__20667\,
            in3 => \N__23130\,
            lcout => \c0.n17813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27111\,
            in1 => \N__23586\,
            in2 => \_gnd_net_\,
            in3 => \N__20654\,
            lcout => data_in_frame_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__26343\,
            in1 => \N__27993\,
            in2 => \N__24165\,
            in3 => \N__26358\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27112\,
            in1 => \N__22645\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => data_in_frame_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26496\,
            in1 => \N__25826\,
            in2 => \_gnd_net_\,
            in3 => \N__23625\,
            lcout => data_in_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20640\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_410_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27853\,
            in1 => \N__26870\,
            in2 => \_gnd_net_\,
            in3 => \N__26976\,
            lcout => n12600,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_adj_406_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25678\,
            in1 => \N__23453\,
            in2 => \N__23362\,
            in3 => \N__23210\,
            lcout => n11058,
            ltout => \n11058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26628\,
            in1 => \_gnd_net_\,
            in2 => \N__20862\,
            in3 => \N__26222\,
            lcout => data_in_frame_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26725\,
            in1 => \N__22684\,
            in2 => \_gnd_net_\,
            in3 => \N__26427\,
            lcout => data_in_frame_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_623_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__26550\,
            in1 => \N__23922\,
            in2 => \N__23976\,
            in3 => \N__23982\,
            lcout => n63,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_809_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22336\,
            in2 => \_gnd_net_\,
            in3 => \N__22493\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__33178\,
            in1 => \N__21165\,
            in2 => \_gnd_net_\,
            in3 => \N__21253\,
            lcout => \c0.n1502\,
            ltout => \c0.n1502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_454_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__21371\,
            in1 => \N__20977\,
            in2 => \N__20820\,
            in3 => \N__20817\,
            lcout => \c0.n4_adj_2266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_561_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21169\,
            in1 => \N__21252\,
            in2 => \_gnd_net_\,
            in3 => \N__21370\,
            lcout => \c0.n13033\,
            ltout => \c0.n13033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10975_2_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20769\,
            in3 => \N__20765\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10976_2_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20721\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10977_2_lut_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22282\,
            in2 => \_gnd_net_\,
            in3 => \N__22495\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10986_2_lut_3_lut_4_lut_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21396\,
            in1 => \N__21047\,
            in2 => \N__21289\,
            in3 => \N__21168\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_763_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20984\,
            in2 => \_gnd_net_\,
            in3 => \N__22496\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27121\,
            in1 => \N__25349\,
            in2 => \_gnd_net_\,
            in3 => \N__23636\,
            lcout => data_in_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_609_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23715\,
            in1 => \N__24027\,
            in2 => \N__24054\,
            in3 => \N__24006\,
            lcout => n63_adj_2534,
            ltout => \n63_adj_2534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10988_2_lut_3_lut_4_lut_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21397\,
            in1 => \N__21272\,
            in2 => \N__20883\,
            in3 => \N__24705\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23714\,
            in1 => \N__24015\,
            in2 => \_gnd_net_\,
            in3 => \N__26919\,
            lcout => \c0.n63_adj_2262\,
            ltout => \c0.n63_adj_2262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4650_2_lut_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20871\,
            in3 => \N__21166\,
            lcout => \c0.n7199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_515_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21167\,
            in1 => \N__21398\,
            in2 => \N__21978\,
            in3 => \N__21271\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24599\,
            in2 => \_gnd_net_\,
            in3 => \N__21993\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49711\,
            ce => 'H',
            sr => \N__21987\
        );

    \c0.select_284_Select_5_i3_2_lut_3_lut_4_lut_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21814\,
            in1 => \N__21970\,
            in2 => \N__21717\,
            in3 => \N__21452\,
            lcout => \c0.n3_adj_2336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_599_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__21969\,
            in1 => \N__21735\,
            in2 => \_gnd_net_\,
            in3 => \N__22335\,
            lcout => \c0.n10_adj_2378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_524_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21173\,
            in1 => \N__21276\,
            in2 => \N__21745\,
            in3 => \N__21449\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_3_i3_2_lut_3_lut_4_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21450\,
            in1 => \N__21701\,
            in2 => \N__22343\,
            in3 => \N__21812\,
            lcout => \c0.n3_adj_2340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_284_Select_4_i3_2_lut_3_lut_4_lut_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21813\,
            in1 => \N__21747\,
            in2 => \N__21716\,
            in3 => \N__21451\,
            lcout => \c0.n3_adj_2338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_560_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21448\,
            in1 => \N__25648\,
            in2 => \N__21290\,
            in3 => \N__21174\,
            lcout => \c0.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__0__2184_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32412\,
            in1 => \N__36993\,
            in2 => \_gnd_net_\,
            in3 => \N__37407\,
            lcout => \c0.data_out_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49701\,
            ce => \N__46845\,
            sr => \_gnd_net_\
        );

    \c0.i10993_2_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21104\,
            in2 => \_gnd_net_\,
            in3 => \N__22528\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10994_2_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10997_2_lut_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22224\,
            in2 => \_gnd_net_\,
            in3 => \N__22530\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11001_2_lut_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22168\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_724_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23446\,
            in2 => \_gnd_net_\,
            in3 => \N__22532\,
            lcout => \c0.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i11_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24630\,
            in2 => \_gnd_net_\,
            in3 => \N__22104\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49694\,
            ce => 'H',
            sr => \N__22098\
        );

    \c0.i1_2_lut_adj_600_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__22383\,
            in1 => \N__22056\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n26_adj_2379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_608_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22275\,
            in1 => \N__22617\,
            in2 => \N__22086\,
            in3 => \N__22027\,
            lcout => \c0.n44_adj_2382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10996_2_lut_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22565\,
            in1 => \N__22057\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10985_2_lut_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22028\,
            in2 => \_gnd_net_\,
            in3 => \N__22563\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10995_2_lut_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22619\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10978_2_lut_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22384\,
            in2 => \_gnd_net_\,
            in3 => \N__22561\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10979_2_lut_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22440\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i27_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24631\,
            in2 => \_gnd_net_\,
            in3 => \N__22404\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \N__22368\
        );

    \c0.FRAME_MATCHER_i_i3_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24633\,
            in2 => \_gnd_net_\,
            in3 => \N__22356\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49683\,
            ce => 'H',
            sr => \N__22308\
        );

    \c0.FRAME_MATCHER_i_i28_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22296\,
            in2 => \_gnd_net_\,
            in3 => \N__24644\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49679\,
            ce => 'H',
            sr => \N__22248\
        );

    \i15182_4_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100000"
        )
    port map (
            in0 => \N__24983\,
            in1 => \N__24944\,
            in2 => \N__24966\,
            in3 => \N__24824\,
            lcout => n18043,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15183_4_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011101100"
        )
    port map (
            in0 => \N__24945\,
            in1 => \N__24965\,
            in2 => \N__24828\,
            in3 => \N__24984\,
            lcout => n18044,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15184_3_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__22821\,
            in1 => \N__22815\,
            in2 => \_gnd_net_\,
            in3 => \N__24924\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.PHASES_i3_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__35656\,
            in1 => \N__35461\,
            in2 => \_gnd_net_\,
            in3 => \N__35511\,
            lcout => \PIN_3_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49773\,
            ce => \N__24912\,
            sr => \N__35347\
        );

    \c0.byte_transmit_counter2_i7_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25164\,
            in1 => \N__25225\,
            in2 => \N__30658\,
            in3 => \N__30555\,
            lcout => \c0.byte_transmit_counter2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49842\,
            ce => 'H',
            sr => \N__25026\
        );

    \c0.byte_transmit_counter2_i2_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__24993\,
            in1 => \N__47981\,
            in2 => \N__30657\,
            in3 => \N__30547\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \N__22785\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i3_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25317\,
            in1 => \N__49027\,
            in2 => \N__30643\,
            in3 => \N__30546\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49825\,
            ce => 'H',
            sr => \N__22722\
        );

    \c0.data_in_frame_0__i50_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27106\,
            in1 => \N__22835\,
            in2 => \_gnd_net_\,
            in3 => \N__25860\,
            lcout => data_in_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__22706\,
            in1 => \N__25706\,
            in2 => \N__25785\,
            in3 => \N__25550\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_700_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111101"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__22662\,
            in2 => \N__22656\,
            in3 => \N__26013\,
            lcout => OPEN,
            ltout => \c0.n23_adj_2420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_703_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22893\,
            in1 => \N__22887\,
            in2 => \N__22875\,
            in3 => \N__23061\,
            lcout => \c0.n4494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_adj_412_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__25705\,
            in1 => \N__23466\,
            in2 => \N__23367\,
            in3 => \N__23226\,
            lcout => n16797,
            ltout => \n16797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27211\,
            in1 => \_gnd_net_\,
            in2 => \N__22872\,
            in3 => \N__25416\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__25551\,
            in1 => \N__27212\,
            in2 => \N__25716\,
            in3 => \N__22868\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25861\,
            in1 => \N__25784\,
            in2 => \_gnd_net_\,
            in3 => \N__23537\,
            lcout => data_in_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__25546\,
            in1 => \N__25713\,
            in2 => \N__27627\,
            in3 => \N__22927\,
            lcout => \c0.data_in_frame_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__23461\,
            in1 => \N__23360\,
            in2 => \_gnd_net_\,
            in3 => \N__23220\,
            lcout => \c0.rx.n129\,
            ltout => \c0.rx.n129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__22850\,
            in1 => \N__25715\,
            in2 => \N__22854\,
            in3 => \N__24178\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__25712\,
            in1 => \N__26303\,
            in2 => \N__25782\,
            in3 => \N__25544\,
            lcout => \c0.data_in_frame_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_642_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22977\,
            in1 => \N__22926\,
            in2 => \N__22836\,
            in3 => \N__23028\,
            lcout => \c0.n16994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__25711\,
            in1 => \N__25477\,
            in2 => \N__26727\,
            in3 => \N__25543\,
            lcout => \c0.data_in_frame_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__25545\,
            in1 => \N__27216\,
            in2 => \N__22985\,
            in3 => \N__25714\,
            lcout => \c0.data_in_frame_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24177\,
            in1 => \N__23052\,
            in2 => \_gnd_net_\,
            in3 => \N__25863\,
            lcout => data_in_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_628_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23039\,
            in1 => \N__26297\,
            in2 => \N__25478\,
            in3 => \N__25872\,
            lcout => \c0.n10761\,
            ltout => \c0.n10761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_629_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23010\,
            in2 => \N__22992\,
            in3 => \N__23514\,
            lcout => \c0.n17733\,
            ltout => \c0.n17733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_632_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22976\,
            in2 => \N__22953\,
            in3 => \N__22949\,
            lcout => \c0.n17735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_641_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23481\,
            in1 => \N__26068\,
            in2 => \_gnd_net_\,
            in3 => \N__26042\,
            lcout => \c0.n17722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_645_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23690\,
            in1 => \N__22922\,
            in2 => \_gnd_net_\,
            in3 => \N__22899\,
            lcout => OPEN,
            ltout => \c0.n17734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15141_4_lut_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__23554\,
            in1 => \N__23538\,
            in2 => \N__23523\,
            in3 => \N__23515\,
            lcout => OPEN,
            ltout => \c0.n18000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_672_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23496\,
            in1 => \N__23490\,
            in2 => \N__23484\,
            in3 => \N__26268\,
            lcout => \c0.n29_adj_2408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23480\,
            in1 => \N__26704\,
            in2 => \_gnd_net_\,
            in3 => \N__23633\,
            lcout => data_in_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_4_lut_adj_407_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__23460\,
            in1 => \N__25710\,
            in2 => \N__23361\,
            in3 => \N__23222\,
            lcout => n120,
            ltout => \n120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25763\,
            in1 => \_gnd_net_\,
            in2 => \N__23184\,
            in3 => \N__23179\,
            lcout => data_in_frame_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1012_2_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23159\,
            in2 => \_gnd_net_\,
            in3 => \N__23131\,
            lcout => \c0.n2124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26196\,
            in1 => \N__23589\,
            in2 => \_gnd_net_\,
            in3 => \N__26703\,
            lcout => data_in_frame_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_699_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011111"
        )
    port map (
            in0 => \N__23108\,
            in1 => \N__23091\,
            in2 => \N__23678\,
            in3 => \N__23085\,
            lcout => \c0.n22_adj_2419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27604\,
            in1 => \N__23590\,
            in2 => \_gnd_net_\,
            in3 => \N__25909\,
            lcout => data_in_frame_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23634\,
            in1 => \N__24154\,
            in2 => \_gnd_net_\,
            in3 => \N__23691\,
            lcout => data_in_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27429\,
            in1 => \N__27938\,
            in2 => \N__28135\,
            in3 => \N__26967\,
            lcout => \c0.rx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24153\,
            in1 => \N__23674\,
            in2 => \_gnd_net_\,
            in3 => \N__26425\,
            lcout => data_in_frame_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_423_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27981\,
            lcout => \c0.rx.n17702\,
            ltout => \c0.rx.n17702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011100"
        )
    port map (
            in0 => \N__26733\,
            in1 => \N__26629\,
            in2 => \N__23652\,
            in3 => \N__28106\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_adj_400_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__27796\,
            in2 => \N__23649\,
            in3 => \N__26661\,
            lcout => OPEN,
            ltout => \c0.rx.n17704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27187\,
            in2 => \N__23640\,
            in3 => \N__26367\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25779\,
            in1 => \N__25493\,
            in2 => \_gnd_net_\,
            in3 => \N__23626\,
            lcout => data_in_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__23592\,
            in2 => \_gnd_net_\,
            in3 => \N__25780\,
            lcout => data_in_frame_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15143_4_lut_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23937\,
            in1 => \N__27060\,
            in2 => \N__26574\,
            in3 => \N__23998\,
            lcout => OPEN,
            ltout => \c0.n18002_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_582_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23967\,
            in1 => \N__26545\,
            in2 => \N__23718\,
            in3 => \N__34048\,
            lcout => \c0.n10498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4__2265_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23938\,
            in1 => \_gnd_net_\,
            in2 => \N__34221\,
            in3 => \N__26501\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4__2281_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23968\,
            in1 => \N__34198\,
            in2 => \_gnd_net_\,
            in3 => \N__24080\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__27920\,
            in2 => \N__28154\,
            in3 => \N__26958\,
            lcout => \c0.rx.n10988\,
            ltout => \c0.rx.n10988_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i9849_3_lut_4_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__27854\,
            in1 => \N__27528\,
            in2 => \N__23706\,
            in3 => \N__26863\,
            lcout => OPEN,
            ltout => \c0.rx.n12624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__28148\,
            in1 => \N__24041\,
            in2 => \N__23703\,
            in3 => \N__27855\,
            lcout => \c0.rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5__2288_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23999\,
            in1 => \N__34197\,
            in2 => \_gnd_net_\,
            in3 => \N__24102\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2__2291_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26902\,
            in1 => \N__34212\,
            in2 => \_gnd_net_\,
            in3 => \N__23700\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_570_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__23699\,
            in1 => \N__23948\,
            in2 => \N__26886\,
            in3 => \N__24060\,
            lcout => OPEN,
            ltout => \c0.n20_adj_2371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_580_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__26749\,
            in1 => \N__34280\,
            in2 => \N__24018\,
            in3 => \N__26910\,
            lcout => \c0.n10516\,
            ltout => \c0.n10516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_581_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__26523\,
            in1 => \N__29278\,
            in2 => \N__24009\,
            in3 => \N__26901\,
            lcout => \c0.n10367\,
            ltout => \c0.n10367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_622_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24000\,
            in1 => \N__23939\,
            in2 => \N__23985\,
            in3 => \N__27061\,
            lcout => \c0.n15_adj_2389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4__2289_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23972\,
            in1 => \_gnd_net_\,
            in2 => \N__34228\,
            in3 => \N__23949\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4__2273_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24079\,
            in1 => \N__23940\,
            in2 => \_gnd_net_\,
            in3 => \N__34216\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_619_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__34049\,
            in1 => \N__26571\,
            in2 => \_gnd_net_\,
            in3 => \N__26769\,
            lcout => \c0.n14_adj_2388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3__2282_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34050\,
            in1 => \N__34127\,
            in2 => \_gnd_net_\,
            in3 => \N__27689\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5__2280_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24101\,
            in1 => \N__34186\,
            in2 => \_gnd_net_\,
            in3 => \N__24197\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15770_1_lut_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34126\,
            lcout => \c0.n18631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15148_3_lut_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24213\,
            in1 => \N__24195\,
            in2 => \_gnd_net_\,
            in3 => \N__27658\,
            lcout => \c0.n18008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_569_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__24097\,
            in1 => \N__34297\,
            in2 => \N__24081\,
            in3 => \N__27688\,
            lcout => \c0.n18_adj_2370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_604_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24214\,
            in1 => \N__24196\,
            in2 => \N__26808\,
            in3 => \N__27659\,
            lcout => \c0.n13_adj_2380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3__2266_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34250\,
            in1 => \N__25783\,
            in2 => \_gnd_net_\,
            in3 => \N__34128\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6__2263_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27587\,
            in1 => \N__34187\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011110000"
        )
    port map (
            in0 => \N__26871\,
            in1 => \N__28082\,
            in2 => \N__27540\,
            in3 => \N__24045\,
            lcout => \c0.rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7__2270_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27714\,
            in1 => \N__34185\,
            in2 => \_gnd_net_\,
            in3 => \N__24215\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15146_4_lut_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27254\,
            in1 => \N__27728\,
            in2 => \N__27156\,
            in3 => \N__27712\,
            lcout => OPEN,
            ltout => \c0.n18006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_589_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27031\,
            in1 => \N__27001\,
            in2 => \N__24030\,
            in3 => \N__27675\,
            lcout => \c0.n14_adj_2375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7__2278_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__24216\,
            in1 => \_gnd_net_\,
            in2 => \N__27008\,
            in3 => \N__34183\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5__2272_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34181\,
            in1 => \N__27155\,
            in2 => \_gnd_net_\,
            in3 => \N__24198\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7__2262_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24179\,
            in1 => \N__34182\,
            in2 => \_gnd_net_\,
            in3 => \N__27713\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__0__2293_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27729\,
            in1 => \N__34184\,
            in2 => \_gnd_net_\,
            in3 => \N__26757\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28199\,
            in2 => \_gnd_net_\,
            in3 => \N__24117\,
            lcout => \c0.rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \c0.rx.n16532\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27354\,
            in2 => \_gnd_net_\,
            in3 => \N__24114\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.rx.n16532\,
            carryout => \c0.rx.n16533\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i2_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27336\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.rx.n16533\,
            carryout => \c0.rx.n16534\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27317\,
            in2 => \_gnd_net_\,
            in3 => \N__24108\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.rx.n16534\,
            carryout => \c0.rx.n16535\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i4_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27294\,
            in2 => \_gnd_net_\,
            in3 => \N__24105\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.rx.n16535\,
            carryout => \c0.rx.n16536\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i5_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28253\,
            in2 => \_gnd_net_\,
            in3 => \N__24279\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.rx.n16536\,
            carryout => \c0.rx.n16537\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i6_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29177\,
            in2 => \_gnd_net_\,
            in3 => \N__24276\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.rx.n16537\,
            carryout => \c0.rx.n16538\,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.r_Clock_Count__i7_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29204\,
            in2 => \_gnd_net_\,
            in3 => \N__24273\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49702\,
            ce => \N__24729\,
            sr => \N__24270\
        );

    \c0.rx.i1_2_lut_adj_399_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27447\,
            in2 => \_gnd_net_\,
            in3 => \N__24222\,
            lcout => \c0.rx.n12819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15562_2_lut_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39036\,
            in2 => \_gnd_net_\,
            in3 => \N__47412\,
            lcout => OPEN,
            ltout => \c0.n18225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1__2207_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111010001"
        )
    port map (
            in0 => \N__47689\,
            in1 => \N__47122\,
            in2 => \N__24261\,
            in3 => \N__42498\,
            lcout => \c0.data_out_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49695\,
            ce => \N__43423\,
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_4_lut_adj_408_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29200\,
            in1 => \N__29173\,
            in2 => \N__28196\,
            in3 => \N__28224\,
            lcout => OPEN,
            ltout => \c0.rx.n15905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i21_4_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000111010"
        )
    port map (
            in0 => \N__24258\,
            in1 => \N__24243\,
            in2 => \N__24228\,
            in3 => \N__28250\,
            lcout => OPEN,
            ltout => \c0.rx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13229_4_lut_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__28119\,
            in1 => \N__28161\,
            in2 => \N__24225\,
            in3 => \N__29154\,
            lcout => \c0.rx.n12\,
            ltout => \c0.rx.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15076_4_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__28286\,
            in1 => \N__27876\,
            in2 => \N__24732\,
            in3 => \N__27448\,
            lcout => \c0.rx.n11082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24645\,
            in2 => \_gnd_net_\,
            in3 => \N__24717\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \N__24660\
        );

    \c0.FRAME_MATCHER_i_i13_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24620\,
            in2 => \_gnd_net_\,
            in3 => \N__24393\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49684\,
            ce => 'H',
            sr => \N__24345\
        );

    \blink_counter_2483__i0_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24330\,
            in2 => \_gnd_net_\,
            in3 => \N__24324\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => n16609,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i1_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24321\,
            in2 => \_gnd_net_\,
            in3 => \N__24315\,
            lcout => n25,
            ltout => OPEN,
            carryin => n16609,
            carryout => n16610,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i2_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24312\,
            in2 => \_gnd_net_\,
            in3 => \N__24306\,
            lcout => n24,
            ltout => OPEN,
            carryin => n16610,
            carryout => n16611,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i3_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24303\,
            in2 => \_gnd_net_\,
            in3 => \N__24297\,
            lcout => n23,
            ltout => OPEN,
            carryin => n16611,
            carryout => n16612,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i4_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24294\,
            in2 => \_gnd_net_\,
            in3 => \N__24288\,
            lcout => n22_adj_2481,
            ltout => OPEN,
            carryin => n16612,
            carryout => n16613,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i5_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24285\,
            in2 => \_gnd_net_\,
            in3 => \N__24807\,
            lcout => n21,
            ltout => OPEN,
            carryin => n16613,
            carryout => n16614,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i6_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24804\,
            in2 => \_gnd_net_\,
            in3 => \N__24798\,
            lcout => n20,
            ltout => OPEN,
            carryin => n16614,
            carryout => n16615,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i7_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24795\,
            in2 => \_gnd_net_\,
            in3 => \N__24789\,
            lcout => n19,
            ltout => OPEN,
            carryin => n16615,
            carryout => n16616,
            clk => \N__49703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i8_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24786\,
            in2 => \_gnd_net_\,
            in3 => \N__24780\,
            lcout => n18_adj_2480,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => n16617,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i9_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24777\,
            in2 => \_gnd_net_\,
            in3 => \N__24771\,
            lcout => n17,
            ltout => OPEN,
            carryin => n16617,
            carryout => n16618,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i10_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24768\,
            in2 => \_gnd_net_\,
            in3 => \N__24762\,
            lcout => n16,
            ltout => OPEN,
            carryin => n16618,
            carryout => n16619,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i11_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24759\,
            in2 => \_gnd_net_\,
            in3 => \N__24753\,
            lcout => n15_adj_2479,
            ltout => OPEN,
            carryin => n16619,
            carryout => n16620,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i12_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24750\,
            in2 => \_gnd_net_\,
            in3 => \N__24744\,
            lcout => n14_adj_2478,
            ltout => OPEN,
            carryin => n16620,
            carryout => n16621,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i13_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24741\,
            in2 => \_gnd_net_\,
            in3 => \N__24735\,
            lcout => n13,
            ltout => OPEN,
            carryin => n16621,
            carryout => n16622,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i14_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24891\,
            in2 => \_gnd_net_\,
            in3 => \N__24885\,
            lcout => n12,
            ltout => OPEN,
            carryin => n16622,
            carryout => n16623,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i15_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24882\,
            in2 => \_gnd_net_\,
            in3 => \N__24876\,
            lcout => n11,
            ltout => OPEN,
            carryin => n16623,
            carryout => n16624,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i16_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24873\,
            in2 => \_gnd_net_\,
            in3 => \N__24867\,
            lcout => n10_adj_2467,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => n16625,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i17_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24864\,
            in2 => \_gnd_net_\,
            in3 => \N__24858\,
            lcout => n9,
            ltout => OPEN,
            carryin => n16625,
            carryout => n16626,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i18_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24855\,
            in2 => \_gnd_net_\,
            in3 => \N__24849\,
            lcout => n8,
            ltout => OPEN,
            carryin => n16626,
            carryout => n16627,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i19_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24846\,
            in2 => \_gnd_net_\,
            in3 => \N__24840\,
            lcout => n7_adj_2476,
            ltout => OPEN,
            carryin => n16627,
            carryout => n16628,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i20_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24837\,
            in2 => \_gnd_net_\,
            in3 => \N__24831\,
            lcout => n6,
            ltout => OPEN,
            carryin => n16628,
            carryout => n16629,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i21_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24823\,
            in2 => \_gnd_net_\,
            in3 => \N__24810\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n16629,
            carryout => n16630,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i22_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24982\,
            in2 => \_gnd_net_\,
            in3 => \N__24969\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n16630,
            carryout => n16631,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i23_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24961\,
            in2 => \_gnd_net_\,
            in3 => \N__24948\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n16631,
            carryout => n16632,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i24_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24943\,
            in2 => \_gnd_net_\,
            in3 => \N__24930\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => n16633,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2483__i25_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24923\,
            in2 => \_gnd_net_\,
            in3 => \N__24927\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15760_3_lut_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__28461\,
            in1 => \N__32907\,
            in2 => \_gnd_net_\,
            in3 => \N__32862\,
            lcout => \control.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.PHASES_i1_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35441\,
            lcout => \PIN_1_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49802\,
            ce => \N__35723\,
            sr => \N__28446\
        );

    \c0.byte_transmit_counter2_i6_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25239\,
            in1 => \N__25267\,
            in2 => \N__30659\,
            in3 => \N__30552\,
            lcout => \c0.byte_transmit_counter2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49851\,
            ce => 'H',
            sr => \N__25131\
        );

    \c0.i1_2_lut_4_lut_adj_771_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__25123\,
            in1 => \N__25069\,
            in2 => \N__25305\,
            in3 => \N__33087\,
            lcout => \c0.n4_adj_2203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11047_3_lut_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__48998\,
            in1 => \N__47960\,
            in2 => \_gnd_net_\,
            in3 => \N__48923\,
            lcout => OPEN,
            ltout => \c0.n13808_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_439_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25218\,
            in1 => \N__25299\,
            in2 => \N__25149\,
            in3 => \N__25260\,
            lcout => \c0.n14064\,
            ltout => \c0.n14064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_2_lut_3_lut_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29928\,
            in2 => \N__25146\,
            in3 => \N__30191\,
            lcout => n612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i5_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25281\,
            in1 => \N__25300\,
            in2 => \N__30650\,
            in3 => \N__30551\,
            lcout => \c0.byte_transmit_counter2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__25143\
        );

    \c0.i1_2_lut_4_lut_adj_773_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__33088\,
            in1 => \N__25269\,
            in2 => \N__25074\,
            in3 => \N__25124\,
            lcout => \c0.n4_adj_2201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_774_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__25125\,
            in1 => \N__25073\,
            in2 => \N__25226\,
            in3 => \N__33089\,
            lcout => \c0.n4_adj_2199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11300_1_lut_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30149\,
            lcout => \c0.tx2_transmit_N_1996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_2_lut_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25196\,
            in1 => \N__46160\,
            in2 => \_gnd_net_\,
            in3 => \N__25014\,
            lcout => \c0.n18254\,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \c0.n16479\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_3_lut_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25182\,
            in1 => \N__48622\,
            in2 => \_gnd_net_\,
            in3 => \N__24996\,
            lcout => \c0.n18253\,
            ltout => OPEN,
            carryin => \c0.n16479\,
            carryout => \c0.n16480\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_4_lut_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25200\,
            in1 => \N__47977\,
            in2 => \_gnd_net_\,
            in3 => \N__24987\,
            lcout => \c0.n18314\,
            ltout => OPEN,
            carryin => \c0.n16480\,
            carryout => \c0.n16481\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_5_lut_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25184\,
            in1 => \N__48986\,
            in2 => \_gnd_net_\,
            in3 => \N__25311\,
            lcout => \c0.n18315\,
            ltout => OPEN,
            carryin => \c0.n16481\,
            carryout => \c0.n16482\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_6_lut_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25197\,
            in1 => \N__48925\,
            in2 => \_gnd_net_\,
            in3 => \N__25308\,
            lcout => \c0.n18362\,
            ltout => OPEN,
            carryin => \c0.n16482\,
            carryout => \c0.n16483\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_7_lut_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25183\,
            in1 => \N__25301\,
            in2 => \_gnd_net_\,
            in3 => \N__25272\,
            lcout => \c0.n18316\,
            ltout => OPEN,
            carryin => \c0.n16483\,
            carryout => \c0.n16484\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_8_lut_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__25199\,
            in1 => \N__25268\,
            in2 => \_gnd_net_\,
            in3 => \N__25230\,
            lcout => \c0.n18317\,
            ltout => OPEN,
            carryin => \c0.n16484\,
            carryout => \c0.n16485\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_9_lut_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__25227\,
            in1 => \N__25198\,
            in2 => \_gnd_net_\,
            in3 => \N__25167\,
            lcout => \c0.n18318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15239_4_lut_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__28892\,
            in1 => \N__28815\,
            in2 => \N__40462\,
            in3 => \N__28868\,
            lcout => OPEN,
            ltout => \c0.n18100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__28818\,
            in1 => \N__28989\,
            in2 => \N__25155\,
            in3 => \N__28920\,
            lcout => \c0.data_out_frame2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15242_4_lut_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__28893\,
            in1 => \N__28816\,
            in2 => \N__41613\,
            in3 => \N__28869\,
            lcout => OPEN,
            ltout => \c0.n18103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__28988\,
            in2 => \N__25152\,
            in3 => \N__28919\,
            lcout => \c0.data_out_frame2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_665_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__25442\,
            in1 => \N__26205\,
            in2 => \N__25415\,
            in3 => \N__25398\,
            lcout => \c0.n27_adj_2405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__25391\,
            in1 => \N__25700\,
            in2 => \N__26726\,
            in3 => \N__25557\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11390_2_lut_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30070\,
            in2 => \_gnd_net_\,
            in3 => \N__30132\,
            lcout => \c0.n14161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27622\,
            in1 => \N__25370\,
            in2 => \_gnd_net_\,
            in3 => \N__25862\,
            lcout => data_in_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_4_lut_adj_403_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__27435\,
            in1 => \N__27549\,
            in2 => \N__28155\,
            in3 => \N__27944\,
            lcout => n158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_633_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25356\,
            in1 => \N__26012\,
            in2 => \_gnd_net_\,
            in3 => \N__26069\,
            lcout => \c0.n16982\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__26111\,
            in1 => \N__25552\,
            in2 => \N__26494\,
            in3 => \N__25677\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_416_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__27943\,
            in1 => \N__28150\,
            in2 => \_gnd_net_\,
            in3 => \N__27434\,
            lcout => n135_adj_2463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26718\,
            in1 => \N__25331\,
            in2 => \_gnd_net_\,
            in3 => \N__25865\,
            lcout => data_in_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__25553\,
            in1 => \N__27623\,
            in2 => \N__25704\,
            in3 => \N__26093\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26475\,
            in1 => \N__26240\,
            in2 => \_gnd_net_\,
            in3 => \N__25866\,
            lcout => data_in_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_635_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25830\,
            in1 => \N__25476\,
            in2 => \_gnd_net_\,
            in3 => \N__26298\,
            lcout => \c0.n17725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__30372\,
            in1 => \N__30783\,
            in2 => \N__30416\,
            in3 => \N__29850\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__25812\,
            in1 => \N__28020\,
            in2 => \N__25781\,
            in3 => \N__25806\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__25702\,
            in1 => \N__25556\,
            in2 => \N__26646\,
            in3 => \N__26070\,
            lcout => \c0.data_in_frame_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__25555\,
            in1 => \N__25703\,
            in2 => \N__26505\,
            in3 => \N__25945\,
            lcout => \c0.data_in_frame_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__25701\,
            in1 => \N__25554\,
            in2 => \N__27135\,
            in3 => \N__26038\,
            lcout => \c0.data_in_frame_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_631_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25494\,
            in1 => \N__25475\,
            in2 => \_gnd_net_\,
            in3 => \N__26037\,
            lcout => OPEN,
            ltout => \c0.n16981_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_652_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__26322\,
            in1 => \N__26302\,
            in2 => \N__26271\,
            in3 => \N__25944\,
            lcout => \c0.n20_adj_2397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_516_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111111111001"
        )
    port map (
            in0 => \N__26067\,
            in1 => \N__26247\,
            in2 => \N__26393\,
            in3 => \N__26142\,
            lcout => \c0.n20_adj_2350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1016_2_lut_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26004\,
            lcout => \c0.n2128\,
            ltout => \c0.n2128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_643_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26241\,
            in1 => \N__26226\,
            in2 => \N__26208\,
            in3 => \N__26141\,
            lcout => \c0.n22_adj_2392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1008_2_lut_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__26192\,
            in1 => \_gnd_net_\,
            in2 => \N__26174\,
            in3 => \_gnd_net_\,
            lcout => \c0.n2120\,
            ltout => \c0.n2120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_690_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26131\,
            in1 => \N__26112\,
            in2 => \N__26097\,
            in3 => \N__26094\,
            lcout => \c0.n19_adj_2415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_624_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26066\,
            in2 => \_gnd_net_\,
            in3 => \N__26036\,
            lcout => OPEN,
            ltout => \c0.n17721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_626_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26003\,
            in1 => \N__25940\,
            in2 => \N__25917\,
            in3 => \N__25900\,
            lcout => \c0.n10_adj_2390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26500\,
            in1 => \N__26389\,
            in2 => \_gnd_net_\,
            in3 => \N__26424\,
            lcout => data_in_frame_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101000101010"
        )
    port map (
            in0 => \N__27926\,
            in1 => \N__26956\,
            in2 => \N__28136\,
            in3 => \N__26354\,
            lcout => OPEN,
            ltout => \c0.rx.n18729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.n18729_bdd_4_lut_4_lut_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011100101"
        )
    port map (
            in0 => \N__28149\,
            in1 => \N__28287\,
            in2 => \N__26373\,
            in3 => \N__28005\,
            lcout => OPEN,
            ltout => \c0.rx.n18732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26370\,
            in3 => \N__27428\,
            lcout => \c0.rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__27542\,
            in1 => \N__28107\,
            in2 => \N__27807\,
            in3 => \N__26660\,
            lcout => \c0.rx.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100011001000"
        )
    port map (
            in0 => \N__27797\,
            in1 => \N__26864\,
            in2 => \N__28137\,
            in3 => \N__26957\,
            lcout => \c0.rx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_409_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27541\,
            in2 => \_gnd_net_\,
            in3 => \N__26659\,
            lcout => n12582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_418_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26339\,
            in1 => \N__27543\,
            in2 => \_gnd_net_\,
            in3 => \N__27856\,
            lcout => OPEN,
            ltout => \n4_adj_2471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__26689\,
            in1 => \N__28006\,
            in2 => \N__26325\,
            in3 => \N__27753\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__0__2285_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27039\,
            in1 => \N__26750\,
            in2 => \_gnd_net_\,
            in3 => \N__34195\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27846\,
            in1 => \N__27809\,
            in2 => \N__27548\,
            in3 => \N__27748\,
            lcout => \c0.rx.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2__2267_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26705\,
            in1 => \N__34194\,
            in2 => \_gnd_net_\,
            in3 => \N__26572\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_420_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__28200\,
            in1 => \N__29143\,
            in2 => \N__28260\,
            in3 => \N__28223\,
            lcout => \c0.rx.r_SM_Main_2_N_2088_2\,
            ltout => \c0.rx.r_SM_Main_2_N_2088_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_411_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27845\,
            in2 => \N__26664\,
            in3 => \N__26851\,
            lcout => \c0.rx.n161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0__2269_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34193\,
            in1 => \N__26637\,
            in2 => \_gnd_net_\,
            in3 => \N__27062\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2__2275_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26807\,
            in1 => \N__26573\,
            in2 => \_gnd_net_\,
            in3 => \N__34196\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__6__2287_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__26549\,
            in2 => \_gnd_net_\,
            in3 => \N__27258\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6__2271_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27276\,
            in1 => \N__26527\,
            in2 => \_gnd_net_\,
            in3 => \N__34219\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_613_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__29279\,
            in1 => \N__26903\,
            in2 => \N__26529\,
            in3 => \N__26768\,
            lcout => \c0.n8_adj_2385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_573_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__27274\,
            lcout => \c0.n15_adj_2372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2__2283_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34218\,
            in1 => \N__26904\,
            in2 => \_gnd_net_\,
            in3 => \N__26802\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_422_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__26865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26954\,
            lcout => n12527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7__2286_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34217\,
            in1 => \N__27009\,
            in2 => \_gnd_net_\,
            in3 => \N__26885\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_417_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__26866\,
            in1 => \_gnd_net_\,
            in2 => \N__27857\,
            in3 => \N__26955\,
            lcout => n151,
            ltout => \n151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15541_3_lut_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__27529\,
            in1 => \_gnd_net_\,
            in2 => \N__26811\,
            in3 => \N__27808\,
            lcout => \c0.rx.n18194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_563_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__26778\,
            in2 => \N__27035\,
            in3 => \N__27696\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_565_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__27150\,
            in1 => \N__26982\,
            in2 => \N__26772\,
            in3 => \N__27252\,
            lcout => \c0.n10493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6__2279_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27253\,
            in1 => \N__27275\,
            in2 => \_gnd_net_\,
            in3 => \N__34211\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010101"
        )
    port map (
            in0 => \N__27455\,
            in1 => \N__27234\,
            in2 => \N__28118\,
            in3 => \N__28269\,
            lcout => \c0.rx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5__2264_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27219\,
            in1 => \N__34210\,
            in2 => \_gnd_net_\,
            in3 => \N__27151\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1__2268_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34208\,
            in1 => \N__27134\,
            in2 => \_gnd_net_\,
            in3 => \N__34301\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0__2277_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27030\,
            in1 => \N__34209\,
            in2 => \_gnd_net_\,
            in3 => \N__27066\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_3_lut_4_lut_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27352\,
            in1 => \N__27334\,
            in2 => \N__27318\,
            in3 => \N__27292\,
            lcout => \c0.rx.n15902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10932_2_lut_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27000\,
            in2 => \_gnd_net_\,
            in3 => \N__27673\,
            lcout => \c0.n13693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_3_lut_4_lut_4_lut_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__27948\,
            in1 => \N__27450\,
            in2 => \N__28138\,
            in3 => \N__26974\,
            lcout => OPEN,
            ltout => \c0.rx.n11041_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__27451\,
            in1 => \N__34188\,
            in2 => \N__26922\,
            in3 => \N__28117\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15577_3_lut_4_lut_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__27858\,
            in1 => \N__27810\,
            in2 => \N__27547\,
            in3 => \N__27752\,
            lcout => \c0.rx.n18196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_559_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27711\,
            lcout => \c0.n6_adj_2368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3__2290_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27674\,
            in1 => \N__34180\,
            in2 => \_gnd_net_\,
            in3 => \N__27690\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1__2292_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34179\,
            in1 => \N__29283\,
            in2 => \_gnd_net_\,
            in3 => \N__27660\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i9777_4_lut_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011100000"
        )
    port map (
            in0 => \N__27645\,
            in1 => \N__28023\,
            in2 => \N__27586\,
            in3 => \N__27639\,
            lcout => OPEN,
            ltout => \c0.rx.n12552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27572\,
            in2 => \N__27630\,
            in3 => \N__28123\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_4_lut_adj_404_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27510\,
            in1 => \N__27456\,
            in2 => \N__28139\,
            in3 => \N__27947\,
            lcout => n164_adj_2464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15131_2_lut_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27353\,
            in2 => \_gnd_net_\,
            in3 => \N__27335\,
            lcout => OPEN,
            ltout => \c0.rx.n17990_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15163_4_lut_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28197\,
            in1 => \N__27316\,
            in2 => \N__27297\,
            in3 => \N__27293\,
            lcout => OPEN,
            ltout => \c0.rx.n18024_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__28252\,
            in1 => \_gnd_net_\,
            in2 => \N__28290\,
            in3 => \N__29150\,
            lcout => \c0.rx.n12828\,
            ltout => \c0.rx.n12828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15639_3_lut_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28022\,
            in2 => \N__28272\,
            in3 => \N__27946\,
            lcout => \c0.rx.n18303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15551_2_lut_3_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28251\,
            in1 => \N__28222\,
            in2 => \_gnd_net_\,
            in3 => \N__28198\,
            lcout => \c0.rx.n18211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_adj_419_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__28086\,
            in1 => \N__28021\,
            in2 => \_gnd_net_\,
            in3 => \N__27945\,
            lcout => \c0.rx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28334\,
            in1 => \N__28349\,
            in2 => \N__28386\,
            in3 => \N__28400\,
            lcout => \c0.tx.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__28494\,
            in1 => \N__28304\,
            in2 => \_gnd_net_\,
            in3 => \N__28319\,
            lcout => \c0.tx.n54\,
            ltout => \c0.tx.n54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i11043_2_lut_4_lut_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__28366\,
            in1 => \N__28417\,
            in2 => \N__27870\,
            in3 => \N__27866\,
            lcout => \c0.tx.r_SM_Main_2_N_2031_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5_3_lut_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__27867\,
            in1 => \_gnd_net_\,
            in2 => \N__28422\,
            in3 => \N__28367\,
            lcout => OPEN,
            ltout => \c0.tx.n47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__29400\,
            in1 => \N__28431\,
            in2 => \N__28425\,
            in3 => \N__29472\,
            lcout => \c0.tx.n11297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28421\,
            in2 => \_gnd_net_\,
            in3 => \N__28404\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \c0.tx.n16524\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28401\,
            in2 => \_gnd_net_\,
            in3 => \N__28389\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx.n16524\,
            carryout => \c0.tx.n16525\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28385\,
            in2 => \_gnd_net_\,
            in3 => \N__28371\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx.n16525\,
            carryout => \c0.tx.n16526\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i3_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28368\,
            in2 => \_gnd_net_\,
            in3 => \N__28353\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx.n16526\,
            carryout => \c0.tx.n16527\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28350\,
            in2 => \_gnd_net_\,
            in3 => \N__28338\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx.n16527\,
            carryout => \c0.tx.n16528\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28335\,
            in2 => \_gnd_net_\,
            in3 => \N__28323\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx.n16528\,
            carryout => \c0.tx.n16529\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i6_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28320\,
            in2 => \_gnd_net_\,
            in3 => \N__28308\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx.n16529\,
            carryout => \c0.tx.n16530\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i7_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28305\,
            in2 => \_gnd_net_\,
            in3 => \N__28293\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx.n16530\,
            carryout => \c0.tx.n16531\,
            clk => \N__49696\,
            ce => \N__29484\,
            sr => \N__28475\
        );

    \c0.tx.r_Clock_Count__i8_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28493\,
            in2 => \_gnd_net_\,
            in3 => \N__28497\,
            lcout => \c0.tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => \N__29483\,
            sr => \N__28479\
        );

    \control.i15748_2_lut_3_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__28460\,
            in1 => \N__32906\,
            in2 => \_gnd_net_\,
            in3 => \N__32858\,
            lcout => \control.n6_adj_2460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i19_3_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__35663\,
            in1 => \N__35444\,
            in2 => \_gnd_net_\,
            in3 => \N__35512\,
            lcout => \control.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i5146_2_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35664\,
            lcout => \control.PHASES_5_N_2152_1\,
            ltout => \control.PHASES_5_N_2152_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i1_2_lut_4_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110010"
        )
    port map (
            in0 => \N__35559\,
            in1 => \N__35442\,
            in2 => \N__28449\,
            in3 => \N__35337\,
            lcout => \control.n10356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__48032\,
            in1 => \N__48171\,
            in2 => \N__45336\,
            in3 => \N__28437\,
            lcout => \c0.n22_adj_2239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15978_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__28575\,
            in1 => \N__49045\,
            in2 => \N__40602\,
            in3 => \N__48031\,
            lcout => \c0.n18843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15914_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__31761\,
            in1 => \N__48604\,
            in2 => \N__46212\,
            in3 => \N__37872\,
            lcout => OPEN,
            ltout => \c0.n18801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18801_bdd_4_lut_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48605\,
            in1 => \N__31809\,
            in2 => \N__28440\,
            in3 => \N__40991\,
            lcout => \c0.n18804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18843_bdd_4_lut_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__49046\,
            in1 => \N__31644\,
            in2 => \N__29799\,
            in3 => \N__28563\,
            lcout => OPEN,
            ltout => \c0.n18846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__48926\,
            in1 => \N__49047\,
            in2 => \N__28557\,
            in3 => \N__28554\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49866\,
            ce => \N__48796\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15814_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__33999\,
            in1 => \N__48482\,
            in2 => \N__36087\,
            in3 => \N__46017\,
            lcout => OPEN,
            ltout => \c0.n18675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18675_bdd_4_lut_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48483\,
            in1 => \N__32991\,
            in2 => \N__28530\,
            in3 => \N__45454\,
            lcout => OPEN,
            ltout => \c0.n18678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__48029\,
            in1 => \N__35877\,
            in2 => \N__28527\,
            in3 => \N__48168\,
            lcout => \c0.n22_adj_2242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15879_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__28581\,
            in1 => \N__49048\,
            in2 => \N__29784\,
            in3 => \N__48030\,
            lcout => OPEN,
            ltout => \c0.n18741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18741_bdd_4_lut_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49049\,
            in1 => \N__29742\,
            in2 => \N__28524\,
            in3 => \N__31743\,
            lcout => OPEN,
            ltout => \c0.n18744_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__28521\,
            in1 => \N__49050\,
            in2 => \N__28515\,
            in3 => \N__48924\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49859\,
            ce => \N__48786\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i4_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__28987\,
            in1 => \N__28656\,
            in2 => \N__45092\,
            in3 => \N__28719\,
            lcout => \c0.data_out_frame2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15710_4_lut_4_lut_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001110000000"
        )
    port map (
            in0 => \N__29841\,
            in1 => \N__30340\,
            in2 => \N__30441\,
            in3 => \N__29926\,
            lcout => OPEN,
            ltout => \n17689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010111010"
        )
    port map (
            in0 => \N__30184\,
            in1 => \N__30762\,
            in2 => \N__28584\,
            in3 => \N__30435\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18681_bdd_4_lut_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48481\,
            in1 => \N__44806\,
            in2 => \N__44171\,
            in3 => \N__37929\,
            lcout => \c0.n18684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29925\,
            in1 => \N__30434\,
            in2 => \N__30355\,
            in3 => \N__30761\,
            lcout => \c0.tx2.n9639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18855_bdd_4_lut_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__48480\,
            in1 => \N__29733\,
            in2 => \N__41678\,
            in3 => \N__41154\,
            lcout => \c0.n18072\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i34_2_lut_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30430\,
            lcout => OPEN,
            ltout => \c0.tx2.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_4_lut_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__29876\,
            in1 => \N__30781\,
            in2 => \N__28566\,
            in3 => \N__30810\,
            lcout => \c0.tx2.n11312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_630_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30067\,
            in2 => \_gnd_net_\,
            in3 => \N__28696\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15633_3_lut_4_lut_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__28698\,
            in1 => \N__30071\,
            in2 => \N__37741\,
            in3 => \N__28861\,
            lcout => OPEN,
            ltout => \c0.n18284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i5_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__37721\,
            in1 => \N__28984\,
            in2 => \N__28746\,
            in3 => \N__28655\,
            lcout => \c0.data_out_frame2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_680_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__30068\,
            in1 => \N__28743\,
            in2 => \N__28593\,
            in3 => \N__28734\,
            lcout => \c0.n12704\,
            ltout => \c0.n12704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15621_3_lut_4_lut_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__30069\,
            in2 => \N__28722\,
            in3 => \N__28697\,
            lcout => \c0.n18287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15636_3_lut_4_lut_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__28699\,
            in1 => \N__30072\,
            in2 => \N__50664\,
            in3 => \N__28862\,
            lcout => OPEN,
            ltout => \c0.n18289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i3_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__50655\,
            in1 => \N__28983\,
            in2 => \N__28659\,
            in3 => \N__28654\,
            lcout => \c0.data_out_frame2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6035_bdd_4_lut_4_lut_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011111000"
        )
    port map (
            in0 => \N__28982\,
            in1 => \N__28924\,
            in2 => \N__28804\,
            in3 => \N__33083\,
            lcout => \c0.n18831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15218_4_lut_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__28859\,
            in1 => \N__37843\,
            in2 => \N__28803\,
            in3 => \N__28824\,
            lcout => OPEN,
            ltout => \c0.n18079_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i8_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__28793\,
            in2 => \N__28641\,
            in3 => \N__28986\,
            lcout => \c0.data_out_frame2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_661_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28638\,
            in1 => \N__28629\,
            in2 => \N__28617\,
            in3 => \N__28605\,
            lcout => \c0.n28_adj_2403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15224_4_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__28883\,
            in1 => \N__28791\,
            in2 => \N__44367\,
            in3 => \N__28860\,
            lcout => OPEN,
            ltout => \c0.n18085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i6_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__28792\,
            in1 => \N__28985\,
            in2 => \N__28938\,
            in3 => \N__28933\,
            lcout => \c0.data_out_frame2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15221_4_lut_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__28882\,
            in1 => \N__28787\,
            in2 => \N__41811\,
            in3 => \N__28858\,
            lcout => \c0.n18082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15527_3_lut_4_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__30161\,
            in1 => \N__37842\,
            in2 => \N__30599\,
            in3 => \N__30049\,
            lcout => \c0.n18270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_707_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__33176\,
            in1 => \N__33283\,
            in2 => \N__30066\,
            in3 => \N__30124\,
            lcout => \c0.n6035\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30213\,
            in2 => \_gnd_net_\,
            in3 => \N__28758\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \c0.tx2.n16539\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30227\,
            in2 => \_gnd_net_\,
            in3 => \N__28755\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx2.n16539\,
            carryout => \c0.tx2.n16540\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30240\,
            in2 => \_gnd_net_\,
            in3 => \N__28752\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx2.n16540\,
            carryout => \c0.tx2.n16541\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30830\,
            in2 => \_gnd_net_\,
            in3 => \N__28749\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx2.n16541\,
            carryout => \c0.tx2.n16542\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30252\,
            in2 => \_gnd_net_\,
            in3 => \N__29100\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx2.n16542\,
            carryout => \c0.tx2.n16543\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30854\,
            in2 => \_gnd_net_\,
            in3 => \N__29097\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx2.n16543\,
            carryout => \c0.tx2.n16544\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29087\,
            in2 => \_gnd_net_\,
            in3 => \N__29073\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx2.n16544\,
            carryout => \c0.tx2.n16545\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29063\,
            in2 => \_gnd_net_\,
            in3 => \N__29049\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx2.n16545\,
            carryout => \c0.tx2.n16546\,
            clk => \N__49827\,
            ce => \N__30726\,
            sr => \N__29021\
        );

    \c0.tx2.r_Clock_Count__i8_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29036\,
            in2 => \_gnd_net_\,
            in3 => \N__29046\,
            lcout => \c0.tx2.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49815\,
            ce => \N__30725\,
            sr => \N__29022\
        );

    \c0.add_2506_2_lut_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29127\,
            in2 => \N__42799\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_transmit_N_1947_0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \c0.n16517\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_3_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34774\,
            in2 => \_gnd_net_\,
            in3 => \N__28998\,
            lcout => \c0.tx_transmit_N_1947_1\,
            ltout => OPEN,
            carryin => \c0.n16517\,
            carryout => \c0.n16518\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_4_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35144\,
            in2 => \_gnd_net_\,
            in3 => \N__28995\,
            lcout => \c0.tx_transmit_N_1947_2\,
            ltout => OPEN,
            carryin => \c0.n16518\,
            carryout => \c0.n16519\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_5_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35049\,
            in2 => \_gnd_net_\,
            in3 => \N__28992\,
            lcout => \tx_transmit_N_1947_3\,
            ltout => OPEN,
            carryin => \c0.n16519\,
            carryout => \c0.n16520\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_6_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32484\,
            in2 => \_gnd_net_\,
            in3 => \N__29250\,
            lcout => \tx_transmit_N_1947_4\,
            ltout => OPEN,
            carryin => \c0.n16520\,
            carryout => \c0.n16521\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_7_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30927\,
            in2 => \_gnd_net_\,
            in3 => \N__29247\,
            lcout => \c0.tx_transmit_N_1947_5\,
            ltout => OPEN,
            carryin => \c0.n16521\,
            carryout => \c0.n16522\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_8_lut_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30887\,
            in2 => \_gnd_net_\,
            in3 => \N__29244\,
            lcout => \tx_transmit_N_1947_6\,
            ltout => OPEN,
            carryin => \c0.n16522\,
            carryout => \c0.n16523\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_9_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31035\,
            in2 => \_gnd_net_\,
            in3 => \N__29241\,
            lcout => \tx_transmit_N_1947_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__30554\,
            in1 => \N__29238\,
            in2 => \N__30642\,
            in3 => \N__45952\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49791\,
            ce => 'H',
            sr => \N__29223\
        );

    \c0.i1_2_lut_adj_759_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36051\,
            in2 => \_gnd_net_\,
            in3 => \N__31911\,
            lcout => \c0.n10782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29208\,
            in2 => \_gnd_net_\,
            in3 => \N__29181\,
            lcout => \c0.rx.n73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29289\,
            in2 => \_gnd_net_\,
            in3 => \N__32120\,
            lcout => \c0.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29354\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_4_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__32180\,
            in1 => \N__31347\,
            in2 => \N__31294\,
            in3 => \N__31398\,
            lcout => n9667,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__3__2253_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__43411\,
            in1 => \N__36584\,
            in2 => \_gnd_net_\,
            in3 => \N__46960\,
            lcout => data_out_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_2167_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32130\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1__2284_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__29274\,
            in2 => \_gnd_net_\,
            in3 => \N__34281\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__7__2241_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__46959\,
            in1 => \N__43412\,
            in2 => \_gnd_net_\,
            in3 => \N__29322\,
            lcout => data_out_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_585_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__47228\,
            in1 => \N__47685\,
            in2 => \_gnd_net_\,
            in3 => \N__46958\,
            lcout => n10973,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001100"
        )
    port map (
            in0 => \N__29328\,
            in1 => \N__30906\,
            in2 => \N__31295\,
            in3 => \N__32129\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__33706\,
            in1 => \N__33748\,
            in2 => \_gnd_net_\,
            in3 => \N__33914\,
            lcout => \r_Bit_Index_0_adj_2519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15180_3_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32322\,
            in1 => \N__31632\,
            in2 => \_gnd_net_\,
            in3 => \N__31149\,
            lcout => \c0.tx.n18041\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18747_bdd_4_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__35220\,
            in1 => \N__29493\,
            in2 => \N__31578\,
            in3 => \N__34359\,
            lcout => n18750,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011001"
        )
    port map (
            in0 => \N__31348\,
            in1 => \N__31285\,
            in2 => \_gnd_net_\,
            in3 => \N__29301\,
            lcout => OPEN,
            ltout => \n3_adj_2525_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29353\,
            in2 => \N__29370\,
            in3 => \N__29479\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_3_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31349\,
            in1 => \N__31399\,
            in2 => \_gnd_net_\,
            in3 => \N__31215\,
            lcout => \c0.tx.n17697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15687_2_lut_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42707\,
            in2 => \_gnd_net_\,
            in3 => \N__29321\,
            lcout => \c0.n18354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_4_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__31350\,
            in1 => \N__31400\,
            in2 => \N__31296\,
            in3 => \N__31216\,
            lcout => OPEN,
            ltout => \c0.tx.n11030_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101001001010"
        )
    port map (
            in0 => \N__31150\,
            in1 => \N__31289\,
            in2 => \N__29310\,
            in3 => \N__31074\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n18711_bdd_4_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__31413\,
            in1 => \N__29307\,
            in2 => \N__31461\,
            in3 => \N__31434\,
            lcout => \c0.tx.o_Tx_Serial_N_2062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15306_3_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31154\,
            in1 => \N__29381\,
            in2 => \_gnd_net_\,
            in3 => \N__29408\,
            lcout => \c0.tx.n18167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_817_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__35230\,
            in1 => \N__29295\,
            in2 => \N__30897\,
            in3 => \N__35081\,
            lcout => OPEN,
            ltout => \n10_adj_2532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__32523\,
            in1 => \N__32570\,
            in2 => \N__29412\,
            in3 => \N__29409\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_528_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32352\,
            in2 => \_gnd_net_\,
            in3 => \N__37335\,
            lcout => \c0.n10749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__31214\,
            in1 => \N__31327\,
            in2 => \N__31293\,
            in3 => \N__31395\,
            lcout => \c0.tx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__31396\,
            in1 => \N__31275\,
            in2 => \N__31345\,
            in3 => \N__31213\,
            lcout => \c0.tx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15125_2_lut_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31252\,
            in2 => \_gnd_net_\,
            in3 => \N__31326\,
            lcout => \c0.tx.n17984\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__4__2188_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46847\,
            in1 => \N__38058\,
            in2 => \_gnd_net_\,
            in3 => \N__36708\,
            lcout => data_out_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__42812\,
            in1 => \N__31407\,
            in2 => \N__36663\,
            in3 => \N__34870\,
            lcout => OPEN,
            ltout => \n10_adj_2537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_815_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__35092\,
            in1 => \N__29433\,
            in2 => \N__29388\,
            in3 => \N__35246\,
            lcout => OPEN,
            ltout => \n10_adj_2535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__32585\,
            in1 => \N__29382\,
            in2 => \N__29385\,
            in3 => \N__32529\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15574_2_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29427\,
            in2 => \_gnd_net_\,
            in3 => \N__42808\,
            lcout => \c0.n18188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__7__2185_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46855\,
            in1 => \N__38748\,
            in2 => \_gnd_net_\,
            in3 => \N__32357\,
            lcout => data_out_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_603_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32681\,
            in1 => \N__42606\,
            in2 => \_gnd_net_\,
            in3 => \N__34565\,
            lcout => \c0.n17883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_1_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31380\,
            lcout => n5155,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18753_bdd_4_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__29538\,
            in1 => \N__31554\,
            in2 => \N__29445\,
            in3 => \N__35245\,
            lcout => n18756,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__6__2226_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__47668\,
            in1 => \N__29426\,
            in2 => \N__43409\,
            in3 => \N__47121\,
            lcout => \c0.data_out_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42800\,
            in1 => \N__39908\,
            in2 => \_gnd_net_\,
            in3 => \N__36776\,
            lcout => \c0.n5_adj_2241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42801\,
            in1 => \N__31610\,
            in2 => \_gnd_net_\,
            in3 => \N__31698\,
            lcout => \c0.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__7__2233_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__47115\,
            in1 => \_gnd_net_\,
            in2 => \N__29550\,
            in3 => \N__43372\,
            lcout => data_out_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__6__2242_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__31599\,
            in1 => \N__47400\,
            in2 => \N__43410\,
            in3 => \N__47117\,
            lcout => data_out_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__7__2225_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__47116\,
            in1 => \N__43376\,
            in2 => \N__29562\,
            in3 => \N__47401\,
            lcout => data_out_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42811\,
            in1 => \N__29558\,
            in2 => \_gnd_net_\,
            in3 => \N__29546\,
            lcout => \c0.n2_adj_2229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_1266_i1_3_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47677\,
            in1 => \N__47394\,
            in2 => \_gnd_net_\,
            in3 => \N__47111\,
            lcout => n2837,
            ltout => \n2837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__5__2251_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43319\,
            in2 => \N__29529\,
            in3 => \N__29526\,
            lcout => data_out_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49690\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15651_2_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29525\,
            in2 => \_gnd_net_\,
            in3 => \N__42860\,
            lcout => \c0.n18189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i2658_4_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__29642\,
            in1 => \N__29627\,
            in2 => \N__29661\,
            in3 => \N__29675\,
            lcout => OPEN,
            ltout => \control.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i2661_4_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__29597\,
            in1 => \N__29583\,
            in2 => \N__29514\,
            in3 => \N__29612\,
            lcout => \control.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i0_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29511\,
            in2 => \_gnd_net_\,
            in3 => \N__29505\,
            lcout => \control.n10\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \control.n16647\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29502\,
            in2 => \_gnd_net_\,
            in3 => \N__29496\,
            lcout => \control.n9_adj_2459\,
            ltout => OPEN,
            carryin => \control.n16647\,
            carryout => \control.n16648\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i2_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29676\,
            in2 => \_gnd_net_\,
            in3 => \N__29664\,
            lcout => \control.pwm_delay_2\,
            ltout => OPEN,
            carryin => \control.n16648\,
            carryout => \control.n16649\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29660\,
            in2 => \_gnd_net_\,
            in3 => \N__29646\,
            lcout => \control.pwm_delay_3\,
            ltout => OPEN,
            carryin => \control.n16649\,
            carryout => \control.n16650\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i4_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29643\,
            in2 => \_gnd_net_\,
            in3 => \N__29631\,
            lcout => \control.pwm_delay_4\,
            ltout => OPEN,
            carryin => \control.n16650\,
            carryout => \control.n16651\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i5_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29628\,
            in2 => \_gnd_net_\,
            in3 => \N__29616\,
            lcout => \control.pwm_delay_5\,
            ltout => OPEN,
            carryin => \control.n16651\,
            carryout => \control.n16652\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i6_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29613\,
            in2 => \_gnd_net_\,
            in3 => \N__29601\,
            lcout => \control.pwm_delay_6\,
            ltout => OPEN,
            carryin => \control.n16652\,
            carryout => \control.n16653\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i7_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29598\,
            in2 => \_gnd_net_\,
            in3 => \N__29586\,
            lcout => \control.pwm_delay_7\,
            ltout => OPEN,
            carryin => \control.n16653\,
            carryout => \control.n16654\,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i8_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29582\,
            in2 => \_gnd_net_\,
            in3 => \N__29568\,
            lcout => \control.pwm_delay_8\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \control.n16655\,
            clk => \N__49778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.pwm_delay_2485__i9_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32900\,
            in2 => \_gnd_net_\,
            in3 => \N__29565\,
            lcout => \control.pwm_delay_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18885_bdd_4_lut_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__49075\,
            in1 => \N__29754\,
            in2 => \N__31731\,
            in3 => \N__29694\,
            lcout => OPEN,
            ltout => \c0.n18888_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_10_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__29700\,
            in1 => \N__49076\,
            in2 => \N__29709\,
            in3 => \N__48927\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49867\,
            ce => \N__48812\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15904_LC_10_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__31827\,
            in1 => \N__48602\,
            in2 => \N__31659\,
            in3 => \N__46162\,
            lcout => OPEN,
            ltout => \c0.n18789_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18789_bdd_4_lut_LC_10_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48603\,
            in1 => \N__29724\,
            in2 => \N__29706\,
            in3 => \N__35904\,
            lcout => OPEN,
            ltout => \c0.n18792_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_10_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__48035\,
            in1 => \N__37899\,
            in2 => \N__29703\,
            in3 => \N__48170\,
            lcout => \c0.n22_adj_2270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_10_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__33531\,
            in1 => \N__49074\,
            in2 => \N__29685\,
            in3 => \N__48034\,
            lcout => \c0.n18885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_494_LC_10_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43661\,
            in1 => \N__40751\,
            in2 => \N__45801\,
            in3 => \N__40976\,
            lcout => \c0.n10816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_758_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41082\,
            in2 => \_gnd_net_\,
            in3 => \N__46415\,
            lcout => OPEN,
            ltout => \c0.n10861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_775_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45357\,
            in1 => \N__40437\,
            in2 => \N__29688\,
            in3 => \N__40803\,
            lcout => \c0.n20_adj_2442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18795_bdd_4_lut_LC_10_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48623\,
            in1 => \N__31767\,
            in2 => \N__41722\,
            in3 => \N__33333\,
            lcout => \c0.n18798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_780_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31857\,
            in2 => \_gnd_net_\,
            in3 => \N__45202\,
            lcout => \c0.n10893\,
            ltout => \c0.n10893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_781_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41674\,
            in1 => \N__36335\,
            in2 => \N__29727\,
            in3 => \N__44167\,
            lcout => \c0.n17886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_705_LC_10_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33383\,
            in2 => \_gnd_net_\,
            in3 => \N__31856\,
            lcout => \c0.n18_adj_2423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_483_LC_10_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45815\,
            in1 => \N__41036\,
            in2 => \_gnd_net_\,
            in3 => \N__43662\,
            lcout => \c0.n17911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__46090\,
            in1 => \N__40844\,
            in2 => \N__50743\,
            in3 => \_gnd_net_\,
            lcout => \c0.n5_adj_2433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__48161\,
            in1 => \N__31773\,
            in2 => \N__48033\,
            in3 => \N__31716\,
            lcout => \c0.n22_adj_2373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_788_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37139\,
            lcout => \c0.n17748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_508_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37138\,
            in1 => \N__41077\,
            in2 => \_gnd_net_\,
            in3 => \N__45206\,
            lcout => \c0.n10688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__30773\,
            in1 => \N__29889\,
            in2 => \N__30366\,
            in3 => \N__29842\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i138_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38660\,
            in1 => \N__29723\,
            in2 => \_gnd_net_\,
            in3 => \N__50451\,
            lcout => data_out_frame2_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46091\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__41190\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__48624\,
            in1 => \N__44660\,
            in2 => \N__29802\,
            in3 => \N__46092\,
            lcout => \c0.n6_adj_2223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30439\,
            in1 => \N__30774\,
            in2 => \N__29849\,
            in3 => \N__30368\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15828_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__46187\,
            in1 => \N__36049\,
            in2 => \N__48649\,
            in3 => \N__45248\,
            lcout => OPEN,
            ltout => \c0.n18687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18687_bdd_4_lut_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48556\,
            in1 => \N__44624\,
            in2 => \N__29787\,
            in3 => \N__36314\,
            lcout => \c0.n18690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_518_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44742\,
            in1 => \N__44899\,
            in2 => \N__44805\,
            in3 => \N__41405\,
            lcout => \c0.n17795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__48557\,
            in1 => \N__31854\,
            in2 => \N__29772\,
            in3 => \N__46188\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__46189\,
            in1 => \N__44820\,
            in2 => \N__37792\,
            in3 => \N__48558\,
            lcout => \c0.n6_adj_2354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15973_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__43656\,
            in1 => \N__44741\,
            in2 => \N__48648\,
            in3 => \N__46186\,
            lcout => \c0.n18855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i46_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37785\,
            in1 => \N__39354\,
            in2 => \_gnd_net_\,
            in3 => \N__50445\,
            lcout => data_out_frame2_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10936_2_lut_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29918\,
            in2 => \_gnd_net_\,
            in3 => \N__30192\,
            lcout => \c0.n12359\,
            ltout => \c0.n12359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_782_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30162\,
            in1 => \N__33175\,
            in2 => \N__30138\,
            in3 => \N__33290\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_2261_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33177\,
            in2 => \N__30135\,
            in3 => \N__30050\,
            lcout => \c0.r_SM_Main_2_N_2034_0_adj_2213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49836\,
            ce => 'H',
            sr => \N__30131\
        );

    \c0.i1_2_lut_adj_448_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30045\,
            in2 => \_gnd_net_\,
            in3 => \N__33174\,
            lcout => \c0.n10958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4167_4_lut_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__30450\,
            in1 => \N__29828\,
            in2 => \N__29927\,
            in3 => \N__30438\,
            lcout => n6707,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11346_2_lut_4_lut_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__29877\,
            in1 => \N__30855\,
            in2 => \N__30831\,
            in3 => \N__30201\,
            lcout => \r_SM_Main_2_N_2031_1\,
            ltout => \r_SM_Main_2_N_2031_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15154_3_lut_4_lut_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__30356\,
            in1 => \N__30436\,
            in2 => \N__29808\,
            in3 => \N__30769\,
            lcout => n18014,
            ltout => \n18014_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15159_3_lut_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__30437\,
            in1 => \_gnd_net_\,
            in2 => \N__29805\,
            in3 => \N__30449\,
            lcout => n11545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i4_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__30675\,
            in1 => \N__48891\,
            in2 => \N__30600\,
            in3 => \N__30553\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__30459\
        );

    \c0.tx2.i1_2_lut_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33885\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33938\,
            lcout => n4_adj_2472,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33937\,
            in1 => \N__33680\,
            in2 => \_gnd_net_\,
            in3 => \N__33884\,
            lcout => \c0.tx2.n13800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15201_3_lut_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42387\,
            in1 => \N__43074\,
            in2 => \_gnd_net_\,
            in3 => \N__33936\,
            lcout => \c0.tx2.n18062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110011001"
        )
    port map (
            in0 => \N__30440\,
            in1 => \N__30367\,
            in2 => \_gnd_net_\,
            in3 => \N__30258\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_1__bdd_4_lut_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__33883\,
            in1 => \N__30294\,
            in2 => \N__33681\,
            in3 => \N__30282\,
            lcout => OPEN,
            ltout => \c0.tx2.n18717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18717_bdd_4_lut_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__30267\,
            in1 => \N__30789\,
            in2 => \N__30261\,
            in3 => \N__33679\,
            lcout => \c0.tx2.o_Tx_Serial_N_2062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4_4_lut_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30251\,
            in1 => \N__30239\,
            in2 => \N__30228\,
            in3 => \N__30212\,
            lcout => \c0.tx2.n10\,
            ltout => \c0.tx2.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5_3_lut_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__30853\,
            in1 => \_gnd_net_\,
            in2 => \N__30834\,
            in3 => \N__30829\,
            lcout => \c0.tx2.n12775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15200_3_lut_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30798\,
            in1 => \N__49179\,
            in2 => \_gnd_net_\,
            in3 => \N__33939\,
            lcout => \c0.tx2.n18061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i13_1_lut_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30782\,
            lcout => n11096,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15706_3_lut_4_lut_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001111"
        )
    port map (
            in0 => \N__33834\,
            in1 => \N__33450\,
            in2 => \N__47672\,
            in3 => \N__33794\,
            lcout => OPEN,
            ltout => \c0.n18260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_2168_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000010011"
        )
    port map (
            in0 => \N__30690\,
            in1 => \N__30696\,
            in2 => \N__30699\,
            in3 => \N__33765\,
            lcout => \c0.r_SM_Main_2_N_2034_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__30684\
        );

    \c0.i1_2_lut_3_lut_adj_637_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__32132\,
            in1 => \_gnd_net_\,
            in2 => \N__32178\,
            in3 => \N__47291\,
            lcout => \c0.n130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10860_2_lut_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32164\,
            in2 => \_gnd_net_\,
            in3 => \N__32131\,
            lcout => n12227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__47292\,
            in1 => \_gnd_net_\,
            in2 => \N__47691\,
            in3 => \N__47059\,
            lcout => \c0.n3465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__47058\,
            in1 => \N__47681\,
            in2 => \_gnd_net_\,
            in3 => \N__47293\,
            lcout => \c0.n4806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33515\,
            in1 => \N__33490\,
            in2 => \_gnd_net_\,
            in3 => \N__33469\,
            lcout => \c0.n85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__30876\,
            in1 => \N__30888\,
            in2 => \N__31005\,
            in3 => \N__30950\,
            lcout => byte_transmit_counter_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_533_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31016\,
            in1 => \N__30875\,
            in2 => \N__30867\,
            in3 => \N__31046\,
            lcout => \c0.n14068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__30866\,
            in2 => \N__31004\,
            in3 => \N__30949\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__32019\,
            in1 => \N__33402\,
            in2 => \N__31920\,
            in3 => \N__32187\,
            lcout => \UART_TRANSMITTER_state_7_N_1223_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__30993\,
            in1 => \N__35071\,
            in2 => \N__33858\,
            in3 => \N__30948\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__30951\,
            in1 => \N__30989\,
            in2 => \N__34856\,
            in3 => \N__33491\,
            lcout => byte_transmit_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__35190\,
            in1 => \N__33470\,
            in2 => \N__31003\,
            in3 => \N__30952\,
            lcout => byte_transmit_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__33516\,
            in1 => \N__42798\,
            in2 => \N__31001\,
            in3 => \N__30953\,
            lcout => byte_transmit_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_437_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47260\,
            in2 => \_gnd_net_\,
            in3 => \N__32293\,
            lcout => OPEN,
            ltout => \c0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__30982\,
            in1 => \N__34376\,
            in2 => \N__31056\,
            in3 => \N__30912\,
            lcout => n5341,
            ltout => \n5341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__31000\,
            in1 => \N__31034\,
            in2 => \N__31053\,
            in3 => \N__31050\,
            lcout => byte_transmit_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__30926\,
            in1 => \N__31020\,
            in2 => \N__31002\,
            in3 => \N__30954\,
            lcout => \c0.byte_transmit_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15139_4_lut_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__32024\,
            in1 => \N__47259\,
            in2 => \N__47615\,
            in3 => \N__32193\,
            lcout => \c0.n17998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15079_2_lut_3_lut_3_lut_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__31346\,
            in2 => \_gnd_net_\,
            in3 => \N__31397\,
            lcout => \c0.tx.n17938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011011000110"
        )
    port map (
            in0 => \N__46962\,
            in1 => \N__47257\,
            in2 => \N__47614\,
            in3 => \N__32262\,
            lcout => \UART_TRANSMITTER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__32241\,
            in2 => \N__47669\,
            in3 => \N__32280\,
            lcout => \UART_TRANSMITTER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__37101\,
            in1 => \N__34844\,
            in2 => \N__31083\,
            in3 => \N__42708\,
            lcout => n10_adj_2536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2723_2_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31487\,
            lcout => OPEN,
            ltout => \n5440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110000000000"
        )
    port map (
            in0 => \N__31170\,
            in1 => \N__31459\,
            in2 => \N__31095\,
            in3 => \N__31092\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15156_2_lut_3_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__31291\,
            in1 => \N__31073\,
            in2 => \_gnd_net_\,
            in3 => \N__31168\,
            lcout => n18016,
            ltout => \n18016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__31169\,
            in1 => \N__31488\,
            in2 => \N__31086\,
            in3 => \N__31153\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_636_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47536\,
            in2 => \_gnd_net_\,
            in3 => \N__46961\,
            lcout => n9_adj_2477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42781\,
            in1 => \N__34492\,
            in2 => \_gnd_net_\,
            in3 => \N__37443\,
            lcout => \c0.n8_adj_2207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31427\,
            in1 => \N__32226\,
            in2 => \N__32600\,
            in3 => \N__32524\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31151\,
            in1 => \N__31486\,
            in2 => \_gnd_net_\,
            in3 => \N__31455\,
            lcout => \c0.tx.n13802\,
            ltout => \c0.tx.n13802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4255_4_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__31292\,
            in1 => \N__31217\,
            in2 => \N__31062\,
            in3 => \N__32181\,
            lcout => OPEN,
            ltout => \c0.tx.n6796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__31218\,
            in1 => \N__31401\,
            in2 => \N__31059\,
            in3 => \N__31344\,
            lcout => \c0.tx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__31485\,
            in1 => \N__31467\,
            in2 => \N__31460\,
            in3 => \N__31101\,
            lcout => \c0.tx.n18711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15179_3_lut_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31428\,
            in1 => \N__32457\,
            in2 => \_gnd_net_\,
            in3 => \N__31148\,
            lcout => \c0.tx.n18040\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31110\,
            in1 => \N__31521\,
            in2 => \N__32613\,
            in3 => \N__32530\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42804\,
            in1 => \N__34728\,
            in2 => \_gnd_net_\,
            in3 => \N__32353\,
            lcout => \c0.n8_adj_2205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__5__2187_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46846\,
            in1 => \N__38034\,
            in2 => \_gnd_net_\,
            in3 => \N__37390\,
            lcout => data_out_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42803\,
            in1 => \N__34336\,
            in2 => \_gnd_net_\,
            in3 => \N__36557\,
            lcout => \c0.n8_adj_2232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32674\,
            in1 => \N__37389\,
            in2 => \_gnd_net_\,
            in3 => \N__42802\,
            lcout => \c0.n8_adj_2209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15152_3_lut_4_lut_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__31379\,
            in1 => \N__31325\,
            in2 => \N__31290\,
            in3 => \N__31207\,
            lcout => n18012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15305_3_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31155\,
            in1 => \N__31109\,
            in2 => \_gnd_net_\,
            in3 => \N__32646\,
            lcout => \c0.tx.n18166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15948_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__32625\,
            in1 => \N__35192\,
            in2 => \N__31563\,
            in3 => \N__34833\,
            lcout => \c0.n18753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18873_bdd_4_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__35193\,
            in1 => \N__31548\,
            in2 => \N__31539\,
            in3 => \N__31512\,
            lcout => OPEN,
            ltout => \n18876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_819_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__31494\,
            in1 => \N__35080\,
            in2 => \N__31524\,
            in3 => \N__35194\,
            lcout => n10_adj_2531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39941\,
            in1 => \N__42821\,
            in2 => \_gnd_net_\,
            in3 => \N__36745\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__31683\,
            in1 => \N__35191\,
            in2 => \N__31515\,
            in3 => \N__34834\,
            lcout => \c0.n18873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i5_3_lut_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36854\,
            in1 => \N__42820\,
            in2 => \_gnd_net_\,
            in3 => \N__34563\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i43_4_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__42822\,
            in1 => \N__37336\,
            in2 => \N__31506\,
            in3 => \N__34832\,
            lcout => n24_adj_2523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__34835\,
            in1 => \N__42823\,
            in2 => \N__31503\,
            in3 => \N__34683\,
            lcout => n10_adj_2533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15533_3_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__37340\,
            in1 => \N__47646\,
            in2 => \_gnd_net_\,
            in3 => \N__39837\,
            lcout => \c0.n18230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_825_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__34923\,
            in1 => \N__35093\,
            in2 => \N__32370\,
            in3 => \N__35247\,
            lcout => OPEN,
            ltout => \n10_adj_2528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__32614\,
            in1 => \N__31628\,
            in2 => \N__31635\,
            in3 => \N__32531\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15731_2_lut_3_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__43368\,
            in1 => \N__47634\,
            in2 => \_gnd_net_\,
            in3 => \N__47072\,
            lcout => \c0.n11016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_549_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34347\,
            in2 => \_gnd_net_\,
            in3 => \N__37284\,
            lcout => \c0.n10558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__5__2227_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__47345\,
            in1 => \N__43346\,
            in2 => \N__31614\,
            in3 => \N__47073\,
            lcout => data_out_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6__2250_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__47680\,
            in1 => \N__47118\,
            in2 => \N__43393\,
            in3 => \N__31587\,
            lcout => \c0.data_out_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31598\,
            in1 => \N__31586\,
            in2 => \_gnd_net_\,
            in3 => \N__42810\,
            lcout => \c0.n1_adj_2272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15707_3_lut_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__47679\,
            in1 => \N__36891\,
            in2 => \_gnd_net_\,
            in3 => \N__37485\,
            lcout => \c0.n18184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15958_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__32718\,
            in1 => \N__35195\,
            in2 => \N__32655\,
            in3 => \N__34867\,
            lcout => \c0.n18849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15604_2_lut_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42809\,
            lcout => \c0.n18377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__5__2235_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__43269\,
            in1 => \N__47119\,
            in2 => \_gnd_net_\,
            in3 => \N__31697\,
            lcout => data_out_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15657_2_lut_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37484\,
            in2 => \_gnd_net_\,
            in3 => \N__42712\,
            lcout => \c0.n18335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3__2237_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__47678\,
            in1 => \N__31674\,
            in2 => \N__43318\,
            in3 => \N__47120\,
            lcout => \c0.data_out_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15068_2_lut_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35574\,
            in2 => \_gnd_net_\,
            in3 => \N__35665\,
            lcout => \control.n17926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15091_2_lut_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35575\,
            in2 => \_gnd_net_\,
            in3 => \N__32921\,
            lcout => \control.n17950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37859\,
            in1 => \N__37653\,
            in2 => \N__40406\,
            in3 => \N__33332\,
            lcout => OPEN,
            ltout => \c0.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i154_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__32964\,
            in1 => \_gnd_net_\,
            in2 => \N__31662\,
            in3 => \N__31650\,
            lcout => \c0.data_out_frame2_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__50444\,
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41724\,
            in1 => \N__40791\,
            in2 => \N__36012\,
            in3 => \N__45455\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15649_3_lut_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46205\,
            in2 => \N__48682\,
            in3 => \N__37858\,
            lcout => \c0.n18266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15206_3_lut_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001011000010"
        )
    port map (
            in0 => \N__37740\,
            in1 => \N__48591\,
            in2 => \N__46210\,
            in3 => \_gnd_net_\,
            lcout => \c0.n18067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15557_2_lut_3_lut_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46201\,
            in2 => \N__48681\,
            in3 => \N__50671\,
            lcout => \c0.n18221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15606_3_lut_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110010"
        )
    port map (
            in0 => \N__44374\,
            in1 => \N__48595\,
            in2 => \N__46211\,
            in3 => \_gnd_net_\,
            lcout => \c0.n18360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15608_3_lut_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46206\,
            in2 => \N__48683\,
            in3 => \N__40468\,
            lcout => \c0.n18256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40940\,
            in1 => \N__40983\,
            in2 => \N__44172\,
            in3 => \N__37559\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i161_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31704\,
            in1 => \N__31710\,
            in2 => \N__31719\,
            in3 => \N__37761\,
            lcout => \c0.data_out_frame2_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49868\,
            ce => \N__50426\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_721_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44973\,
            in1 => \N__46262\,
            in2 => \N__44589\,
            in3 => \N__45669\,
            lcout => \c0.n15_adj_2429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_527_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44286\,
            in1 => \N__43819\,
            in2 => \_gnd_net_\,
            in3 => \N__43865\,
            lcout => \c0.n17847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_798_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__43818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33324\,
            lcout => \c0.n10867\,
            ltout => \c0.n10867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_806_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33644\,
            in1 => \N__36153\,
            in2 => \N__31791\,
            in3 => \N__45696\,
            lcout => \c0.n17_adj_2449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i59_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50263\,
            in1 => \N__38568\,
            in2 => \_gnd_net_\,
            in3 => \N__50742\,
            lcout => data_out_frame2_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_789_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46638\,
            in1 => \N__43745\,
            in2 => \_gnd_net_\,
            in3 => \N__50703\,
            lcout => OPEN,
            ltout => \c0.n17739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_709_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31866\,
            in1 => \N__44659\,
            in2 => \N__31788\,
            in3 => \N__43892\,
            lcout => \c0.n28_adj_2425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i137_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38720\,
            in1 => \N__31784\,
            in2 => \_gnd_net_\,
            in3 => \N__50261\,
            lcout => data_out_frame2_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18837_bdd_4_lut_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48487\,
            in1 => \N__31833\,
            in2 => \N__31785\,
            in3 => \N__37188\,
            lcout => \c0.n18840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i136_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42098\,
            in1 => \N__40984\,
            in2 => \_gnd_net_\,
            in3 => \N__50260\,
            lcout => data_out_frame2_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15909_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__35985\,
            in1 => \N__40389\,
            in2 => \N__48606\,
            in3 => \N__46190\,
            lcout => \c0.n18795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i152_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42099\,
            in1 => \N__31757\,
            in2 => \_gnd_net_\,
            in3 => \N__50262\,
            lcout => data_out_frame2_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i88_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50137\,
            in1 => \_gnd_net_\,
            in2 => \N__39633\,
            in3 => \N__44749\,
            lcout => data_out_frame2_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i42_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39503\,
            in1 => \N__31855\,
            in2 => \_gnd_net_\,
            in3 => \N__50134\,
            lcout => data_out_frame2_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i54_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50135\,
            in1 => \N__38846\,
            in2 => \_gnd_net_\,
            in3 => \N__44888\,
            lcout => data_out_frame2_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i114_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39087\,
            in1 => \N__40396\,
            in2 => \_gnd_net_\,
            in3 => \N__50131\,
            lcout => data_out_frame2_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15953_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__46185\,
            in1 => \N__48524\,
            in2 => \N__37602\,
            in3 => \N__33344\,
            lcout => \c0.n18837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i83_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40891\,
            in1 => \N__36183\,
            in2 => \_gnd_net_\,
            in3 => \N__50136\,
            lcout => data_out_frame2_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i146_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50133\,
            in1 => \N__38336\,
            in2 => \_gnd_net_\,
            in3 => \N__31823\,
            lcout => data_out_frame2_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i144_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39232\,
            in1 => \N__31805\,
            in2 => \_gnd_net_\,
            in3 => \N__50132\,
            lcout => data_out_frame2_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i50_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50254\,
            in1 => \N__39085\,
            in2 => \_gnd_net_\,
            in3 => \N__44040\,
            lcout => data_out_frame2_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i84_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50256\,
            in1 => \N__38982\,
            in2 => \_gnd_net_\,
            in3 => \N__41406\,
            lcout => data_out_frame2_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i99_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38271\,
            in1 => \N__41076\,
            in2 => \_gnd_net_\,
            in3 => \N__50259\,
            lcout => data_out_frame2_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i96_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50258\,
            in1 => \N__39234\,
            in2 => \_gnd_net_\,
            in3 => \N__43660\,
            lcout => data_out_frame2_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i128_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39233\,
            in1 => \N__40928\,
            in2 => \_gnd_net_\,
            in3 => \N__50253\,
            lcout => data_out_frame2_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i53_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50255\,
            in1 => \N__38907\,
            in2 => \_gnd_net_\,
            in3 => \N__36220\,
            lcout => data_out_frame2_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i87_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39705\,
            in1 => \N__50789\,
            in2 => \_gnd_net_\,
            in3 => \N__50257\,
            lcout => data_out_frame2_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_682_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41624\,
            in1 => \N__44967\,
            in2 => \N__36363\,
            in3 => \N__37128\,
            lcout => \c0.n16_adj_2412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_479_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45789\,
            in1 => \N__43655\,
            in2 => \_gnd_net_\,
            in3 => \N__40739\,
            lcout => \c0.n17727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i110_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50313\,
            in1 => \N__39343\,
            in2 => \_gnd_net_\,
            in3 => \N__44792\,
            lcout => data_out_frame2_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i151_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50314\,
            in1 => \N__41284\,
            in2 => \_gnd_net_\,
            in3 => \N__42368\,
            lcout => data_out_frame2_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__36216\,
            in1 => \_gnd_net_\,
            in2 => \N__44972\,
            in3 => \N__46139\,
            lcout => \c0.n5_adj_2436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i82_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50316\,
            in1 => \_gnd_net_\,
            in2 => \N__40750\,
            in3 => \N__39086\,
            lcout => data_out_frame2_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i58_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38650\,
            in1 => \N__31903\,
            in2 => \_gnd_net_\,
            in3 => \N__50315\,
            lcout => data_out_frame2_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32097\,
            in2 => \N__33573\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \c0.n16634\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33420\,
            in2 => \_gnd_net_\,
            in3 => \N__31884\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n16634\,
            carryout => \c0.n16635\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31952\,
            in2 => \_gnd_net_\,
            in3 => \N__31881\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n16635\,
            carryout => \c0.n16636\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33617\,
            in2 => \_gnd_net_\,
            in3 => \N__31878\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n16636\,
            carryout => \c0.n16637\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32060\,
            in2 => \_gnd_net_\,
            in3 => \N__31875\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n16637\,
            carryout => \c0.n16638\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31934\,
            in2 => \_gnd_net_\,
            in3 => \N__31872\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n16638\,
            carryout => \c0.n16639\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33543\,
            in2 => \_gnd_net_\,
            in3 => \N__31869\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n16639\,
            carryout => \c0.n16640\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32045\,
            in2 => \_gnd_net_\,
            in3 => \N__31974\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \c0.n16640\,
            carryout => \c0.n16641\,
            clk => \N__49829\,
            ce => \N__36516\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i8_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33603\,
            in2 => \_gnd_net_\,
            in3 => \N__31971\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \c0.n16642\,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i9_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33432\,
            in2 => \_gnd_net_\,
            in3 => \N__31968\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \c0.n16642\,
            carryout => \c0.n16643\,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i10_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33585\,
            in2 => \_gnd_net_\,
            in3 => \N__31965\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \c0.n16643\,
            carryout => \c0.n16644\,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32088\,
            in2 => \_gnd_net_\,
            in3 => \N__31962\,
            lcout => \c0.delay_counter_11\,
            ltout => OPEN,
            carryin => \c0.n16644\,
            carryout => \c0.n16645\,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i12_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32076\,
            in2 => \_gnd_net_\,
            in3 => \N__31959\,
            lcout => \c0.delay_counter_12\,
            ltout => OPEN,
            carryin => \c0.n16645\,
            carryout => \c0.n16646\,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2484__i13_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33557\,
            in2 => \_gnd_net_\,
            in3 => \N__31956\,
            lcout => \c0.delay_counter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49816\,
            ce => \N__36512\,
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31953\,
            in1 => \N__33591\,
            in2 => \N__31938\,
            in3 => \N__32031\,
            lcout => n26_adj_2466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_438_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__33789\,
            in1 => \N__32023\,
            in2 => \_gnd_net_\,
            in3 => \N__33851\,
            lcout => \c0.n98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15158_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__33852\,
            in1 => \N__33446\,
            in2 => \N__47128\,
            in3 => \N__33790\,
            lcout => \c0.n18019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_441_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33788\,
            in1 => \N__33850\,
            in2 => \_gnd_net_\,
            in3 => \N__33806\,
            lcout => n129,
            ltout => \n129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_567_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32168\,
            in2 => \N__32139\,
            in3 => \N__32136\,
            lcout => \c0.n1707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__32075\,
            in2 => \N__32064\,
            in3 => \N__32046\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__33853\,
            in1 => \N__33445\,
            in2 => \N__32025\,
            in3 => \N__33787\,
            lcout => n574,
            ltout => \n574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_618_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011011100"
        )
    port map (
            in0 => \N__47258\,
            in1 => \N__47085\,
            in2 => \N__31998\,
            in3 => \N__31995\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3__2205_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38931\,
            in1 => \N__47237\,
            in2 => \N__31989\,
            in3 => \N__46974\,
            lcout => \c0.data_out_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49793\,
            ce => \N__43425\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2__2206_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46973\,
            in1 => \N__39006\,
            in2 => \N__32235\,
            in3 => \N__47255\,
            lcout => \c0.data_out_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49793\,
            ce => \N__43425\,
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_587_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__47254\,
            in1 => \N__46970\,
            in2 => \_gnd_net_\,
            in3 => \N__32295\,
            lcout => n6_adj_2470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15119_2_lut_3_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__46968\,
            in1 => \N__32270\,
            in2 => \_gnd_net_\,
            in3 => \N__32256\,
            lcout => OPEN,
            ltout => \n17978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15531_4_lut_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100011111"
        )
    port map (
            in0 => \N__47550\,
            in1 => \N__46971\,
            in2 => \N__32298\,
            in3 => \N__32294\,
            lcout => n18202,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15708_4_lut_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__32258\,
            in1 => \N__47236\,
            in2 => \N__32274\,
            in3 => \N__46972\,
            lcout => n18368,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__46969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32257\,
            lcout => n22_adj_2522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15560_3_lut_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__47549\,
            in1 => \N__42493\,
            in2 => \_gnd_net_\,
            in3 => \N__37341\,
            lcout => \c0.n18226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i42_4_lut_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__33957\,
            in1 => \N__35072\,
            in2 => \N__32769\,
            in3 => \N__35218\,
            lcout => n21_adj_2524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000010111010"
        )
    port map (
            in0 => \N__47554\,
            in1 => \N__32220\,
            in2 => \N__47798\,
            in3 => \N__32214\,
            lcout => \UART_TRANSMITTER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15963_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__34008\,
            in1 => \N__34852\,
            in2 => \N__42561\,
            in3 => \N__35216\,
            lcout => OPEN,
            ltout => \c0.n18861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18861_bdd_4_lut_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__35217\,
            in1 => \N__36570\,
            in2 => \N__32208\,
            in3 => \N__32205\,
            lcout => OPEN,
            ltout => \n18864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_823_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__32307\,
            in1 => \N__35073\,
            in2 => \N__32328\,
            in3 => \N__35219\,
            lcout => OPEN,
            ltout => \n10_adj_2529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__32601\,
            in1 => \N__32321\,
            in2 => \N__32325\,
            in3 => \N__32513\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_496_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34701\,
            in2 => \_gnd_net_\,
            in3 => \N__32424\,
            lcout => \c0.n17850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_727_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34679\,
            in1 => \N__34593\,
            in2 => \N__37368\,
            in3 => \N__42494\,
            lcout => \c0.n6_adj_2276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i10_4_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__34699\,
            in1 => \N__34851\,
            in2 => \N__36603\,
            in3 => \N__42780\,
            lcout => n10_adj_2499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_543_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39834\,
            in1 => \N__36858\,
            in2 => \N__34525\,
            in3 => \N__36777\,
            lcout => \c0.n10550\,
            ltout => \c0.n10550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_712_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34700\,
            in1 => \N__32682\,
            in2 => \N__32301\,
            in3 => \N__32438\,
            lcout => \c0.n14_adj_2320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_540_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34678\,
            lcout => \c0.n10524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32712\,
            in1 => \N__43437\,
            in2 => \_gnd_net_\,
            in3 => \N__42779\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_545_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__32439\,
            in2 => \N__36659\,
            in3 => \N__32423\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_537_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34408\,
            in2 => \_gnd_net_\,
            in3 => \N__43148\,
            lcout => \c0.n6_adj_2361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_531_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36462\,
            in2 => \_gnd_net_\,
            in3 => \N__36709\,
            lcout => \c0.n10746\,
            ltout => \c0.n10746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_538_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32397\,
            in1 => \N__32385\,
            in2 => \N__32391\,
            in3 => \N__34439\,
            lcout => n17758,
            ltout => \n17758_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__2__2182_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__46853\,
            in1 => \N__34343\,
            in2 => \N__32388\,
            in3 => \N__37097\,
            lcout => data_out_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49752\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_666_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37442\,
            in1 => \N__37388\,
            in2 => \_gnd_net_\,
            in3 => \N__42469\,
            lcout => \c0.n10734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__34409\,
            in1 => \N__34871\,
            in2 => \N__32379\,
            in3 => \N__42830\,
            lcout => n10_adj_2461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_487_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34533\,
            in1 => \N__39751\,
            in2 => \N__37047\,
            in3 => \N__32358\,
            lcout => \c0.n17742\,
            ltout => \c0.n17742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__4__2180_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34962\,
            in1 => \N__36485\,
            in2 => \N__32331\,
            in3 => \N__43152\,
            lcout => \c0.data_out_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49739\,
            ce => \N__46854\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__5__2179_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32697\,
            in1 => \N__34656\,
            in2 => \N__32691\,
            in3 => \N__42540\,
            lcout => \c0.data_out_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49739\,
            ce => \N__46854\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_621_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34337\,
            in1 => \N__39750\,
            in2 => \_gnd_net_\,
            in3 => \N__37282\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_551_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34968\,
            in1 => \N__42937\,
            in2 => \N__32658\,
            in3 => \N__36746\,
            lcout => \c0.n17768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37537\,
            in1 => \N__43147\,
            in2 => \_gnd_net_\,
            in3 => \N__42817\,
            lcout => \c0.n5_adj_2220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42818\,
            in1 => \N__50924\,
            in2 => \_gnd_net_\,
            in3 => \N__34532\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32525\,
            in1 => \N__32618\,
            in2 => \N__32645\,
            in3 => \N__35019\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_579_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39984\,
            in1 => \N__50925\,
            in2 => \_gnd_net_\,
            in3 => \N__39893\,
            lcout => \c0.n10537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15584_2_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43527\,
            in2 => \_gnd_net_\,
            in3 => \N__42816\,
            lcout => \c0.n18265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__32748\,
            in2 => \N__32619\,
            in3 => \N__32535\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10351_3_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34590\,
            in1 => \N__39985\,
            in2 => \_gnd_net_\,
            in3 => \N__34857\,
            lcout => OPEN,
            ltout => \c0.n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i29_4_lut_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__42819\,
            in1 => \N__34858\,
            in2 => \N__32772\,
            in3 => \N__37043\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18849_bdd_4_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__40236\,
            in1 => \N__32757\,
            in2 => \N__32742\,
            in3 => \N__35234\,
            lcout => OPEN,
            ltout => \n18852_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__35235\,
            in1 => \N__32724\,
            in2 => \N__32751\,
            in3 => \N__35088\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15580_2_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32945\,
            in2 => \_gnd_net_\,
            in3 => \N__42814\,
            lcout => \c0.n18264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i10_4_lut_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__42815\,
            in1 => \N__34632\,
            in2 => \N__32733\,
            in3 => \N__34878\,
            lcout => n10_adj_2527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__4__2244_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__47632\,
            in1 => \N__47081\,
            in2 => \N__43317\,
            in3 => \N__35003\,
            lcout => \c0.data_out_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15643_2_lut_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42485\,
            in2 => \_gnd_net_\,
            in3 => \N__42813\,
            lcout => \c0.n18322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__1__2255_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__43260\,
            in1 => \N__47080\,
            in2 => \_gnd_net_\,
            in3 => \N__32711\,
            lcout => data_out_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15737_4_lut_4_lut_4_lut_3_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__47625\,
            in1 => \N__47320\,
            in2 => \_gnd_net_\,
            in3 => \N__47070\,
            lcout => n11017,
            ltout => \n11017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__0__2256_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__47071\,
            in1 => \N__32946\,
            in2 => \N__32949\,
            in3 => \N__47346\,
            lcout => data_out_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49705\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__4__2228_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32934\,
            in1 => \N__40277\,
            in2 => \_gnd_net_\,
            in3 => \N__43270\,
            lcout => data_out_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15603_2_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32933\,
            in2 => \_gnd_net_\,
            in3 => \N__42861\,
            lcout => \c0.n18191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i1_2_lut_4_lut_adj_814_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111111111"
        )
    port map (
            in0 => \N__35679\,
            in1 => \N__32905\,
            in2 => \N__35471\,
            in3 => \N__32857\,
            lcout => \control.n17251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i1_3_lut_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__35567\,
            in1 => \N__32925\,
            in2 => \_gnd_net_\,
            in3 => \N__35315\,
            lcout => \control.n10490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15757_2_lut_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32904\,
            in2 => \_gnd_net_\,
            in3 => \N__32856\,
            lcout => \control.PHASES_5__N_2160\,
            ltout => \control.PHASES_5__N_2160_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15769_4_lut_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111110"
        )
    port map (
            in0 => \N__35463\,
            in1 => \N__32823\,
            in2 => \N__32817\,
            in3 => \N__32813\,
            lcout => \control.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i1_2_lut_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35566\,
            lcout => \control.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.i15762_4_lut_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110010"
        )
    port map (
            in0 => \N__35462\,
            in1 => \N__32814\,
            in2 => \N__32802\,
            in3 => \N__35324\,
            lcout => \control.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i57_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50425\,
            in1 => \_gnd_net_\,
            in2 => \N__38724\,
            in3 => \N__40536\,
            lcout => data_out_frame2_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i122_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38661\,
            in1 => \N__35980\,
            in2 => \_gnd_net_\,
            in3 => \N__50423\,
            lcout => data_out_frame2_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i130_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50424\,
            in1 => \N__38340\,
            in2 => \_gnd_net_\,
            in3 => \N__35898\,
            lcout => data_out_frame2_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15784_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__48488\,
            in1 => \N__50711\,
            in2 => \N__50621\,
            in3 => \N__46197\,
            lcout => OPEN,
            ltout => \c0.n18639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18639_bdd_4_lut_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__37221\,
            in1 => \N__41089\,
            in2 => \N__32970\,
            in3 => \N__48489\,
            lcout => \c0.n18642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_689_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35979\,
            in2 => \_gnd_net_\,
            in3 => \N__44853\,
            lcout => \c0.n10700\,
            ltout => \c0.n10700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_535_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42054\,
            in1 => \N__43950\,
            in2 => \N__32967\,
            in3 => \N__35897\,
            lcout => \c0.n17841\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33030\,
            in1 => \N__33645\,
            in2 => \N__32958\,
            in3 => \N__33024\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46261\,
            in2 => \_gnd_net_\,
            in3 => \N__37183\,
            lcout => \c0.n17804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_710_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36104\,
            in1 => \N__40355\,
            in2 => \N__37622\,
            in3 => \N__45146\,
            lcout => \c0.n29_adj_2427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_432_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36184\,
            in1 => \N__33320\,
            in2 => \_gnd_net_\,
            in3 => \N__48220\,
            lcout => \c0.n10849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_426_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44898\,
            in2 => \_gnd_net_\,
            in3 => \N__41415\,
            lcout => \c0.n17874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_757_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45627\,
            in1 => \N__44457\,
            in2 => \_gnd_net_\,
            in3 => \N__45695\,
            lcout => \c0.n17908\,
            ltout => \c0.n17908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_706_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33018\,
            in1 => \N__45486\,
            in2 => \N__33009\,
            in3 => \N__44490\,
            lcout => OPEN,
            ltout => \c0.n30_adj_2424_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_717_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36387\,
            in1 => \N__33006\,
            in2 => \N__33000\,
            in3 => \N__32997\,
            lcout => \c0.n10577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i62_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50141\,
            in1 => \N__38460\,
            in2 => \_gnd_net_\,
            in3 => \N__44852\,
            lcout => data_out_frame2_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i142_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38459\,
            in1 => \N__32984\,
            in2 => \_gnd_net_\,
            in3 => \N__50139\,
            lcout => data_out_frame2_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i74_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50142\,
            in1 => \N__39510\,
            in2 => \_gnd_net_\,
            in3 => \N__43949\,
            lcout => data_out_frame2_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i147_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38277\,
            in1 => \N__43052\,
            in2 => \_gnd_net_\,
            in3 => \N__50140\,
            lcout => data_out_frame2_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i98_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50143\,
            in1 => \N__38335\,
            in2 => \_gnd_net_\,
            in3 => \N__33328\,
            lcout => data_out_frame2_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_800_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36306\,
            in2 => \_gnd_net_\,
            in3 => \N__40664\,
            lcout => \c0.n10829\,
            ltout => \c0.n10829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_747_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36255\,
            in1 => \N__37637\,
            in2 => \N__33294\,
            in3 => \N__46562\,
            lcout => \c0.n17755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i115_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40899\,
            in1 => \N__50613\,
            in2 => \_gnd_net_\,
            in3 => \N__50138\,
            lcout => data_out_frame2_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i97_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50123\,
            in1 => \N__38400\,
            in2 => \_gnd_net_\,
            in3 => \N__45766\,
            lcout => data_out_frame2_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i131_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38275\,
            in1 => \N__46637\,
            in2 => \_gnd_net_\,
            in3 => \N__50120\,
            lcout => data_out_frame2_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i61_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50121\,
            in1 => \N__50529\,
            in2 => \_gnd_net_\,
            in3 => \N__44949\,
            lcout => data_out_frame2_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_430_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__33289\,
            in1 => \N__33192\,
            in2 => \N__33183\,
            in3 => \N__33090\,
            lcout => n11114,
            ltout => \n11114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i123_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38563\,
            in1 => \_gnd_net_\,
            in2 => \N__33033\,
            in3 => \N__50710\,
            lcout => data_out_frame2_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i106_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39502\,
            in1 => \N__41703\,
            in2 => \_gnd_net_\,
            in3 => \N__50118\,
            lcout => data_out_frame2_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i127_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50119\,
            in1 => \N__39287\,
            in2 => \_gnd_net_\,
            in3 => \N__41751\,
            lcout => data_out_frame2_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i70_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44231\,
            in1 => \N__36313\,
            in2 => \_gnd_net_\,
            in3 => \N__50122\,
            lcout => data_out_frame2_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i71_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50148\,
            in1 => \N__41289\,
            in2 => \_gnd_net_\,
            in3 => \N__37129\,
            lcout => data_out_frame2_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i145_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38392\,
            in1 => \N__33345\,
            in2 => \_gnd_net_\,
            in3 => \N__50144\,
            lcout => data_out_frame2_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i86_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50150\,
            in1 => \N__38847\,
            in2 => \_gnd_net_\,
            in3 => \N__36039\,
            lcout => data_out_frame2_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i56_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39625\,
            in1 => \N__33372\,
            in2 => \_gnd_net_\,
            in3 => \N__50147\,
            lcout => data_out_frame2_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i148_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50145\,
            in1 => \N__38186\,
            in2 => \_gnd_net_\,
            in3 => \N__41999\,
            lcout => data_out_frame2_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i89_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38719\,
            in1 => \N__46467\,
            in2 => \_gnd_net_\,
            in3 => \N__50151\,
            lcout => data_out_frame2_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i45_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50146\,
            in1 => \_gnd_net_\,
            in2 => \N__41508\,
            in3 => \N__46697\,
            lcout => data_out_frame2_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i72_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42091\,
            in1 => \N__41657\,
            in2 => \_gnd_net_\,
            in3 => \N__50149\,
            lcout => data_out_frame2_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_744_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45394\,
            in2 => \_gnd_net_\,
            in3 => \N__42165\,
            lcout => \c0.n10887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i134_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50299\,
            in1 => \N__44232\,
            in2 => \_gnd_net_\,
            in3 => \N__45444\,
            lcout => data_out_frame2_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i111_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40149\,
            in1 => \N__42166\,
            in2 => \_gnd_net_\,
            in3 => \N__50297\,
            lcout => data_out_frame2_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i69_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50301\,
            in1 => \N__38107\,
            in2 => \_gnd_net_\,
            in3 => \N__50869\,
            lcout => data_out_frame2_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i67_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38276\,
            in1 => \N__43759\,
            in2 => \_gnd_net_\,
            in3 => \N__50300\,
            lcout => data_out_frame2_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i126_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50298\,
            in1 => \_gnd_net_\,
            in2 => \N__45403\,
            in3 => \N__38450\,
            lcout => data_out_frame2_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15789_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__45650\,
            in1 => \N__46081\,
            in2 => \N__48490\,
            in3 => \N__36185\,
            lcout => \c0.n18645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i73_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50302\,
            in1 => \N__39555\,
            in2 => \_gnd_net_\,
            in3 => \N__46382\,
            lcout => data_out_frame2_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i156_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__41413\,
            in1 => \N__33382\,
            in2 => \N__36264\,
            in3 => \N__36285\,
            lcout => \c0.data_out_frame2_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49839\,
            ce => \N__50350\,
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_435_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33584\,
            in1 => \N__33569\,
            in2 => \N__33558\,
            in3 => \N__33542\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18807_bdd_4_lut_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__43954\,
            in1 => \N__33390\,
            in2 => \N__48689\,
            in3 => \N__44329\,
            lcout => \c0.n18810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15695_3_lut_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__48635\,
            in1 => \N__45088\,
            in2 => \_gnd_net_\,
            in3 => \N__46089\,
            lcout => \c0.n18371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15704_3_lut_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__46088\,
            in1 => \N__41620\,
            in2 => \_gnd_net_\,
            in3 => \N__48636\,
            lcout => \c0.n18374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i156_2_lut_3_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__33514\,
            in1 => \N__33492\,
            in2 => \_gnd_net_\,
            in3 => \N__33471\,
            lcout => \c0.n155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_436_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33431\,
            in1 => \N__33419\,
            in2 => \_gnd_net_\,
            in3 => \N__33408\,
            lcout => n25_adj_2468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i81_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39155\,
            in1 => \N__46520\,
            in2 => \_gnd_net_\,
            in3 => \N__50429\,
            lcout => data_out_frame2_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15919_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__46117\,
            in1 => \N__45575\,
            in2 => \N__48491\,
            in3 => \N__40746\,
            lcout => \c0.n18807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15207_4_lut_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__33951\,
            in1 => \N__48389\,
            in2 => \N__46708\,
            in3 => \N__46118\,
            lcout => \c0.n18068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4698_2_lut_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__46116\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48372\,
            lcout => \c0.n7263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i101_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38109\,
            in1 => \N__45185\,
            in2 => \_gnd_net_\,
            in3 => \N__50427\,
            lcout => data_out_frame2_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i65_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50428\,
            in1 => \N__38399\,
            in2 => \_gnd_net_\,
            in3 => \N__46345\,
            lcout => data_out_frame2_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011000000000"
        )
    port map (
            in0 => \N__33882\,
            in1 => \N__33940\,
            in2 => \N__33753\,
            in3 => \N__33707\,
            lcout => \r_Bit_Index_1_adj_2518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15579_3_lut_4_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__33857\,
            in1 => \N__33813\,
            in2 => \N__47670\,
            in3 => \N__33795\,
            lcout => \c0.n18259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110000000000"
        )
    port map (
            in0 => \N__33752\,
            in1 => \N__33667\,
            in2 => \N__33723\,
            in3 => \N__33708\,
            lcout => \r_Bit_Index_2_adj_2517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_811_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50871\,
            in1 => \N__41090\,
            in2 => \_gnd_net_\,
            in3 => \N__46341\,
            lcout => \c0.n17715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33618\,
            in2 => \_gnd_net_\,
            in3 => \N__33602\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i52_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38981\,
            in1 => \N__44087\,
            in2 => \_gnd_net_\,
            in3 => \N__50430\,
            lcout => data_out_frame2_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1__2276_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34229\,
            in1 => \N__34273\,
            in2 => \_gnd_net_\,
            in3 => \N__34308\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3__2274_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34257\,
            in1 => \N__34029\,
            in2 => \_gnd_net_\,
            in3 => \N__34230\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15693_2_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39755\,
            in2 => \_gnd_net_\,
            in3 => \N__42797\,
            lcout => \c0.n18365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i100_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38187\,
            in1 => \N__43797\,
            in2 => \_gnd_net_\,
            in3 => \N__50431\,
            lcout => data_out_frame2_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i150_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50433\,
            in1 => \N__44229\,
            in2 => \_gnd_net_\,
            in3 => \N__33989\,
            lcout => data_out_frame2_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i55_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39700\,
            in1 => \N__40657\,
            in2 => \_gnd_net_\,
            in3 => \N__50434\,
            lcout => data_out_frame2_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i113_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50432\,
            in1 => \_gnd_net_\,
            in2 => \N__39159\,
            in3 => \N__46287\,
            lcout => data_out_frame2_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i41_4_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__34869\,
            in1 => \N__33975\,
            in2 => \N__35248\,
            in3 => \N__33969\,
            lcout => n18_adj_2526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__3__2189_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36624\,
            in1 => \N__46851\,
            in2 => \_gnd_net_\,
            in3 => \N__38133\,
            lcout => data_out_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_586_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36539\,
            in2 => \_gnd_net_\,
            in3 => \N__36623\,
            lcout => \c0.n17761\,
            ltout => \c0.n17761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_536_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34630\,
            in1 => \N__40310\,
            in2 => \N__34383\,
            in3 => \N__36802\,
            lcout => \c0.n17844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__2__2190_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__34380\,
            in1 => \N__47313\,
            in2 => \N__38217\,
            in3 => \N__36540\,
            lcout => data_out_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_601_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34365\,
            in1 => \N__34485\,
            in2 => \N__39993\,
            in3 => \N__36803\,
            lcout => \c0.n17826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i44_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42150\,
            in1 => \N__43845\,
            in2 => \_gnd_net_\,
            in3 => \N__50435\,
            lcout => data_out_frame2_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15869_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42897\,
            in1 => \N__35236\,
            in2 => \N__36444\,
            in3 => \N__34868\,
            lcout => \c0.n18747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_555_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35857\,
            in2 => \_gnd_net_\,
            in3 => \N__37545\,
            lcout => OPEN,
            ltout => \c0.n17807_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__2__2174_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34458\,
            in1 => \N__34342\,
            in2 => \N__34350\,
            in3 => \N__42942\,
            lcout => \c0.data_out_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49781\,
            ce => \N__46856\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_715_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34341\,
            in1 => \N__36937\,
            in2 => \_gnd_net_\,
            in3 => \N__37283\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__6__2178_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__37017\,
            in2 => \N__34536\,
            in3 => \N__34519\,
            lcout => \c0.data_out_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49781\,
            ce => \N__46856\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_615_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39942\,
            in1 => \N__47733\,
            in2 => \N__34493\,
            in3 => \N__39907\,
            lcout => \c0.n6_adj_2367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__3__2181_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34452\,
            in1 => \N__36646\,
            in2 => \N__34446\,
            in3 => \N__37361\,
            lcout => \c0.data_out_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49781\,
            ce => \N__46856\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_590_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34723\,
            in2 => \_gnd_net_\,
            in3 => \N__34698\,
            lcout => \c0.n17835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_499_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37093\,
            in2 => \_gnd_net_\,
            in3 => \N__36968\,
            lcout => OPEN,
            ltout => \c0.data_out_9__2__N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_502_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40334\,
            in1 => \N__34710\,
            in2 => \N__34425\,
            in3 => \N__34607\,
            lcout => OPEN,
            ltout => \c0.n15_adj_2319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__7__2177_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34394\,
            in1 => \N__36489\,
            in2 => \N__34422\,
            in3 => \N__34419\,
            lcout => \c0.data_out_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49766\,
            ce => \N__46821\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__6__2170_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34912\,
            in1 => \N__34410\,
            in2 => \N__50923\,
            in3 => \N__34395\,
            lcout => data_out_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49766\,
            ce => \N__46821\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_610_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34631\,
            in1 => \N__34911\,
            in2 => \N__34955\,
            in3 => \N__37544\,
            lcout => \c0.n17718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_564_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50914\,
            in1 => \N__34724\,
            in2 => \N__43533\,
            in3 => \N__39864\,
            lcout => \c0.n17774\,
            ltout => \c0.n17774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__3__2173_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36938\,
            in2 => \N__34704\,
            in3 => \N__34569\,
            lcout => \c0.data_out_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49766\,
            ce => \N__46821\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__5__2171_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36831\,
            in1 => \N__34591\,
            in2 => \N__36558\,
            in3 => \N__34647\,
            lcout => \c0.data_out_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49753\,
            ce => \N__46843\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_490_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34677\,
            in2 => \_gnd_net_\,
            in3 => \N__36853\,
            lcout => \c0.n6_adj_2314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_568_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34913\,
            in2 => \_gnd_net_\,
            in3 => \N__37534\,
            lcout => OPEN,
            ltout => \c0.n10801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__0__2176_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34646\,
            in1 => \N__36747\,
            in2 => \N__34635\,
            in3 => \N__36897\,
            lcout => \c0.data_out_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49753\,
            ce => \N__46843\,
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_552_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34914\,
            in1 => \N__34608\,
            in2 => \N__34956\,
            in3 => \N__36830\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__1__2175_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35859\,
            in1 => \N__37535\,
            in2 => \N__34596\,
            in3 => \N__36909\,
            lcout => \c0.data_out_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49753\,
            ce => \N__46843\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_577_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42600\,
            in2 => \_gnd_net_\,
            in3 => \N__34564\,
            lcout => \c0.n17819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_485_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39836\,
            in2 => \_gnd_net_\,
            in3 => \N__37433\,
            lcout => \c0.n6_adj_2277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42870\,
            in1 => \N__34948\,
            in2 => \_gnd_net_\,
            in3 => \N__36716\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__34876\,
            in1 => \N__40309\,
            in2 => \N__34932\,
            in3 => \N__42871\,
            lcout => n10_adj_2505,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__6__2186_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37434\,
            in1 => \N__46852\,
            in2 => \_gnd_net_\,
            in3 => \N__38772\,
            lcout => data_out_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15528_2_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39835\,
            in2 => \_gnd_net_\,
            in3 => \N__42868\,
            lcout => OPEN,
            ltout => \c0.n18222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15864_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__34884\,
            in1 => \N__35249\,
            in2 => \N__34929\,
            in3 => \N__34877\,
            lcout => OPEN,
            ltout => \c0.n18693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18693_bdd_4_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__35250\,
            in1 => \N__35802\,
            in2 => \N__34926\,
            in3 => \N__34983\,
            lcout => n18696,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42869\,
            in1 => \N__37071\,
            in2 => \_gnd_net_\,
            in3 => \N__34910\,
            lcout => \c0.n5_adj_2347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15968_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__35231\,
            in1 => \N__34974\,
            in2 => \N__35013\,
            in3 => \N__34872\,
            lcout => OPEN,
            ltout => \c0.n18867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18867_bdd_4_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__35262\,
            in1 => \N__34989\,
            in2 => \N__35253\,
            in3 => \N__35232\,
            lcout => OPEN,
            ltout => \n18870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_821_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__35233\,
            in1 => \N__35106\,
            in2 => \N__35097\,
            in3 => \N__35094\,
            lcout => n10_adj_2530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__7__2193_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__39183\,
            in1 => \N__47871\,
            in2 => \N__47810\,
            in3 => \N__39900\,
            lcout => \c0.data_out_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35853\,
            in1 => \N__36807\,
            in2 => \_gnd_net_\,
            in3 => \N__42872\,
            lcout => \c0.n5_adj_2214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15601_2_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35004\,
            in2 => \_gnd_net_\,
            in3 => \N__42873\,
            lcout => \c0.n18190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__2__2246_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__47142\,
            in1 => \N__43264\,
            in2 => \N__35814\,
            in3 => \N__47690\,
            lcout => \c0.data_out_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15721_2_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__47127\,
            in1 => \N__43259\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n11277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42866\,
            in1 => \N__35822\,
            in2 => \_gnd_net_\,
            in3 => \N__35793\,
            lcout => \c0.n2_adj_2348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15666_2_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37249\,
            in2 => \_gnd_net_\,
            in3 => \N__42865\,
            lcout => \c0.n18334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4__2196_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__38487\,
            in1 => \N__47883\,
            in2 => \N__47814\,
            in3 => \N__35852\,
            lcout => \c0.data_out_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__2__2230_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35823\,
            in1 => \N__40270\,
            in2 => \_gnd_net_\,
            in3 => \N__43265\,
            lcout => data_out_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15665_2_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35810\,
            lcout => \c0.n18223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__2__2238_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__43347\,
            in1 => \N__35792\,
            in2 => \_gnd_net_\,
            in3 => \N__47123\,
            lcout => data_out_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \control.PHASES_i4_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35576\,
            lcout => \PIN_24_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49838\,
            ce => \N__35760\,
            sr => \N__35748\
        );

    \control.PHASES_i5_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35470\,
            in2 => \_gnd_net_\,
            in3 => \N__35545\,
            lcout => \PIN_23_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49847\,
            ce => \N__35727\,
            sr => \N__35700\
        );

    \control.i1_4_lut_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110001"
        )
    port map (
            in0 => \N__35691\,
            in1 => \N__35577\,
            in2 => \N__35472\,
            in3 => \N__35325\,
            lcout => \control.PHASES_5_N_2130_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_786_LC_13_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44437\,
            in1 => \N__50823\,
            in2 => \N__35277\,
            in3 => \N__41324\,
            lcout => \c0.n15_adj_2445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_802_LC_13_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35899\,
            in2 => \_gnd_net_\,
            in3 => \N__35984\,
            lcout => \c0.n10890\,
            ltout => \c0.n10890_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_805_LC_13_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50620\,
            in1 => \N__35961\,
            in2 => \N__35949\,
            in3 => \N__40560\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i155_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35931\,
            in1 => \N__35946\,
            in2 => \N__35934\,
            in3 => \N__41897\,
            lcout => \c0.data_out_frame2_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__50419\,
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_784_LC_13_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35930\,
            in1 => \N__40535\,
            in2 => \_gnd_net_\,
            in3 => \N__36243\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i157_LC_13_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36138\,
            in1 => \N__35913\,
            in2 => \N__35907\,
            in3 => \N__40703\,
            lcout => \c0.data_out_frame2_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__50419\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_693_LC_13_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__35900\,
            in1 => \_gnd_net_\,
            in2 => \N__43958\,
            in3 => \_gnd_net_\,
            lcout => \c0.n10825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i166_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36072\,
            in1 => \N__44913\,
            in2 => \N__35868\,
            in3 => \N__37743\,
            lcout => \c0.data_out_frame2_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49879\,
            ce => \N__50467\,
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_adj_532_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37802\,
            in1 => \N__44160\,
            in2 => \_gnd_net_\,
            in3 => \N__46475\,
            lcout => \c0.n16_adj_2358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_428_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36228\,
            in2 => \_gnd_net_\,
            in3 => \N__40777\,
            lcout => OPEN,
            ltout => \c0.n10720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_783_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36149\,
            in1 => \N__36070\,
            in2 => \N__36192\,
            in3 => \N__42978\,
            lcout => \c0.n17838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_797_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46535\,
            in2 => \_gnd_net_\,
            in3 => \N__36189\,
            lcout => \c0.n10819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36134\,
            in1 => \N__41564\,
            in2 => \_gnd_net_\,
            in3 => \N__50885\,
            lcout => OPEN,
            ltout => \c0.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i158_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36071\,
            in1 => \N__36117\,
            in2 => \N__36108\,
            in3 => \N__36105\,
            lcout => \c0.data_out_frame2_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49879\,
            ce => \N__50467\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_778_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41950\,
            in2 => \_gnd_net_\,
            in3 => \N__36429\,
            lcout => \c0.n10839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i68_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38182\,
            in1 => \N__40776\,
            in2 => \_gnd_net_\,
            in3 => \N__50244\,
            lcout => data_out_frame2_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i120_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50241\,
            in1 => \N__39632\,
            in2 => \_gnd_net_\,
            in3 => \N__40197\,
            lcout => data_out_frame2_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_792_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36060\,
            in1 => \N__36050\,
            in2 => \N__37583\,
            in3 => \N__36239\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_793_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36011\,
            in1 => \N__45506\,
            in2 => \N__35988\,
            in3 => \N__42052\,
            lcout => \c0.n17792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i112_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40096\,
            in1 => \N__42223\,
            in2 => \_gnd_net_\,
            in3 => \N__50240\,
            lcout => data_out_frame2_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i139_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50243\,
            in1 => \N__38564\,
            in2 => \_gnd_net_\,
            in3 => \N__43019\,
            lcout => data_out_frame2_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_803_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36227\,
            in1 => \N__40775\,
            in2 => \_gnd_net_\,
            in3 => \N__46534\,
            lcout => \c0.n17859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i135_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50242\,
            in1 => \N__41288\,
            in2 => \_gnd_net_\,
            in3 => \N__42261\,
            lcout => data_out_frame2_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i48_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50128\,
            in1 => \N__40098\,
            in2 => \_gnd_net_\,
            in3 => \N__44649\,
            lcout => data_out_frame2_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i107_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39425\,
            in1 => \N__37212\,
            in2 => \_gnd_net_\,
            in3 => \N__50124\,
            lcout => data_out_frame2_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i43_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50127\,
            in1 => \N__39426\,
            in2 => \_gnd_net_\,
            in3 => \N__41555\,
            lcout => data_out_frame2_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i78_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39350\,
            in1 => \N__44613\,
            in2 => \_gnd_net_\,
            in3 => \N__50130\,
            lcout => data_out_frame2_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i132_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50126\,
            in1 => \N__38174\,
            in2 => \_gnd_net_\,
            in3 => \N__41946\,
            lcout => data_out_frame2_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i64_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39231\,
            in1 => \N__41184\,
            in2 => \_gnd_net_\,
            in3 => \N__50129\,
            lcout => data_out_frame2_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i129_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50125\,
            in1 => \_gnd_net_\,
            in2 => \N__38388\,
            in3 => \N__37178\,
            lcout => data_out_frame2_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_506_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43752\,
            in1 => \N__50702\,
            in2 => \N__46645\,
            in3 => \N__41366\,
            lcout => \c0.n10864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i124_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41451\,
            in1 => \N__36426\,
            in2 => \_gnd_net_\,
            in3 => \N__50246\,
            lcout => data_out_frame2_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i66_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50249\,
            in1 => \_gnd_net_\,
            in2 => \N__38320\,
            in3 => \N__44309\,
            lcout => data_out_frame2_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i116_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38980\,
            in1 => \N__45040\,
            in2 => \_gnd_net_\,
            in3 => \N__50245\,
            lcout => data_out_frame2_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i92_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50251\,
            in1 => \N__41452\,
            in2 => \_gnd_net_\,
            in3 => \N__45614\,
            lcout => data_out_frame2_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i47_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40148\,
            in1 => \N__41853\,
            in2 => \_gnd_net_\,
            in3 => \N__50248\,
            lcout => data_out_frame2_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i90_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50250\,
            in1 => \N__38639\,
            in2 => \_gnd_net_\,
            in3 => \N__45574\,
            lcout => data_out_frame2_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i94_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38445\,
            in1 => \N__45234\,
            in2 => \_gnd_net_\,
            in3 => \N__50252\,
            lcout => data_out_frame2_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i133_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50247\,
            in1 => \N__38083\,
            in2 => \_gnd_net_\,
            in3 => \N__48219\,
            lcout => data_out_frame2_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i85_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50402\,
            in1 => \_gnd_net_\,
            in2 => \N__38905\,
            in3 => \N__41025\,
            lcout => data_out_frame2_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i143_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39282\,
            in1 => \N__42290\,
            in2 => \_gnd_net_\,
            in3 => \N__50401\,
            lcout => data_out_frame2_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_678_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45613\,
            in1 => \N__45654\,
            in2 => \N__46474\,
            in3 => \N__45570\,
            lcout => \c0.n10_adj_2411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i105_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39554\,
            in1 => \N__45849\,
            in2 => \_gnd_net_\,
            in3 => \N__50398\,
            lcout => data_out_frame2_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i117_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50399\,
            in1 => \_gnd_net_\,
            in2 => \N__38904\,
            in3 => \N__44418\,
            lcout => data_out_frame2_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i91_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__45655\,
            in1 => \_gnd_net_\,
            in2 => \N__38556\,
            in3 => \N__50403\,
            lcout => data_out_frame2_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i125_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50400\,
            in1 => \N__50505\,
            in2 => \_gnd_net_\,
            in3 => \N__45003\,
            lcout => data_out_frame2_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_762_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45039\,
            in1 => \N__45233\,
            in2 => \_gnd_net_\,
            in3 => \N__41325\,
            lcout => \c0.n10_adj_2440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_530_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44994\,
            in1 => \N__41357\,
            in2 => \_gnd_net_\,
            in3 => \N__45435\,
            lcout => \c0.n6_adj_2357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15983_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__41015\,
            in1 => \N__46120\,
            in2 => \N__48688\,
            in3 => \N__50586\,
            lcout => OPEN,
            ltout => \c0.n18879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18879_bdd_4_lut_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__41227\,
            in1 => \N__48631\,
            in2 => \N__36366\,
            in3 => \N__50868\,
            lcout => \c0.n18160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15799_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__36428\,
            in1 => \N__45041\,
            in2 => \N__48687\,
            in3 => \N__46119\,
            lcout => \c0.n18657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_694_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41865\,
            lcout => \c0.n10852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_794_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40689\,
            in1 => \N__44330\,
            in2 => \N__36348\,
            in3 => \N__36315\,
            lcout => \c0.n14_adj_2447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i108_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__42039\,
            in1 => \_gnd_net_\,
            in2 => \N__42148\,
            in3 => \N__50404\,
            lcout => data_out_frame2_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i63_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50405\,
            in1 => \_gnd_net_\,
            in2 => \N__39288\,
            in3 => \N__44683\,
            lcout => data_out_frame2_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15809_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__36398\,
            in1 => \N__48637\,
            in2 => \N__36279\,
            in3 => \N__46122\,
            lcout => \c0.n18669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46121\,
            in1 => \_gnd_net_\,
            in2 => \N__37679\,
            in3 => \N__40551\,
            lcout => \c0.n5_adj_2274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15690_3_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__41815\,
            in1 => \N__48638\,
            in2 => \_gnd_net_\,
            in3 => \N__46123\,
            lcout => \c0.n18308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_702_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37179\,
            in2 => \_gnd_net_\,
            in3 => \N__44677\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_704_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46397\,
            in1 => \N__36427\,
            in2 => \N__36402\,
            in3 => \N__42977\,
            lcout => \c0.n17780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i149_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38108\,
            in1 => \N__36399\,
            in2 => \_gnd_net_\,
            in3 => \N__50463\,
            lcout => data_out_frame2_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i41_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50464\,
            in1 => \_gnd_net_\,
            in2 => \N__39552\,
            in3 => \N__41365\,
            lcout => data_out_frame2_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i49_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37675\,
            in1 => \N__39136\,
            in2 => \_gnd_net_\,
            in3 => \N__50465\,
            lcout => data_out_frame2_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_808_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46331\,
            in2 => \_gnd_net_\,
            in3 => \N__50870\,
            lcout => OPEN,
            ltout => \c0.n10870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_713_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37671\,
            in1 => \N__37213\,
            in2 => \N__36390\,
            in3 => \N__44086\,
            lcout => \c0.n27_adj_2428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_741_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45856\,
            in1 => \N__44810\,
            in2 => \N__46719\,
            in3 => \N__40656\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__48690\,
            in1 => \N__46064\,
            in2 => \N__36375\,
            in3 => \N__41364\,
            lcout => \c0.n6_adj_2275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_594_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39986\,
            in1 => \N__36553\,
            in2 => \_gnd_net_\,
            in3 => \N__36630\,
            lcout => \c0.n10542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15726_2_lut_3_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__47686\,
            in1 => \N__47354\,
            in2 => \_gnd_net_\,
            in3 => \N__47137\,
            lcout => \c0.n11056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15522_2_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38507\,
            in2 => \_gnd_net_\,
            in3 => \N__47353\,
            lcout => OPEN,
            ltout => \c0.n18199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2__2198_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__47138\,
            in1 => \N__47687\,
            in2 => \N__36492\,
            in3 => \N__42941\,
            lcout => \c0.data_out_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49818\,
            ce => \N__47898\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_498_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40311\,
            in2 => \_gnd_net_\,
            in3 => \N__37066\,
            lcout => \c0.n17832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7__2201_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47065\,
            in1 => \N__47358\,
            in2 => \N__39576\,
            in3 => \N__36435\,
            lcout => \c0.data_out_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49807\,
            ce => \N__43424\,
            sr => \_gnd_net_\
        );

    \c0.i15536_3_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__37483\,
            in1 => \N__47603\,
            in2 => \_gnd_net_\,
            in3 => \N__37278\,
            lcout => OPEN,
            ltout => \c0.n18242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6__2202_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__47064\,
            in1 => \N__39654\,
            in2 => \N__36465\,
            in3 => \N__47357\,
            lcout => \c0.data_out_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49807\,
            ce => \N__43424\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47734\,
            in1 => \N__36458\,
            in2 => \_gnd_net_\,
            in3 => \N__42857\,
            lcout => \c0.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15570_3_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__47602\,
            in1 => \N__36890\,
            in2 => \_gnd_net_\,
            in3 => \N__43529\,
            lcout => \c0.n18247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15535_3_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__47610\,
            in1 => \N__39756\,
            in2 => \_gnd_net_\,
            in3 => \N__37277\,
            lcout => OPEN,
            ltout => \c0.n18238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5__2203_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__47063\,
            in1 => \N__38789\,
            in2 => \N__36810\,
            in3 => \N__47356\,
            lcout => \c0.data_out_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49807\,
            ce => \N__43424\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4__2204_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47355\,
            in1 => \N__38864\,
            in2 => \N__40023\,
            in3 => \N__47066\,
            lcout => \c0.data_out_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49807\,
            ce => \N__43424\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__1__2183_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36626\,
            in1 => \N__36786\,
            in2 => \N__36684\,
            in3 => \N__36769\,
            lcout => \c0.data_out_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49795\,
            ce => \N__46844\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_592_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36735\,
            in2 => \_gnd_net_\,
            in3 => \N__36717\,
            lcout => \c0.n17745\,
            ltout => \c0.n17745_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__7__2169_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36675\,
            in1 => \N__37005\,
            in2 => \N__36666\,
            in3 => \N__42605\,
            lcout => \c0.data_out_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49795\,
            ce => \N__46844\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36933\,
            in1 => \N__36625\,
            in2 => \_gnd_net_\,
            in3 => \N__42858\,
            lcout => \c0.n8_adj_2219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15544_2_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__42859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36591\,
            lcout => \c0.n18376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__5__2211_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39305\,
            in2 => \_gnd_net_\,
            in3 => \N__47380\,
            lcout => \c0.data_out_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => \N__43413\,
            sr => \N__43478\
        );

    \c0.i3_4_lut_adj_539_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37092\,
            in1 => \N__37070\,
            in2 => \N__37036\,
            in3 => \N__37469\,
            lcout => \c0.n17730\,
            ltout => \c0.n17730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_544_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37004\,
            in1 => \N__36989\,
            in2 => \N__36972\,
            in3 => \N__36969\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_546_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42536\,
            in2 => \N__36954\,
            in3 => \N__36951\,
            lcout => \c0.n17877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_443_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39741\,
            in1 => \N__43528\,
            in2 => \_gnd_net_\,
            in3 => \N__37275\,
            lcout => \c0.n17816\,
            ltout => \c0.n17816_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36942\,
            in1 => \N__40322\,
            in2 => \N__36912\,
            in3 => \N__36908\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37276\,
            in1 => \N__39742\,
            in2 => \N__37503\,
            in3 => \N__42929\,
            lcout => \c0.n17786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__1__2199_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__47365\,
            in1 => \N__47140\,
            in2 => \N__38595\,
            in3 => \N__36870\,
            lcout => \c0.data_out_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49767\,
            ce => \N__47885\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_572_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36829\,
            lcout => \c0.n17829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0__2208_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__39111\,
            in1 => \N__43382\,
            in2 => \N__47809\,
            in3 => \N__37536\,
            lcout => data_out_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39821\,
            in1 => \N__37313\,
            in2 => \_gnd_net_\,
            in3 => \N__42489\,
            lcout => \c0.n10680\,
            ltout => \c0.n10680_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15682_4_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__37494\,
            in1 => \N__47660\,
            in2 => \N__37488\,
            in3 => \N__37482\,
            lcout => \c0.n18250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_513_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37441\,
            in2 => \_gnd_net_\,
            in3 => \N__37403\,
            lcout => \c0.n17771\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1__2215_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__47139\,
            in1 => \N__47688\,
            in2 => \N__39453\,
            in3 => \N__47402\,
            lcout => data_out_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49742\,
            ce => \N__43396\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__4__2212_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39381\,
            in2 => \_gnd_net_\,
            in3 => \N__47398\,
            lcout => \c0.data_out_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49728\,
            ce => \N__43383\,
            sr => \N__43462\
        );

    \c0.i1_3_lut_4_lut_adj_505_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37220\,
            in1 => \N__46233\,
            in2 => \N__42275\,
            in3 => \N__37187\,
            lcout => \c0.n17880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15894_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__50819\,
            in1 => \N__46165\,
            in2 => \N__48703\,
            in3 => \N__41323\,
            lcout => OPEN,
            ltout => \c0.n18759_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18759_bdd_4_lut_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__37140\,
            in1 => \N__40589\,
            in2 => \N__37692\,
            in3 => \N__48678\,
            lcout => \c0.n18762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_14_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40590\,
            in1 => \N__41229\,
            in2 => \N__37689\,
            in3 => \N__41189\,
            lcout => \c0.n10778\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i121_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46234\,
            in1 => \N__38715\,
            in2 => \_gnd_net_\,
            in3 => \N__50473\,
            lcout => data_out_frame2_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49887\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15938_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__40941\,
            in1 => \N__40198\,
            in2 => \N__48704\,
            in3 => \N__46166\,
            lcout => \c0.n18813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_429_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40199\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40942\,
            lcout => \c0.n10920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_431_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46303\,
            in1 => \N__42265\,
            in2 => \N__45861\,
            in3 => \N__41766\,
            lcout => \c0.n17783\,
            ltout => \c0.n17783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37821\,
            in1 => \N__43675\,
            in2 => \N__37644\,
            in3 => \N__37641\,
            lcout => OPEN,
            ltout => \c0.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i153_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37626\,
            in1 => \N__44709\,
            in2 => \N__37605\,
            in3 => \N__40173\,
            lcout => \c0.data_out_frame2_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__50474\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_751_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41035\,
            lcout => OPEN,
            ltout => \c0.n10813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_687_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37587\,
            in1 => \N__46487\,
            in2 => \N__37563\,
            in3 => \N__37560\,
            lcout => OPEN,
            ltout => \c0.n15_adj_2414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i162_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37908\,
            in1 => \N__41109\,
            in2 => \N__37902\,
            in3 => \N__40550\,
            lcout => \c0.data_out_frame2_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__50474\,
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_739_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45540\,
            in1 => \N__41882\,
            in2 => \N__40629\,
            in3 => \N__37754\,
            lcout => OPEN,
            ltout => \c0.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i160_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40164\,
            in1 => \N__37887\,
            in2 => \N__37875\,
            in3 => \N__40671\,
            lcout => \c0.data_out_frame2_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49880\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_725_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40475\,
            lcout => \c0.n6_adj_2430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_433_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__41817\,
            in1 => \N__37860\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17777\,
            ltout => \c0.n17777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_726_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50672\,
            in1 => \N__37812\,
            in2 => \N__37806\,
            in3 => \N__44513\,
            lcout => \c0.n10617\,
            ltout => \c0.n10617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_731_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37803\,
            in2 => \N__37764\,
            in3 => \N__41577\,
            lcout => \c0.n17765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_723_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37742\,
            in2 => \_gnd_net_\,
            in3 => \N__44375\,
            lcout => \c0.n17853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i60_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41454\,
            in1 => \N__45107\,
            in2 => \_gnd_net_\,
            in3 => \N__50356\,
            lcout => data_out_frame2_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i95_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50360\,
            in1 => \N__39278\,
            in2 => \_gnd_net_\,
            in3 => \N__41322\,
            lcout => data_out_frame2_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i118_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38839\,
            in1 => \N__43603\,
            in2 => \_gnd_net_\,
            in3 => \N__50354\,
            lcout => data_out_frame2_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i80_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50359\,
            in1 => \N__40097\,
            in2 => \_gnd_net_\,
            in3 => \N__41149\,
            lcout => data_out_frame2_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i75_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39424\,
            in1 => \N__46594\,
            in2 => \_gnd_net_\,
            in3 => \N__50357\,
            lcout => data_out_frame2_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i79_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50358\,
            in1 => \N__40147\,
            in2 => \_gnd_net_\,
            in3 => \N__40576\,
            lcout => data_out_frame2_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i119_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39704\,
            in1 => \N__43699\,
            in2 => \_gnd_net_\,
            in3 => \N__50355\,
            lcout => data_out_frame2_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15819_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__43602\,
            in1 => \N__46161\,
            in2 => \N__48691\,
            in3 => \N__45410\,
            lcout => \c0.n18681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38369\,
            in2 => \_gnd_net_\,
            in3 => \N__37914\,
            lcout => rand_data_0,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => n16547,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38309\,
            in2 => \_gnd_net_\,
            in3 => \N__37911\,
            lcout => rand_data_1,
            ltout => OPEN,
            carryin => n16547,
            carryout => n16548,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38251\,
            in2 => \_gnd_net_\,
            in3 => \N__37956\,
            lcout => rand_data_2,
            ltout => OPEN,
            carryin => n16548,
            carryout => n16549,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i3_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38164\,
            in2 => \_gnd_net_\,
            in3 => \N__37953\,
            lcout => rand_data_3,
            ltout => OPEN,
            carryin => n16549,
            carryout => n16550,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i4_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38082\,
            in2 => \_gnd_net_\,
            in3 => \N__37950\,
            lcout => rand_data_4,
            ltout => OPEN,
            carryin => n16550,
            carryout => n16551,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i5_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44203\,
            in2 => \_gnd_net_\,
            in3 => \N__37947\,
            lcout => rand_data_5,
            ltout => OPEN,
            carryin => n16551,
            carryout => n16552,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i6_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41258\,
            in2 => \_gnd_net_\,
            in3 => \N__37944\,
            lcout => rand_data_6,
            ltout => OPEN,
            carryin => n16552,
            carryout => n16553,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i7_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42080\,
            in2 => \_gnd_net_\,
            in3 => \N__37941\,
            lcout => rand_data_7,
            ltout => OPEN,
            carryin => n16553,
            carryout => n16554,
            clk => \N__49871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i8_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38693\,
            in2 => \_gnd_net_\,
            in3 => \N__37938\,
            lcout => rand_data_8,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => n16555,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38626\,
            in2 => \_gnd_net_\,
            in3 => \N__37935\,
            lcout => rand_data_9,
            ltout => OPEN,
            carryin => n16555,
            carryout => n16556,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38542\,
            in2 => \_gnd_net_\,
            in3 => \N__37932\,
            lcout => rand_data_10,
            ltout => OPEN,
            carryin => n16556,
            carryout => n16557,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i11_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41446\,
            in2 => \_gnd_net_\,
            in3 => \N__37983\,
            lcout => rand_data_11,
            ltout => OPEN,
            carryin => n16557,
            carryout => n16558,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i12_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50504\,
            in2 => \_gnd_net_\,
            in3 => \N__37980\,
            lcout => rand_data_12,
            ltout => OPEN,
            carryin => n16558,
            carryout => n16559,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i13_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38441\,
            in2 => \_gnd_net_\,
            in3 => \N__37977\,
            lcout => rand_data_13,
            ltout => OPEN,
            carryin => n16559,
            carryout => n16560,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i14_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39265\,
            in2 => \_gnd_net_\,
            in3 => \N__37974\,
            lcout => rand_data_14,
            ltout => OPEN,
            carryin => n16560,
            carryout => n16561,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i15_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39207\,
            in2 => \_gnd_net_\,
            in3 => \N__37971\,
            lcout => rand_data_15,
            ltout => OPEN,
            carryin => n16561,
            carryout => n16562,
            clk => \N__49863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i16_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39135\,
            in2 => \_gnd_net_\,
            in3 => \N__37968\,
            lcout => rand_data_16,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => n16563,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i17_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39055\,
            in2 => \_gnd_net_\,
            in3 => \N__37965\,
            lcout => rand_data_17,
            ltout => OPEN,
            carryin => n16563,
            carryout => n16564,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i18_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40869\,
            in2 => \_gnd_net_\,
            in3 => \N__37962\,
            lcout => rand_data_18,
            ltout => OPEN,
            carryin => n16564,
            carryout => n16565,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i19_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38960\,
            in2 => \_gnd_net_\,
            in3 => \N__37959\,
            lcout => rand_data_19,
            ltout => OPEN,
            carryin => n16565,
            carryout => n16566,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i20_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38891\,
            in2 => \_gnd_net_\,
            in3 => \N__38010\,
            lcout => rand_data_20,
            ltout => OPEN,
            carryin => n16566,
            carryout => n16567,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i21_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38816\,
            in2 => \_gnd_net_\,
            in3 => \N__38007\,
            lcout => rand_data_21,
            ltout => OPEN,
            carryin => n16567,
            carryout => n16568,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i22_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39680\,
            in2 => \_gnd_net_\,
            in3 => \N__38004\,
            lcout => rand_data_22,
            ltout => OPEN,
            carryin => n16568,
            carryout => n16569,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i23_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39602\,
            in2 => \_gnd_net_\,
            in3 => \N__38001\,
            lcout => rand_data_23,
            ltout => OPEN,
            carryin => n16569,
            carryout => n16570,
            clk => \N__49857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i24_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39539\,
            in2 => \_gnd_net_\,
            in3 => \N__37998\,
            lcout => rand_data_24,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => n16571,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i25_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39477\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => rand_data_25,
            ltout => OPEN,
            carryin => n16571,
            carryout => n16572,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i26_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39411\,
            in2 => \_gnd_net_\,
            in3 => \N__37992\,
            lcout => rand_data_26,
            ltout => OPEN,
            carryin => n16572,
            carryout => n16573,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i27_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42128\,
            in2 => \_gnd_net_\,
            in3 => \N__37989\,
            lcout => rand_data_27,
            ltout => OPEN,
            carryin => n16573,
            carryout => n16574,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i28_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41478\,
            in2 => \_gnd_net_\,
            in3 => \N__37986\,
            lcout => rand_data_28,
            ltout => OPEN,
            carryin => n16574,
            carryout => n16575,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i29_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39325\,
            in2 => \_gnd_net_\,
            in3 => \N__38409\,
            lcout => rand_data_29,
            ltout => OPEN,
            carryin => n16575,
            carryout => n16576,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i30_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40125\,
            in2 => \_gnd_net_\,
            in3 => \N__38406\,
            lcout => rand_data_30,
            ltout => OPEN,
            carryin => n16576,
            carryout => n16577,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2481__i31_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40076\,
            in2 => \_gnd_net_\,
            in3 => \N__38403\,
            lcout => rand_data_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i0_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38381\,
            in2 => \N__50945\,
            in3 => \_gnd_net_\,
            lcout => rand_setpoint_0,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => n16578,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38316\,
            in2 => \N__40010\,
            in3 => \N__38280\,
            lcout => rand_setpoint_1,
            ltout => OPEN,
            carryin => n16578,
            carryout => n16579,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38261\,
            in2 => \N__38207\,
            in3 => \N__38190\,
            lcout => rand_setpoint_2,
            ltout => OPEN,
            carryin => n16579,
            carryout => n16580,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i3_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38175\,
            in2 => \N__38129\,
            in3 => \N__38112\,
            lcout => rand_setpoint_3,
            ltout => OPEN,
            carryin => n16580,
            carryout => n16581,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i4_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38048\,
            in2 => \N__38090\,
            in3 => \N__38037\,
            lcout => rand_setpoint_4,
            ltout => OPEN,
            carryin => n16581,
            carryout => n16582,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i5_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38024\,
            in2 => \N__44228\,
            in3 => \N__38013\,
            lcout => rand_setpoint_5,
            ltout => OPEN,
            carryin => n16582,
            carryout => n16583,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i6_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38762\,
            in2 => \N__41280\,
            in3 => \N__38751\,
            lcout => rand_setpoint_6,
            ltout => OPEN,
            carryin => n16583,
            carryout => n16584,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i7_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38738\,
            in2 => \N__42097\,
            in3 => \N__38727\,
            lcout => rand_setpoint_7,
            ltout => OPEN,
            carryin => n16584,
            carryout => n16585,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i8_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38702\,
            in2 => \N__43169\,
            in3 => \N__38664\,
            lcout => rand_setpoint_8,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => n16586,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i9_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38649\,
            in2 => \N__38588\,
            in3 => \N__38571\,
            lcout => rand_setpoint_9,
            ltout => OPEN,
            carryin => n16586,
            carryout => n16587,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i10_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38552\,
            in2 => \N__38508\,
            in3 => \N__38493\,
            lcout => rand_setpoint_10,
            ltout => OPEN,
            carryin => n16587,
            carryout => n16588,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i11_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41453\,
            in2 => \N__42888\,
            in3 => \N__38490\,
            lcout => rand_setpoint_11,
            ltout => OPEN,
            carryin => n16588,
            carryout => n16589,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i12_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50523\,
            in2 => \N__38480\,
            in3 => \N__38463\,
            lcout => rand_setpoint_12,
            ltout => OPEN,
            carryin => n16589,
            carryout => n16590,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i13_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38449\,
            in2 => \N__40040\,
            in3 => \N__38412\,
            lcout => rand_setpoint_13,
            ltout => OPEN,
            carryin => n16590,
            carryout => n16591,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i14_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39283\,
            in2 => \N__47915\,
            in3 => \N__39237\,
            lcout => rand_setpoint_14,
            ltout => OPEN,
            carryin => n16591,
            carryout => n16592,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i15_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39173\,
            in2 => \N__39230\,
            in3 => \N__39162\,
            lcout => rand_setpoint_15,
            ltout => OPEN,
            carryin => n16592,
            carryout => n16593,
            clk => \N__49831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i16_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39148\,
            in2 => \N__39107\,
            in3 => \N__39090\,
            lcout => rand_setpoint_16,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => n16594,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i17_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39070\,
            in2 => \N__39026\,
            in3 => \N__39009\,
            lcout => rand_setpoint_17,
            ltout => OPEN,
            carryin => n16594,
            carryout => n16595,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i18_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40876\,
            in2 => \N__39002\,
            in3 => \N__38985\,
            lcout => rand_setpoint_18,
            ltout => OPEN,
            carryin => n16595,
            carryout => n16596,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i19_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38979\,
            in2 => \N__38927\,
            in3 => \N__38910\,
            lcout => rand_setpoint_19,
            ltout => OPEN,
            carryin => n16596,
            carryout => n16597,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i20_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38906\,
            in2 => \N__38865\,
            in3 => \N__38850\,
            lcout => rand_setpoint_20,
            ltout => OPEN,
            carryin => n16597,
            carryout => n16598,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i21_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38838\,
            in2 => \N__38790\,
            in3 => \N__38775\,
            lcout => rand_setpoint_21,
            ltout => OPEN,
            carryin => n16598,
            carryout => n16599,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i22_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39699\,
            in2 => \N__39653\,
            in3 => \N__39636\,
            lcout => rand_setpoint_22,
            ltout => OPEN,
            carryin => n16599,
            carryout => n16600,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i23_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39624\,
            in2 => \N__39575\,
            in3 => \N__39558\,
            lcout => rand_setpoint_23,
            ltout => OPEN,
            carryin => n16600,
            carryout => n16601,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i24_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39553\,
            in2 => \N__42513\,
            in3 => \N__39513\,
            lcout => rand_setpoint_24,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => n16602,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i25_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39492\,
            in2 => \N__39446\,
            in3 => \N__39429\,
            lcout => rand_setpoint_25,
            ltout => OPEN,
            carryin => n16602,
            carryout => n16603,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i26_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39415\,
            in2 => \N__39854\,
            in3 => \N__39387\,
            lcout => rand_setpoint_26,
            ltout => OPEN,
            carryin => n16603,
            carryout => n16604,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i27_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42138\,
            in2 => \N__39773\,
            in3 => \N__39384\,
            lcout => rand_setpoint_27,
            ltout => OPEN,
            carryin => n16604,
            carryout => n16605,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i28_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41499\,
            in2 => \N__39374\,
            in3 => \N__39357\,
            lcout => rand_setpoint_28,
            ltout => OPEN,
            carryin => n16605,
            carryout => n16606,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i29_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39342\,
            in2 => \N__39306\,
            in3 => \N__39291\,
            lcout => rand_setpoint_29,
            ltout => OPEN,
            carryin => n16606,
            carryout => n16607,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i30_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40146\,
            in2 => \N__39791\,
            in3 => \N__40101\,
            lcout => rand_setpoint_30,
            ltout => OPEN,
            carryin => n16607,
            carryout => n16608,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2482__i31_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40092\,
            in1 => \N__43545\,
            in2 => \_gnd_net_\,
            in3 => \N__40044\,
            lcout => rand_setpoint_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5__2195_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__39931\,
            in1 => \N__40041\,
            in2 => \N__47799\,
            in3 => \N__47886\,
            lcout => \c0.data_out_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15534_3_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__47661\,
            in1 => \N__39743\,
            in2 => \_gnd_net_\,
            in3 => \N__39822\,
            lcout => \c0.n18234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__1__2191_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46814\,
            in1 => \N__40011\,
            in2 => \_gnd_net_\,
            in3 => \N__39972\,
            lcout => \c0.data_out_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_562_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39930\,
            in1 => \N__47735\,
            in2 => \_gnd_net_\,
            in3 => \N__39909\,
            lcout => \c0.n10533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2__2214_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39855\,
            lcout => \c0.data_out_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49783\,
            ce => \N__43418\,
            sr => \N__43477\
        );

    \c0.data_out_5__6__2210_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39792\,
            in2 => \_gnd_net_\,
            in3 => \N__47409\,
            lcout => \c0.data_out_7__2__N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49783\,
            ce => \N__43418\,
            sr => \N__43477\
        );

    \c0.data_out_5__3__2213_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39774\,
            in2 => \_gnd_net_\,
            in3 => \N__47408\,
            lcout => \c0.data_out_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49783\,
            ce => \N__43418\,
            sr => \N__43477\
        );

    \c0.data_out_10__4__2172_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40341\,
            in2 => \_gnd_net_\,
            in3 => \N__40323\,
            lcout => \c0.data_out_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49768\,
            ce => \N__46857\,
            sr => \_gnd_net_\
        );

    \c0.data_out_3__0__2232_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40245\,
            in1 => \N__40281\,
            in2 => \_gnd_net_\,
            in3 => \N__43395\,
            lcout => data_out_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40244\,
            in1 => \N__40226\,
            in2 => \_gnd_net_\,
            in3 => \N__42862\,
            lcout => \c0.n2_adj_2221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__0__2240_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__40227\,
            in1 => \N__43394\,
            in2 => \_gnd_net_\,
            in3 => \N__47141\,
            lcout => data_out_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_15_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__46164\,
            in1 => \N__40218\,
            in2 => \N__48702\,
            in3 => \N__41568\,
            lcout => \c0.n6_adj_2227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15874_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__41763\,
            in1 => \N__43708\,
            in2 => \N__48700\,
            in3 => \N__46163\,
            lcout => \c0.n18705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_810_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45305\,
            in1 => \N__40949\,
            in2 => \_gnd_net_\,
            in3 => \N__40203\,
            lcout => \c0.n17899\,
            ltout => \c0.n17899_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_738_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41864\,
            in1 => \N__44010\,
            in2 => \N__40167\,
            in3 => \N__42180\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_796_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40840\,
            in2 => \_gnd_net_\,
            in3 => \N__44324\,
            lcout => \c0.n17736\,
            ltout => \c0.n17736_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_541_LC_15_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41863\,
            in1 => \N__41218\,
            in2 => \N__40611\,
            in3 => \N__40587\,
            lcout => \c0.n17914\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18813_bdd_4_lut_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__42231\,
            in1 => \N__44268\,
            in2 => \N__48701\,
            in3 => \N__40608\,
            lcout => \c0.n18816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_501_LC_15_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44325\,
            in1 => \_gnd_net_\,
            in2 => \N__40845\,
            in3 => \N__40588\,
            lcout => \c0.n10725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_683_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40549\,
            in1 => \N__41883\,
            in2 => \N__40509\,
            in3 => \N__46308\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i163_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43979\,
            in1 => \N__40491\,
            in2 => \N__40479\,
            in3 => \N__40371\,
            lcout => \c0.data_out_frame2_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49888\,
            ce => \N__50462\,
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_681_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40476\,
            in1 => \N__45267\,
            in2 => \N__40436\,
            in3 => \N__40407\,
            lcout => \c0.n17862\,
            ltout => \c0.n17862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_676_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40905\,
            in1 => \N__45536\,
            in2 => \N__40365\,
            in3 => \N__40362\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i164_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41679\,
            in1 => \N__50553\,
            in2 => \N__40344\,
            in3 => \N__43776\,
            lcout => \c0.data_out_frame2_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49888\,
            ce => \N__50462\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_719_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40992\,
            in2 => \_gnd_net_\,
            in3 => \N__40950\,
            lcout => \c0.n17889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_790_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41145\,
            lcout => \c0.n17868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i51_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40892\,
            in1 => \N__40839\,
            in2 => \_gnd_net_\,
            in3 => \N__50436\,
            lcout => data_out_frame2_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18645_bdd_4_lut_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__43761\,
            in1 => \N__48686\,
            in2 => \N__46595\,
            in3 => \N__40815\,
            lcout => \c0.n18648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_770_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45814\,
            in1 => \N__41331\,
            in2 => \N__44535\,
            in3 => \N__40787\,
            lcout => \c0.n18_adj_2441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18663_bdd_4_lut_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__40786\,
            in1 => \N__41376\,
            in2 => \N__44581\,
            in3 => \N__48685\,
            lcout => \c0.n18666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_520_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__43610\,
            in1 => \_gnd_net_\,
            in2 => \N__43679\,
            in3 => \N__40752\,
            lcout => \c0.n17917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_740_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40707\,
            in1 => \N__40688\,
            in2 => \N__41523\,
            in3 => \N__44523\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46191\,
            in1 => \N__40665\,
            in2 => \_gnd_net_\,
            in3 => \N__44690\,
            lcout => \c0.n5_adj_2439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15804_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__45625\,
            in1 => \N__41414\,
            in2 => \N__48693\,
            in3 => \N__46192\,
            lcout => \c0.n18663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_769_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41370\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45015\,
            lcout => \c0.n10911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_772_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50571\,
            in1 => \N__45244\,
            in2 => \_gnd_net_\,
            in3 => \N__41312\,
            lcout => \c0.n17810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i103_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41262\,
            in1 => \N__43579\,
            in2 => \_gnd_net_\,
            in3 => \N__50446\,
            lcout => data_out_frame2_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i77_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50447\,
            in1 => \N__41507\,
            in2 => \_gnd_net_\,
            in3 => \N__41217\,
            lcout => data_out_frame2_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_812_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41185\,
            in1 => \N__44053\,
            in2 => \N__41150\,
            in3 => \N__44614\,
            lcout => \c0.n10703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i93_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50448\,
            in1 => \_gnd_net_\,
            in2 => \N__50581\,
            in3 => \N__50525\,
            lcout => data_out_frame2_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_542_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46590\,
            in1 => \N__46707\,
            in2 => \N__41121\,
            in3 => \N__43575\,
            lcout => \c0.n14_adj_2362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_522_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46411\,
            in1 => \N__41567\,
            in2 => \N__41094\,
            in3 => \N__41037\,
            lcout => \c0.n17892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_728_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46589\,
            in1 => \N__41901\,
            in2 => \_gnd_net_\,
            in3 => \N__41765\,
            lcout => \c0.n17789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__41859\,
            in1 => \N__48609\,
            in2 => \N__41826\,
            in3 => \N__46193\,
            lcout => \c0.n6_adj_2218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_adj_646_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41816\,
            in2 => \_gnd_net_\,
            in3 => \N__41764\,
            lcout => \c0.n18_adj_2393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_730_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41723\,
            in1 => \N__41670\,
            in2 => \N__41625\,
            in3 => \N__50821\,
            lcout => \c0.n10_adj_2431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__46194\,
            in1 => \N__44067\,
            in2 => \N__48684\,
            in3 => \N__43855\,
            lcout => \c0.n6_adj_2360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_766_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41566\,
            in2 => \_gnd_net_\,
            in3 => \N__50881\,
            lcout => \c0.n17865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i109_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41500\,
            in1 => \N__42969\,
            in2 => \_gnd_net_\,
            in3 => \N__50453\,
            lcout => data_out_frame2_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i140_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50454\,
            in1 => \N__41447\,
            in2 => \_gnd_net_\,
            in3 => \N__41973\,
            lcout => data_out_frame2_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_696_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42230\,
            in2 => \_gnd_net_\,
            in3 => \N__41954\,
            lcout => \c0.n17902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_679_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__42201\,
            in1 => \N__44754\,
            in2 => \_gnd_net_\,
            in3 => \N__50820\,
            lcout => \c0.n10583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18705_bdd_4_lut_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__48607\,
            in1 => \N__42192\,
            in2 => \N__43584\,
            in3 => \N__42173\,
            lcout => \c0.n18708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i76_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50455\,
            in1 => \N__42149\,
            in2 => \_gnd_net_\,
            in3 => \N__44571\,
            lcout => data_out_frame2_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i104_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42087\,
            in1 => \N__44267\,
            in2 => \_gnd_net_\,
            in3 => \N__50452\,
            lcout => data_out_frame2_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18657_bdd_4_lut_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__42053\,
            in1 => \N__48608\,
            in2 => \N__43821\,
            in3 => \N__42015\,
            lcout => \c0.n18660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15794_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42003\,
            in1 => \N__48618\,
            in2 => \N__41985\,
            in3 => \N__46159\,
            lcout => OPEN,
            ltout => \c0.n18651_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18651_bdd_4_lut_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48619\,
            in1 => \N__41972\,
            in2 => \N__41961\,
            in3 => \N__41958\,
            lcout => OPEN,
            ltout => \c0.n18654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__48076\,
            in1 => \N__41916\,
            in2 => \N__41904\,
            in3 => \N__48139\,
            lcout => \c0.n22_adj_2259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15859_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42438\,
            in1 => \N__49097\,
            in2 => \N__42429\,
            in3 => \N__48077\,
            lcout => OPEN,
            ltout => \c0.n18735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18735_bdd_4_lut_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49098\,
            in1 => \N__42417\,
            in2 => \N__42408\,
            in3 => \N__42405\,
            lcout => OPEN,
            ltout => \c0.n18738_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__42396\,
            in1 => \N__49099\,
            in2 => \N__42390\,
            in3 => \N__48950\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49864\,
            ce => \N__48828\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15833_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__46150\,
            in1 => \N__42372\,
            in2 => \N__43881\,
            in3 => \N__48402\,
            lcout => \c0.n18699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15943_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__42354\,
            in1 => \N__49094\,
            in2 => \N__42345\,
            in3 => \N__48079\,
            lcout => OPEN,
            ltout => \c0.n18777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18777_bdd_4_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49095\,
            in1 => \N__42327\,
            in2 => \N__42315\,
            in3 => \N__42312\,
            lcout => \c0.n18780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18699_bdd_4_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__48403\,
            in1 => \N__42303\,
            in2 => \N__42297\,
            in3 => \N__42276\,
            lcout => OPEN,
            ltout => \c0.n18702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__48080\,
            in1 => \N__44469\,
            in2 => \N__42234\,
            in3 => \N__48138\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__43002\,
            in1 => \N__49096\,
            in2 => \N__42996\,
            in3 => \N__48949\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49858\,
            ce => \N__48824\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15899_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__48620\,
            in1 => \N__46080\,
            in2 => \N__44439\,
            in3 => \N__45013\,
            lcout => OPEN,
            ltout => \c0.n18783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18783_bdd_4_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__45201\,
            in1 => \N__48621\,
            in2 => \N__42981\,
            in3 => \N__42976\,
            lcout => \c0.n18161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11016_2_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47399\,
            in2 => \_gnd_net_\,
            in3 => \N__47129\,
            lcout => n2732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15645_2_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42933\,
            in2 => \_gnd_net_\,
            in3 => \N__42863\,
            lcout => \c0.n18311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15532_2_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42887\,
            in2 => \_gnd_net_\,
            in3 => \N__47404\,
            lcout => \c0.n18201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42864\,
            in1 => \N__42524\,
            in2 => \_gnd_net_\,
            in3 => \N__42604\,
            lcout => \c0.n5_adj_2217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__3__2197_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__47671\,
            in1 => \N__47130\,
            in2 => \N__42549\,
            in3 => \N__43514\,
            lcout => \c0.data_out_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49820\,
            ce => \N__47893\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__0__2216_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42512\,
            in2 => \_gnd_net_\,
            in3 => \N__47405\,
            lcout => \c0.data_out_6__1__N_537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49809\,
            ce => \N__43417\,
            sr => \N__43479\
        );

    \c0.data_out_5__7__2209_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43544\,
            lcout => \c0.data_out_7__3__N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49809\,
            ce => \N__43417\,
            sr => \N__43479\
        );

    \c0.data_out_1__1__2247_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__47676\,
            in1 => \N__47410\,
            in2 => \_gnd_net_\,
            in3 => \N__47144\,
            lcout => \c0.data_out_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49797\,
            ce => \N__43419\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0__2200_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__43185\,
            in1 => \N__47411\,
            in2 => \N__43176\,
            in3 => \N__47145\,
            lcout => \c0.data_out_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49784\,
            ce => \N__47884\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15884_LC_16_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__43122\,
            in1 => \N__49108\,
            in2 => \N__43113\,
            in3 => \N__48071\,
            lcout => OPEN,
            ltout => \c0.n18765_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18765_bdd_4_lut_LC_16_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49109\,
            in1 => \N__43101\,
            in2 => \N__43089\,
            in3 => \N__43086\,
            lcout => OPEN,
            ltout => \c0.n18768_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_16_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__43989\,
            in1 => \N__49110\,
            in2 => \N__43077\,
            in3 => \N__48951\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49892\,
            ce => \N__48811\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15779_LC_16_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__43056\,
            in1 => \N__48679\,
            in2 => \N__43038\,
            in3 => \N__46184\,
            lcout => OPEN,
            ltout => \c0.n18633_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18633_bdd_4_lut_LC_16_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48680\,
            in1 => \N__43026\,
            in2 => \N__43005\,
            in3 => \N__46654\,
            lcout => OPEN,
            ltout => \c0.n18636_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_16_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__48070\,
            in1 => \N__43998\,
            in2 => \N__43992\,
            in3 => \N__48169\,
            lcout => \c0.n22_adj_2268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_753_LC_16_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50763\,
            in1 => \N__43583\,
            in2 => \N__43983\,
            in3 => \N__43959\,
            lcout => OPEN,
            ltout => \c0.n20_adj_2438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i159_LC_16_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43911\,
            in1 => \N__43767\,
            in2 => \N__43902\,
            in3 => \N__43899\,
            lcout => \c0.data_out_frame2_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => \N__50475\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_750_LC_16_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__43866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43820\,
            lcout => \c0.n10905\,
            ltout => \c0.n10905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_4_lut_LC_16_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44150\,
            in1 => \N__44284\,
            in2 => \N__43770\,
            in3 => \N__46486\,
            lcout => \c0.n16_adj_2391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_801_LC_16_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43710\,
            in1 => \N__43760\,
            in2 => \_gnd_net_\,
            in3 => \N__45790\,
            lcout => \c0.n17920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_427_LC_16_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43709\,
            lcout => \c0.n10788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_756_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__43680\,
            in1 => \N__43614\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_767_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43574\,
            in2 => \_gnd_net_\,
            in3 => \N__48221\,
            lcout => \c0.n10929\,
            ltout => \c0.n10929_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_734_LC_16_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44857\,
            in2 => \N__44526\,
            in3 => \N__44928\,
            lcout => \c0.n17823\,
            ltout => \c0.n17823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_656_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44433\,
            in1 => \N__44517\,
            in2 => \N__44502\,
            in3 => \N__46485\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i167_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44499\,
            in1 => \N__46545\,
            in2 => \N__44493\,
            in3 => \N__44489\,
            lcout => \c0.data_out_frame2_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => \N__50466\,
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_660_LC_16_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44453\,
            in1 => \N__44582\,
            in2 => \N__44438\,
            in3 => \N__44388\,
            lcout => \c0.n18_adj_2402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_649_LC_16_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44376\,
            in1 => \N__44331\,
            in2 => \N__44285\,
            in3 => \N__44858\,
            lcout => \c0.n22_adj_2395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i102_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44140\,
            in1 => \N__44230\,
            in2 => \_gnd_net_\,
            in3 => \N__50449\,
            lcout => data_out_frame2_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45115\,
            in1 => \N__44103\,
            in2 => \_gnd_net_\,
            in3 => \N__46196\,
            lcout => \c0.n5_adj_2381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_735_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44900\,
            in1 => \N__46416\,
            in2 => \N__44061\,
            in3 => \N__45117\,
            lcout => \c0.n30_adj_2434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_667_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45116\,
            in1 => \N__45093\,
            in2 => \_gnd_net_\,
            in3 => \N__45045\,
            lcout => \c0.n17871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_733_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46353\,
            in1 => \N__45014\,
            in2 => \N__44971\,
            in3 => \N__45546\,
            lcout => \c0.n10710\,
            ltout => \c0.n10710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_662_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44718\,
            in1 => \N__45287\,
            in2 => \N__44922\,
            in3 => \N__44919\,
            lcout => \c0.n20_adj_2404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46195\,
            in1 => \N__44901\,
            in2 => \_gnd_net_\,
            in3 => \N__44859\,
            lcout => \c0.n5_adj_2386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_764_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44811\,
            in2 => \_gnd_net_\,
            in3 => \N__44753\,
            lcout => \c0.n10877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_711_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45668\,
            in1 => \N__45621\,
            in2 => \_gnd_net_\,
            in3 => \N__45683\,
            lcout => OPEN,
            ltout => \c0.n10593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45380\,
            in2 => \N__44712\,
            in3 => \N__44697\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_729_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44696\,
            in1 => \N__44661\,
            in2 => \N__44625\,
            in3 => \N__44564\,
            lcout => \c0.n17751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_534_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45682\,
            in1 => \N__45667\,
            in2 => \N__45626\,
            in3 => \N__45576\,
            lcout => \c0.n17798\,
            ltout => \c0.n17798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_648_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45523\,
            in1 => \N__45507\,
            in2 => \N__45489\,
            in3 => \N__45482\,
            lcout => OPEN,
            ltout => \c0.n24_adj_2394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_651_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45468\,
            in1 => \N__45462\,
            in2 => \N__45417\,
            in3 => \N__45414\,
            lcout => OPEN,
            ltout => \c0.n26_adj_2396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i168_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45381\,
            in1 => \N__45369\,
            in2 => \N__45360\,
            in3 => \N__45353\,
            lcout => \c0.data_out_frame2_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49882\,
            ce => \N__50469\,
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_668_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__46656\,
            in1 => \_gnd_net_\,
            in2 => \N__50552\,
            in3 => \N__45315\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i165_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45288\,
            in1 => \N__46662\,
            in2 => \N__45270\,
            in3 => \N__45123\,
            lcout => \c0.data_out_frame2_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__50468\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_670_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45263\,
            in1 => \N__45249\,
            in2 => \N__45207\,
            in3 => \N__45147\,
            lcout => \c0.n15_adj_2407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_685_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46715\,
            in2 => \_gnd_net_\,
            in3 => \N__46604\,
            lcout => \c0.n17856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_654_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46655\,
            in1 => \N__46536\,
            in2 => \N__46608\,
            in3 => \N__46563\,
            lcout => \c0.n16_adj_2399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15988_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__48694\,
            in1 => \N__46533\,
            in2 => \N__46488\,
            in3 => \N__46157\,
            lcout => OPEN,
            ltout => \c0.n18891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18891_bdd_4_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48692\,
            in1 => \N__46410\,
            in2 => \N__46356\,
            in3 => \N__46352\,
            lcout => \c0.n18060\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__48695\,
            in1 => \N__46304\,
            in2 => \N__46263\,
            in3 => \N__46158\,
            lcout => OPEN,
            ltout => \c0.n18897_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18897_bdd_4_lut_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__45857\,
            in1 => \N__48696\,
            in2 => \N__45819\,
            in3 => \N__45816\,
            lcout => OPEN,
            ltout => \c0.n18057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15854_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__45732\,
            in1 => \N__49111\,
            in2 => \N__45726\,
            in3 => \N__48081\,
            lcout => OPEN,
            ltout => \c0.n18723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18723_bdd_4_lut_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49112\,
            in1 => \N__45723\,
            in2 => \N__45714\,
            in3 => \N__45711\,
            lcout => OPEN,
            ltout => \c0.n18726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__49200\,
            in1 => \N__49113\,
            in2 => \N__49182\,
            in3 => \N__48948\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49873\,
            ce => \N__48816\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15889_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__49170\,
            in1 => \N__48078\,
            in2 => \N__49158\,
            in3 => \N__49114\,
            lcout => OPEN,
            ltout => \c0.n18771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18771_bdd_4_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49115\,
            in1 => \N__49149\,
            in2 => \N__49131\,
            in3 => \N__49128\,
            lcout => OPEN,
            ltout => \c0.n18774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__47925\,
            in1 => \N__49116\,
            in2 => \N__48954\,
            in3 => \N__48947\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49865\,
            ce => \N__48823\,
            sr => \_gnd_net_\
        );

    \c0.n18669_bdd_4_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__48717\,
            in1 => \N__48705\,
            in2 => \N__49914\,
            in3 => \N__48222\,
            lcout => OPEN,
            ltout => \c0.n18672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__48180\,
            in1 => \N__48157\,
            in2 => \N__48084\,
            in3 => \N__48075\,
            lcout => \c0.n22_adj_2243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6__2194_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__47919\,
            in1 => \N__47894\,
            in2 => \N__47791\,
            in3 => \N__47723\,
            lcout => \c0.data_out_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15718_2_lut_3_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47633\,
            in1 => \N__47403\,
            in2 => \_gnd_net_\,
            in3 => \N__47143\,
            lcout => \data_out_10__7__N_110\,
            ltout => \data_out_10__7__N_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__0__2192_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50949\,
            in2 => \N__50928\,
            in3 => \N__50910\,
            lcout => data_out_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_752_LC_17_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50757\,
            in1 => \N__50886\,
            in2 => \N__50832\,
            in3 => \N__50822\,
            lcout => \c0.n18_adj_2437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_674_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50756\,
            in2 => \_gnd_net_\,
            in3 => \N__50712\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_675_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50676\,
            in1 => \N__50625\,
            in2 => \N__50589\,
            in3 => \N__50585\,
            lcout => \c0.n17905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i141_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50524\,
            in1 => \N__49907\,
            in2 => \_gnd_net_\,
            in3 => \N__50450\,
            lcout => data_out_frame2_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
