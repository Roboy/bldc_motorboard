// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 16 2019 18:45:02

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    inout PIN_6;
    inout PIN_5;
    inout PIN_4;
    output PIN_3;
    output PIN_24;
    output PIN_23;
    output PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    inout PIN_11;
    inout PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__73031;
    wire N__73030;
    wire N__73029;
    wire N__73022;
    wire N__73021;
    wire N__73020;
    wire N__73013;
    wire N__73012;
    wire N__73011;
    wire N__73004;
    wire N__73003;
    wire N__73002;
    wire N__72995;
    wire N__72994;
    wire N__72993;
    wire N__72986;
    wire N__72985;
    wire N__72984;
    wire N__72977;
    wire N__72976;
    wire N__72975;
    wire N__72968;
    wire N__72967;
    wire N__72966;
    wire N__72959;
    wire N__72958;
    wire N__72957;
    wire N__72950;
    wire N__72949;
    wire N__72948;
    wire N__72941;
    wire N__72940;
    wire N__72939;
    wire N__72932;
    wire N__72931;
    wire N__72930;
    wire N__72923;
    wire N__72922;
    wire N__72921;
    wire N__72914;
    wire N__72913;
    wire N__72912;
    wire N__72905;
    wire N__72904;
    wire N__72903;
    wire N__72896;
    wire N__72895;
    wire N__72894;
    wire N__72887;
    wire N__72886;
    wire N__72885;
    wire N__72878;
    wire N__72877;
    wire N__72876;
    wire N__72859;
    wire N__72858;
    wire N__72855;
    wire N__72852;
    wire N__72851;
    wire N__72848;
    wire N__72845;
    wire N__72844;
    wire N__72841;
    wire N__72838;
    wire N__72835;
    wire N__72834;
    wire N__72833;
    wire N__72832;
    wire N__72831;
    wire N__72828;
    wire N__72827;
    wire N__72824;
    wire N__72819;
    wire N__72812;
    wire N__72809;
    wire N__72806;
    wire N__72803;
    wire N__72800;
    wire N__72795;
    wire N__72790;
    wire N__72781;
    wire N__72778;
    wire N__72775;
    wire N__72774;
    wire N__72771;
    wire N__72768;
    wire N__72767;
    wire N__72766;
    wire N__72761;
    wire N__72756;
    wire N__72755;
    wire N__72754;
    wire N__72749;
    wire N__72748;
    wire N__72745;
    wire N__72744;
    wire N__72741;
    wire N__72740;
    wire N__72739;
    wire N__72738;
    wire N__72737;
    wire N__72734;
    wire N__72733;
    wire N__72730;
    wire N__72729;
    wire N__72726;
    wire N__72723;
    wire N__72720;
    wire N__72717;
    wire N__72712;
    wire N__72711;
    wire N__72710;
    wire N__72707;
    wire N__72704;
    wire N__72701;
    wire N__72700;
    wire N__72699;
    wire N__72698;
    wire N__72697;
    wire N__72694;
    wire N__72691;
    wire N__72686;
    wire N__72681;
    wire N__72678;
    wire N__72677;
    wire N__72674;
    wire N__72673;
    wire N__72672;
    wire N__72669;
    wire N__72666;
    wire N__72661;
    wire N__72660;
    wire N__72659;
    wire N__72656;
    wire N__72653;
    wire N__72650;
    wire N__72649;
    wire N__72646;
    wire N__72641;
    wire N__72636;
    wire N__72633;
    wire N__72630;
    wire N__72627;
    wire N__72622;
    wire N__72615;
    wire N__72614;
    wire N__72613;
    wire N__72612;
    wire N__72611;
    wire N__72610;
    wire N__72607;
    wire N__72604;
    wire N__72601;
    wire N__72598;
    wire N__72595;
    wire N__72592;
    wire N__72589;
    wire N__72584;
    wire N__72575;
    wire N__72572;
    wire N__72569;
    wire N__72566;
    wire N__72563;
    wire N__72558;
    wire N__72549;
    wire N__72546;
    wire N__72541;
    wire N__72538;
    wire N__72535;
    wire N__72532;
    wire N__72531;
    wire N__72528;
    wire N__72525;
    wire N__72522;
    wire N__72517;
    wire N__72510;
    wire N__72505;
    wire N__72502;
    wire N__72499;
    wire N__72496;
    wire N__72491;
    wire N__72486;
    wire N__72475;
    wire N__72474;
    wire N__72473;
    wire N__72468;
    wire N__72467;
    wire N__72466;
    wire N__72463;
    wire N__72460;
    wire N__72455;
    wire N__72452;
    wire N__72449;
    wire N__72446;
    wire N__72439;
    wire N__72438;
    wire N__72437;
    wire N__72434;
    wire N__72429;
    wire N__72426;
    wire N__72425;
    wire N__72424;
    wire N__72421;
    wire N__72418;
    wire N__72415;
    wire N__72412;
    wire N__72409;
    wire N__72404;
    wire N__72397;
    wire N__72394;
    wire N__72393;
    wire N__72392;
    wire N__72389;
    wire N__72386;
    wire N__72385;
    wire N__72382;
    wire N__72379;
    wire N__72376;
    wire N__72373;
    wire N__72370;
    wire N__72369;
    wire N__72366;
    wire N__72359;
    wire N__72356;
    wire N__72349;
    wire N__72346;
    wire N__72343;
    wire N__72342;
    wire N__72339;
    wire N__72338;
    wire N__72337;
    wire N__72336;
    wire N__72335;
    wire N__72332;
    wire N__72329;
    wire N__72324;
    wire N__72319;
    wire N__72316;
    wire N__72309;
    wire N__72304;
    wire N__72301;
    wire N__72298;
    wire N__72295;
    wire N__72294;
    wire N__72293;
    wire N__72292;
    wire N__72291;
    wire N__72288;
    wire N__72287;
    wire N__72286;
    wire N__72285;
    wire N__72284;
    wire N__72283;
    wire N__72280;
    wire N__72277;
    wire N__72274;
    wire N__72271;
    wire N__72270;
    wire N__72267;
    wire N__72262;
    wire N__72261;
    wire N__72260;
    wire N__72257;
    wire N__72256;
    wire N__72255;
    wire N__72254;
    wire N__72251;
    wire N__72248;
    wire N__72243;
    wire N__72242;
    wire N__72241;
    wire N__72238;
    wire N__72235;
    wire N__72232;
    wire N__72231;
    wire N__72228;
    wire N__72225;
    wire N__72222;
    wire N__72221;
    wire N__72218;
    wire N__72217;
    wire N__72214;
    wire N__72211;
    wire N__72208;
    wire N__72207;
    wire N__72206;
    wire N__72205;
    wire N__72202;
    wire N__72201;
    wire N__72200;
    wire N__72199;
    wire N__72196;
    wire N__72193;
    wire N__72190;
    wire N__72187;
    wire N__72184;
    wire N__72181;
    wire N__72178;
    wire N__72175;
    wire N__72172;
    wire N__72165;
    wire N__72162;
    wire N__72159;
    wire N__72156;
    wire N__72153;
    wire N__72150;
    wire N__72149;
    wire N__72146;
    wire N__72145;
    wire N__72144;
    wire N__72141;
    wire N__72136;
    wire N__72133;
    wire N__72132;
    wire N__72129;
    wire N__72128;
    wire N__72125;
    wire N__72122;
    wire N__72117;
    wire N__72114;
    wire N__72105;
    wire N__72100;
    wire N__72097;
    wire N__72092;
    wire N__72085;
    wire N__72082;
    wire N__72079;
    wire N__72074;
    wire N__72071;
    wire N__72066;
    wire N__72059;
    wire N__72054;
    wire N__72051;
    wire N__72046;
    wire N__72043;
    wire N__72036;
    wire N__72031;
    wire N__72024;
    wire N__72019;
    wire N__72014;
    wire N__72009;
    wire N__71998;
    wire N__71995;
    wire N__71994;
    wire N__71993;
    wire N__71992;
    wire N__71989;
    wire N__71982;
    wire N__71977;
    wire N__71974;
    wire N__71973;
    wire N__71972;
    wire N__71971;
    wire N__71970;
    wire N__71969;
    wire N__71966;
    wire N__71965;
    wire N__71964;
    wire N__71963;
    wire N__71962;
    wire N__71961;
    wire N__71960;
    wire N__71959;
    wire N__71958;
    wire N__71955;
    wire N__71952;
    wire N__71949;
    wire N__71948;
    wire N__71947;
    wire N__71942;
    wire N__71941;
    wire N__71938;
    wire N__71935;
    wire N__71934;
    wire N__71933;
    wire N__71932;
    wire N__71929;
    wire N__71922;
    wire N__71917;
    wire N__71912;
    wire N__71907;
    wire N__71902;
    wire N__71899;
    wire N__71898;
    wire N__71895;
    wire N__71890;
    wire N__71883;
    wire N__71876;
    wire N__71871;
    wire N__71870;
    wire N__71869;
    wire N__71868;
    wire N__71863;
    wire N__71860;
    wire N__71857;
    wire N__71854;
    wire N__71851;
    wire N__71846;
    wire N__71839;
    wire N__71836;
    wire N__71833;
    wire N__71830;
    wire N__71825;
    wire N__71822;
    wire N__71817;
    wire N__71806;
    wire N__71803;
    wire N__71802;
    wire N__71801;
    wire N__71800;
    wire N__71797;
    wire N__71794;
    wire N__71793;
    wire N__71792;
    wire N__71791;
    wire N__71788;
    wire N__71787;
    wire N__71786;
    wire N__71783;
    wire N__71782;
    wire N__71781;
    wire N__71780;
    wire N__71779;
    wire N__71778;
    wire N__71777;
    wire N__71776;
    wire N__71775;
    wire N__71770;
    wire N__71767;
    wire N__71766;
    wire N__71763;
    wire N__71762;
    wire N__71759;
    wire N__71756;
    wire N__71755;
    wire N__71754;
    wire N__71749;
    wire N__71746;
    wire N__71745;
    wire N__71744;
    wire N__71741;
    wire N__71740;
    wire N__71739;
    wire N__71738;
    wire N__71735;
    wire N__71734;
    wire N__71729;
    wire N__71726;
    wire N__71723;
    wire N__71718;
    wire N__71713;
    wire N__71710;
    wire N__71707;
    wire N__71704;
    wire N__71701;
    wire N__71698;
    wire N__71693;
    wire N__71688;
    wire N__71681;
    wire N__71678;
    wire N__71671;
    wire N__71668;
    wire N__71665;
    wire N__71662;
    wire N__71659;
    wire N__71656;
    wire N__71653;
    wire N__71650;
    wire N__71647;
    wire N__71644;
    wire N__71641;
    wire N__71636;
    wire N__71633;
    wire N__71630;
    wire N__71625;
    wire N__71624;
    wire N__71623;
    wire N__71620;
    wire N__71615;
    wire N__71612;
    wire N__71607;
    wire N__71604;
    wire N__71601;
    wire N__71594;
    wire N__71591;
    wire N__71586;
    wire N__71583;
    wire N__71580;
    wire N__71573;
    wire N__71570;
    wire N__71563;
    wire N__71548;
    wire N__71547;
    wire N__71544;
    wire N__71543;
    wire N__71540;
    wire N__71537;
    wire N__71536;
    wire N__71535;
    wire N__71534;
    wire N__71531;
    wire N__71528;
    wire N__71527;
    wire N__71526;
    wire N__71525;
    wire N__71524;
    wire N__71521;
    wire N__71518;
    wire N__71513;
    wire N__71510;
    wire N__71507;
    wire N__71506;
    wire N__71505;
    wire N__71504;
    wire N__71503;
    wire N__71500;
    wire N__71497;
    wire N__71496;
    wire N__71493;
    wire N__71492;
    wire N__71489;
    wire N__71488;
    wire N__71487;
    wire N__71486;
    wire N__71485;
    wire N__71480;
    wire N__71473;
    wire N__71470;
    wire N__71467;
    wire N__71466;
    wire N__71465;
    wire N__71464;
    wire N__71459;
    wire N__71456;
    wire N__71453;
    wire N__71450;
    wire N__71445;
    wire N__71442;
    wire N__71437;
    wire N__71436;
    wire N__71433;
    wire N__71430;
    wire N__71427;
    wire N__71420;
    wire N__71419;
    wire N__71412;
    wire N__71409;
    wire N__71404;
    wire N__71399;
    wire N__71394;
    wire N__71393;
    wire N__71390;
    wire N__71385;
    wire N__71380;
    wire N__71377;
    wire N__71376;
    wire N__71375;
    wire N__71374;
    wire N__71369;
    wire N__71362;
    wire N__71359;
    wire N__71356;
    wire N__71353;
    wire N__71350;
    wire N__71349;
    wire N__71348;
    wire N__71347;
    wire N__71344;
    wire N__71341;
    wire N__71336;
    wire N__71333;
    wire N__71330;
    wire N__71323;
    wire N__71320;
    wire N__71315;
    wire N__71312;
    wire N__71307;
    wire N__71302;
    wire N__71295;
    wire N__71284;
    wire N__71283;
    wire N__71280;
    wire N__71277;
    wire N__71274;
    wire N__71273;
    wire N__71270;
    wire N__71267;
    wire N__71266;
    wire N__71265;
    wire N__71262;
    wire N__71259;
    wire N__71256;
    wire N__71251;
    wire N__71248;
    wire N__71245;
    wire N__71240;
    wire N__71233;
    wire N__71232;
    wire N__71231;
    wire N__71230;
    wire N__71229;
    wire N__71228;
    wire N__71227;
    wire N__71226;
    wire N__71225;
    wire N__71224;
    wire N__71223;
    wire N__71222;
    wire N__71221;
    wire N__71220;
    wire N__71219;
    wire N__71218;
    wire N__71217;
    wire N__71216;
    wire N__71215;
    wire N__71214;
    wire N__71213;
    wire N__71212;
    wire N__71211;
    wire N__71210;
    wire N__71209;
    wire N__71208;
    wire N__71207;
    wire N__71206;
    wire N__71205;
    wire N__71204;
    wire N__71203;
    wire N__71202;
    wire N__71201;
    wire N__71200;
    wire N__71199;
    wire N__71198;
    wire N__71197;
    wire N__71196;
    wire N__71195;
    wire N__71194;
    wire N__71193;
    wire N__71192;
    wire N__71191;
    wire N__71190;
    wire N__71189;
    wire N__71188;
    wire N__71187;
    wire N__71186;
    wire N__71185;
    wire N__71184;
    wire N__71183;
    wire N__71182;
    wire N__71181;
    wire N__71180;
    wire N__71179;
    wire N__71178;
    wire N__71177;
    wire N__71176;
    wire N__71175;
    wire N__71174;
    wire N__71173;
    wire N__71172;
    wire N__71171;
    wire N__71170;
    wire N__71169;
    wire N__71168;
    wire N__71167;
    wire N__71166;
    wire N__71165;
    wire N__71164;
    wire N__71163;
    wire N__71162;
    wire N__71161;
    wire N__71160;
    wire N__71159;
    wire N__71158;
    wire N__71157;
    wire N__71156;
    wire N__71155;
    wire N__71154;
    wire N__71153;
    wire N__71152;
    wire N__71151;
    wire N__71150;
    wire N__71149;
    wire N__71148;
    wire N__71147;
    wire N__71146;
    wire N__71145;
    wire N__71144;
    wire N__71143;
    wire N__71142;
    wire N__71141;
    wire N__71140;
    wire N__71139;
    wire N__71138;
    wire N__71137;
    wire N__71136;
    wire N__71135;
    wire N__71134;
    wire N__71133;
    wire N__71132;
    wire N__71131;
    wire N__71130;
    wire N__71129;
    wire N__71128;
    wire N__71127;
    wire N__71126;
    wire N__71125;
    wire N__71124;
    wire N__71123;
    wire N__71122;
    wire N__71121;
    wire N__71120;
    wire N__71119;
    wire N__71118;
    wire N__71117;
    wire N__71116;
    wire N__71115;
    wire N__71114;
    wire N__71113;
    wire N__71112;
    wire N__71111;
    wire N__71110;
    wire N__71109;
    wire N__71108;
    wire N__71107;
    wire N__71106;
    wire N__71105;
    wire N__71104;
    wire N__71103;
    wire N__71102;
    wire N__71101;
    wire N__71100;
    wire N__71099;
    wire N__71098;
    wire N__71097;
    wire N__71096;
    wire N__71095;
    wire N__71094;
    wire N__71093;
    wire N__71092;
    wire N__71091;
    wire N__71090;
    wire N__71089;
    wire N__71088;
    wire N__71087;
    wire N__71086;
    wire N__71085;
    wire N__71084;
    wire N__71083;
    wire N__71082;
    wire N__71081;
    wire N__71080;
    wire N__71079;
    wire N__71078;
    wire N__71077;
    wire N__71076;
    wire N__71075;
    wire N__71074;
    wire N__71073;
    wire N__71072;
    wire N__71071;
    wire N__71070;
    wire N__71069;
    wire N__71068;
    wire N__71067;
    wire N__71066;
    wire N__71065;
    wire N__71064;
    wire N__71063;
    wire N__71062;
    wire N__71061;
    wire N__71060;
    wire N__71059;
    wire N__71058;
    wire N__71057;
    wire N__71056;
    wire N__71055;
    wire N__71054;
    wire N__71053;
    wire N__71052;
    wire N__71051;
    wire N__71050;
    wire N__71049;
    wire N__71048;
    wire N__71047;
    wire N__71046;
    wire N__71045;
    wire N__71044;
    wire N__71043;
    wire N__71042;
    wire N__71041;
    wire N__71040;
    wire N__71039;
    wire N__71038;
    wire N__71037;
    wire N__71036;
    wire N__71035;
    wire N__71034;
    wire N__71033;
    wire N__71032;
    wire N__71031;
    wire N__71030;
    wire N__71029;
    wire N__71028;
    wire N__71027;
    wire N__71026;
    wire N__71025;
    wire N__71024;
    wire N__71023;
    wire N__71022;
    wire N__71021;
    wire N__71020;
    wire N__71019;
    wire N__71018;
    wire N__71017;
    wire N__71016;
    wire N__71015;
    wire N__71014;
    wire N__71013;
    wire N__71012;
    wire N__71011;
    wire N__71010;
    wire N__71009;
    wire N__71008;
    wire N__71007;
    wire N__71006;
    wire N__71005;
    wire N__71004;
    wire N__71003;
    wire N__71002;
    wire N__71001;
    wire N__71000;
    wire N__70999;
    wire N__70998;
    wire N__70997;
    wire N__70996;
    wire N__70995;
    wire N__70994;
    wire N__70993;
    wire N__70992;
    wire N__70991;
    wire N__70504;
    wire N__70501;
    wire N__70498;
    wire N__70495;
    wire N__70494;
    wire N__70491;
    wire N__70488;
    wire N__70485;
    wire N__70482;
    wire N__70481;
    wire N__70478;
    wire N__70475;
    wire N__70472;
    wire N__70465;
    wire N__70464;
    wire N__70461;
    wire N__70460;
    wire N__70457;
    wire N__70456;
    wire N__70451;
    wire N__70448;
    wire N__70445;
    wire N__70442;
    wire N__70439;
    wire N__70438;
    wire N__70435;
    wire N__70432;
    wire N__70429;
    wire N__70428;
    wire N__70425;
    wire N__70420;
    wire N__70417;
    wire N__70414;
    wire N__70405;
    wire N__70402;
    wire N__70399;
    wire N__70396;
    wire N__70393;
    wire N__70390;
    wire N__70389;
    wire N__70386;
    wire N__70383;
    wire N__70382;
    wire N__70379;
    wire N__70376;
    wire N__70375;
    wire N__70374;
    wire N__70371;
    wire N__70368;
    wire N__70365;
    wire N__70362;
    wire N__70359;
    wire N__70354;
    wire N__70351;
    wire N__70348;
    wire N__70339;
    wire N__70338;
    wire N__70337;
    wire N__70334;
    wire N__70331;
    wire N__70328;
    wire N__70325;
    wire N__70324;
    wire N__70321;
    wire N__70318;
    wire N__70315;
    wire N__70314;
    wire N__70311;
    wire N__70308;
    wire N__70303;
    wire N__70300;
    wire N__70291;
    wire N__70288;
    wire N__70285;
    wire N__70282;
    wire N__70279;
    wire N__70276;
    wire N__70273;
    wire N__70270;
    wire N__70267;
    wire N__70264;
    wire N__70261;
    wire N__70258;
    wire N__70257;
    wire N__70254;
    wire N__70251;
    wire N__70248;
    wire N__70243;
    wire N__70242;
    wire N__70239;
    wire N__70236;
    wire N__70233;
    wire N__70230;
    wire N__70225;
    wire N__70224;
    wire N__70221;
    wire N__70218;
    wire N__70213;
    wire N__70210;
    wire N__70209;
    wire N__70208;
    wire N__70205;
    wire N__70202;
    wire N__70199;
    wire N__70196;
    wire N__70189;
    wire N__70188;
    wire N__70183;
    wire N__70180;
    wire N__70177;
    wire N__70174;
    wire N__70171;
    wire N__70168;
    wire N__70165;
    wire N__70162;
    wire N__70161;
    wire N__70158;
    wire N__70155;
    wire N__70154;
    wire N__70151;
    wire N__70148;
    wire N__70147;
    wire N__70144;
    wire N__70139;
    wire N__70134;
    wire N__70131;
    wire N__70126;
    wire N__70125;
    wire N__70124;
    wire N__70123;
    wire N__70120;
    wire N__70117;
    wire N__70114;
    wire N__70111;
    wire N__70108;
    wire N__70105;
    wire N__70102;
    wire N__70099;
    wire N__70096;
    wire N__70091;
    wire N__70084;
    wire N__70083;
    wire N__70080;
    wire N__70077;
    wire N__70074;
    wire N__70069;
    wire N__70066;
    wire N__70063;
    wire N__70060;
    wire N__70057;
    wire N__70056;
    wire N__70053;
    wire N__70050;
    wire N__70045;
    wire N__70044;
    wire N__70041;
    wire N__70038;
    wire N__70037;
    wire N__70032;
    wire N__70029;
    wire N__70026;
    wire N__70021;
    wire N__70018;
    wire N__70017;
    wire N__70016;
    wire N__70013;
    wire N__70010;
    wire N__70007;
    wire N__70004;
    wire N__70001;
    wire N__69998;
    wire N__69991;
    wire N__69988;
    wire N__69987;
    wire N__69986;
    wire N__69983;
    wire N__69980;
    wire N__69977;
    wire N__69974;
    wire N__69971;
    wire N__69968;
    wire N__69967;
    wire N__69966;
    wire N__69965;
    wire N__69964;
    wire N__69961;
    wire N__69958;
    wire N__69955;
    wire N__69946;
    wire N__69937;
    wire N__69934;
    wire N__69933;
    wire N__69930;
    wire N__69927;
    wire N__69922;
    wire N__69919;
    wire N__69918;
    wire N__69913;
    wire N__69910;
    wire N__69907;
    wire N__69904;
    wire N__69903;
    wire N__69900;
    wire N__69897;
    wire N__69896;
    wire N__69893;
    wire N__69890;
    wire N__69889;
    wire N__69886;
    wire N__69883;
    wire N__69880;
    wire N__69879;
    wire N__69876;
    wire N__69873;
    wire N__69870;
    wire N__69867;
    wire N__69862;
    wire N__69853;
    wire N__69850;
    wire N__69849;
    wire N__69848;
    wire N__69845;
    wire N__69840;
    wire N__69835;
    wire N__69834;
    wire N__69831;
    wire N__69828;
    wire N__69827;
    wire N__69826;
    wire N__69825;
    wire N__69822;
    wire N__69819;
    wire N__69818;
    wire N__69817;
    wire N__69812;
    wire N__69809;
    wire N__69804;
    wire N__69801;
    wire N__69798;
    wire N__69787;
    wire N__69784;
    wire N__69781;
    wire N__69778;
    wire N__69777;
    wire N__69774;
    wire N__69773;
    wire N__69772;
    wire N__69769;
    wire N__69766;
    wire N__69761;
    wire N__69758;
    wire N__69753;
    wire N__69748;
    wire N__69747;
    wire N__69746;
    wire N__69745;
    wire N__69744;
    wire N__69739;
    wire N__69734;
    wire N__69731;
    wire N__69726;
    wire N__69723;
    wire N__69718;
    wire N__69715;
    wire N__69714;
    wire N__69711;
    wire N__69708;
    wire N__69707;
    wire N__69704;
    wire N__69701;
    wire N__69698;
    wire N__69695;
    wire N__69688;
    wire N__69685;
    wire N__69684;
    wire N__69683;
    wire N__69682;
    wire N__69679;
    wire N__69676;
    wire N__69673;
    wire N__69670;
    wire N__69661;
    wire N__69658;
    wire N__69657;
    wire N__69656;
    wire N__69653;
    wire N__69652;
    wire N__69649;
    wire N__69648;
    wire N__69645;
    wire N__69642;
    wire N__69637;
    wire N__69636;
    wire N__69633;
    wire N__69630;
    wire N__69625;
    wire N__69622;
    wire N__69619;
    wire N__69614;
    wire N__69607;
    wire N__69606;
    wire N__69603;
    wire N__69602;
    wire N__69599;
    wire N__69596;
    wire N__69595;
    wire N__69592;
    wire N__69589;
    wire N__69586;
    wire N__69583;
    wire N__69580;
    wire N__69577;
    wire N__69572;
    wire N__69565;
    wire N__69564;
    wire N__69561;
    wire N__69558;
    wire N__69557;
    wire N__69556;
    wire N__69555;
    wire N__69552;
    wire N__69547;
    wire N__69544;
    wire N__69543;
    wire N__69540;
    wire N__69537;
    wire N__69534;
    wire N__69529;
    wire N__69526;
    wire N__69517;
    wire N__69514;
    wire N__69511;
    wire N__69510;
    wire N__69509;
    wire N__69506;
    wire N__69501;
    wire N__69496;
    wire N__69493;
    wire N__69492;
    wire N__69489;
    wire N__69486;
    wire N__69483;
    wire N__69480;
    wire N__69475;
    wire N__69472;
    wire N__69469;
    wire N__69466;
    wire N__69465;
    wire N__69462;
    wire N__69459;
    wire N__69458;
    wire N__69455;
    wire N__69450;
    wire N__69445;
    wire N__69444;
    wire N__69443;
    wire N__69442;
    wire N__69439;
    wire N__69438;
    wire N__69437;
    wire N__69436;
    wire N__69435;
    wire N__69432;
    wire N__69429;
    wire N__69426;
    wire N__69425;
    wire N__69424;
    wire N__69423;
    wire N__69422;
    wire N__69421;
    wire N__69418;
    wire N__69415;
    wire N__69414;
    wire N__69411;
    wire N__69410;
    wire N__69409;
    wire N__69408;
    wire N__69405;
    wire N__69402;
    wire N__69399;
    wire N__69396;
    wire N__69393;
    wire N__69390;
    wire N__69385;
    wire N__69382;
    wire N__69381;
    wire N__69380;
    wire N__69377;
    wire N__69376;
    wire N__69371;
    wire N__69364;
    wire N__69363;
    wire N__69360;
    wire N__69357;
    wire N__69352;
    wire N__69349;
    wire N__69342;
    wire N__69339;
    wire N__69336;
    wire N__69331;
    wire N__69328;
    wire N__69325;
    wire N__69320;
    wire N__69317;
    wire N__69316;
    wire N__69315;
    wire N__69314;
    wire N__69311;
    wire N__69308;
    wire N__69301;
    wire N__69298;
    wire N__69293;
    wire N__69288;
    wire N__69287;
    wire N__69284;
    wire N__69279;
    wire N__69278;
    wire N__69277;
    wire N__69274;
    wire N__69271;
    wire N__69264;
    wire N__69261;
    wire N__69256;
    wire N__69253;
    wire N__69248;
    wire N__69247;
    wire N__69242;
    wire N__69239;
    wire N__69236;
    wire N__69233;
    wire N__69228;
    wire N__69225;
    wire N__69222;
    wire N__69219;
    wire N__69218;
    wire N__69217;
    wire N__69216;
    wire N__69215;
    wire N__69212;
    wire N__69207;
    wire N__69204;
    wire N__69201;
    wire N__69194;
    wire N__69189;
    wire N__69184;
    wire N__69169;
    wire N__69168;
    wire N__69167;
    wire N__69164;
    wire N__69161;
    wire N__69158;
    wire N__69155;
    wire N__69152;
    wire N__69151;
    wire N__69150;
    wire N__69147;
    wire N__69146;
    wire N__69143;
    wire N__69140;
    wire N__69139;
    wire N__69138;
    wire N__69133;
    wire N__69130;
    wire N__69127;
    wire N__69124;
    wire N__69121;
    wire N__69116;
    wire N__69111;
    wire N__69108;
    wire N__69105;
    wire N__69102;
    wire N__69097;
    wire N__69092;
    wire N__69089;
    wire N__69082;
    wire N__69081;
    wire N__69080;
    wire N__69079;
    wire N__69078;
    wire N__69071;
    wire N__69066;
    wire N__69063;
    wire N__69060;
    wire N__69057;
    wire N__69056;
    wire N__69055;
    wire N__69050;
    wire N__69045;
    wire N__69040;
    wire N__69037;
    wire N__69036;
    wire N__69035;
    wire N__69032;
    wire N__69031;
    wire N__69026;
    wire N__69025;
    wire N__69024;
    wire N__69023;
    wire N__69022;
    wire N__69019;
    wire N__69016;
    wire N__69015;
    wire N__69014;
    wire N__69013;
    wire N__69012;
    wire N__69011;
    wire N__69008;
    wire N__69007;
    wire N__69006;
    wire N__69003;
    wire N__69002;
    wire N__69001;
    wire N__68998;
    wire N__68995;
    wire N__68994;
    wire N__68991;
    wire N__68986;
    wire N__68981;
    wire N__68980;
    wire N__68977;
    wire N__68974;
    wire N__68973;
    wire N__68970;
    wire N__68967;
    wire N__68964;
    wire N__68961;
    wire N__68956;
    wire N__68953;
    wire N__68950;
    wire N__68945;
    wire N__68938;
    wire N__68935;
    wire N__68932;
    wire N__68929;
    wire N__68928;
    wire N__68927;
    wire N__68924;
    wire N__68923;
    wire N__68920;
    wire N__68917;
    wire N__68912;
    wire N__68909;
    wire N__68904;
    wire N__68903;
    wire N__68898;
    wire N__68895;
    wire N__68890;
    wire N__68887;
    wire N__68882;
    wire N__68879;
    wire N__68872;
    wire N__68867;
    wire N__68866;
    wire N__68863;
    wire N__68860;
    wire N__68855;
    wire N__68854;
    wire N__68853;
    wire N__68850;
    wire N__68845;
    wire N__68844;
    wire N__68843;
    wire N__68840;
    wire N__68837;
    wire N__68834;
    wire N__68827;
    wire N__68826;
    wire N__68825;
    wire N__68824;
    wire N__68821;
    wire N__68818;
    wire N__68813;
    wire N__68808;
    wire N__68803;
    wire N__68800;
    wire N__68797;
    wire N__68794;
    wire N__68789;
    wire N__68786;
    wire N__68781;
    wire N__68776;
    wire N__68771;
    wire N__68758;
    wire N__68755;
    wire N__68752;
    wire N__68751;
    wire N__68750;
    wire N__68747;
    wire N__68746;
    wire N__68745;
    wire N__68744;
    wire N__68741;
    wire N__68740;
    wire N__68737;
    wire N__68734;
    wire N__68731;
    wire N__68728;
    wire N__68727;
    wire N__68726;
    wire N__68725;
    wire N__68724;
    wire N__68723;
    wire N__68722;
    wire N__68719;
    wire N__68716;
    wire N__68713;
    wire N__68712;
    wire N__68711;
    wire N__68708;
    wire N__68701;
    wire N__68698;
    wire N__68695;
    wire N__68692;
    wire N__68691;
    wire N__68688;
    wire N__68683;
    wire N__68682;
    wire N__68675;
    wire N__68674;
    wire N__68671;
    wire N__68668;
    wire N__68657;
    wire N__68656;
    wire N__68655;
    wire N__68652;
    wire N__68649;
    wire N__68648;
    wire N__68647;
    wire N__68646;
    wire N__68645;
    wire N__68644;
    wire N__68641;
    wire N__68638;
    wire N__68635;
    wire N__68632;
    wire N__68629;
    wire N__68626;
    wire N__68623;
    wire N__68622;
    wire N__68619;
    wire N__68616;
    wire N__68613;
    wire N__68612;
    wire N__68609;
    wire N__68604;
    wire N__68601;
    wire N__68598;
    wire N__68595;
    wire N__68594;
    wire N__68593;
    wire N__68590;
    wire N__68587;
    wire N__68584;
    wire N__68581;
    wire N__68576;
    wire N__68573;
    wire N__68570;
    wire N__68565;
    wire N__68562;
    wire N__68559;
    wire N__68554;
    wire N__68553;
    wire N__68546;
    wire N__68543;
    wire N__68540;
    wire N__68535;
    wire N__68532;
    wire N__68529;
    wire N__68526;
    wire N__68523;
    wire N__68522;
    wire N__68521;
    wire N__68518;
    wire N__68515;
    wire N__68512;
    wire N__68509;
    wire N__68506;
    wire N__68503;
    wire N__68500;
    wire N__68495;
    wire N__68492;
    wire N__68489;
    wire N__68484;
    wire N__68481;
    wire N__68476;
    wire N__68473;
    wire N__68470;
    wire N__68463;
    wire N__68456;
    wire N__68447;
    wire N__68434;
    wire N__68431;
    wire N__68430;
    wire N__68429;
    wire N__68428;
    wire N__68425;
    wire N__68422;
    wire N__68419;
    wire N__68416;
    wire N__68413;
    wire N__68410;
    wire N__68405;
    wire N__68398;
    wire N__68395;
    wire N__68392;
    wire N__68391;
    wire N__68388;
    wire N__68385;
    wire N__68384;
    wire N__68383;
    wire N__68378;
    wire N__68375;
    wire N__68374;
    wire N__68371;
    wire N__68368;
    wire N__68365;
    wire N__68364;
    wire N__68361;
    wire N__68356;
    wire N__68355;
    wire N__68352;
    wire N__68349;
    wire N__68348;
    wire N__68345;
    wire N__68342;
    wire N__68339;
    wire N__68336;
    wire N__68333;
    wire N__68330;
    wire N__68327;
    wire N__68324;
    wire N__68317;
    wire N__68308;
    wire N__68307;
    wire N__68304;
    wire N__68301;
    wire N__68300;
    wire N__68299;
    wire N__68296;
    wire N__68293;
    wire N__68290;
    wire N__68289;
    wire N__68286;
    wire N__68283;
    wire N__68278;
    wire N__68275;
    wire N__68274;
    wire N__68271;
    wire N__68266;
    wire N__68263;
    wire N__68260;
    wire N__68257;
    wire N__68252;
    wire N__68245;
    wire N__68242;
    wire N__68239;
    wire N__68236;
    wire N__68235;
    wire N__68234;
    wire N__68229;
    wire N__68228;
    wire N__68227;
    wire N__68224;
    wire N__68221;
    wire N__68218;
    wire N__68217;
    wire N__68214;
    wire N__68213;
    wire N__68208;
    wire N__68203;
    wire N__68200;
    wire N__68197;
    wire N__68196;
    wire N__68195;
    wire N__68192;
    wire N__68185;
    wire N__68180;
    wire N__68173;
    wire N__68170;
    wire N__68169;
    wire N__68166;
    wire N__68165;
    wire N__68162;
    wire N__68159;
    wire N__68158;
    wire N__68157;
    wire N__68154;
    wire N__68151;
    wire N__68148;
    wire N__68143;
    wire N__68140;
    wire N__68133;
    wire N__68130;
    wire N__68125;
    wire N__68124;
    wire N__68121;
    wire N__68120;
    wire N__68119;
    wire N__68114;
    wire N__68113;
    wire N__68112;
    wire N__68109;
    wire N__68106;
    wire N__68105;
    wire N__68104;
    wire N__68101;
    wire N__68096;
    wire N__68093;
    wire N__68090;
    wire N__68085;
    wire N__68084;
    wire N__68081;
    wire N__68076;
    wire N__68071;
    wire N__68070;
    wire N__68067;
    wire N__68064;
    wire N__68059;
    wire N__68056;
    wire N__68047;
    wire N__68044;
    wire N__68043;
    wire N__68040;
    wire N__68037;
    wire N__68034;
    wire N__68031;
    wire N__68026;
    wire N__68023;
    wire N__68022;
    wire N__68019;
    wire N__68018;
    wire N__68017;
    wire N__68014;
    wire N__68011;
    wire N__68008;
    wire N__68005;
    wire N__68002;
    wire N__67993;
    wire N__67990;
    wire N__67987;
    wire N__67984;
    wire N__67983;
    wire N__67982;
    wire N__67981;
    wire N__67980;
    wire N__67979;
    wire N__67976;
    wire N__67973;
    wire N__67972;
    wire N__67971;
    wire N__67968;
    wire N__67965;
    wire N__67964;
    wire N__67961;
    wire N__67958;
    wire N__67953;
    wire N__67952;
    wire N__67951;
    wire N__67950;
    wire N__67949;
    wire N__67948;
    wire N__67947;
    wire N__67946;
    wire N__67945;
    wire N__67944;
    wire N__67941;
    wire N__67940;
    wire N__67939;
    wire N__67936;
    wire N__67933;
    wire N__67932;
    wire N__67929;
    wire N__67926;
    wire N__67923;
    wire N__67922;
    wire N__67921;
    wire N__67920;
    wire N__67919;
    wire N__67916;
    wire N__67913;
    wire N__67912;
    wire N__67911;
    wire N__67908;
    wire N__67905;
    wire N__67900;
    wire N__67897;
    wire N__67890;
    wire N__67889;
    wire N__67886;
    wire N__67883;
    wire N__67880;
    wire N__67877;
    wire N__67872;
    wire N__67869;
    wire N__67866;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67854;
    wire N__67849;
    wire N__67846;
    wire N__67843;
    wire N__67840;
    wire N__67837;
    wire N__67826;
    wire N__67821;
    wire N__67818;
    wire N__67813;
    wire N__67808;
    wire N__67803;
    wire N__67802;
    wire N__67799;
    wire N__67796;
    wire N__67793;
    wire N__67790;
    wire N__67785;
    wire N__67778;
    wire N__67777;
    wire N__67776;
    wire N__67773;
    wire N__67770;
    wire N__67763;
    wire N__67760;
    wire N__67757;
    wire N__67750;
    wire N__67747;
    wire N__67744;
    wire N__67741;
    wire N__67738;
    wire N__67733;
    wire N__67730;
    wire N__67723;
    wire N__67718;
    wire N__67705;
    wire N__67704;
    wire N__67701;
    wire N__67698;
    wire N__67697;
    wire N__67696;
    wire N__67693;
    wire N__67690;
    wire N__67685;
    wire N__67682;
    wire N__67675;
    wire N__67674;
    wire N__67673;
    wire N__67670;
    wire N__67667;
    wire N__67666;
    wire N__67663;
    wire N__67658;
    wire N__67657;
    wire N__67654;
    wire N__67649;
    wire N__67646;
    wire N__67639;
    wire N__67636;
    wire N__67633;
    wire N__67630;
    wire N__67629;
    wire N__67626;
    wire N__67623;
    wire N__67618;
    wire N__67615;
    wire N__67614;
    wire N__67613;
    wire N__67610;
    wire N__67607;
    wire N__67604;
    wire N__67601;
    wire N__67598;
    wire N__67595;
    wire N__67590;
    wire N__67587;
    wire N__67582;
    wire N__67579;
    wire N__67576;
    wire N__67573;
    wire N__67570;
    wire N__67567;
    wire N__67566;
    wire N__67563;
    wire N__67562;
    wire N__67559;
    wire N__67556;
    wire N__67553;
    wire N__67550;
    wire N__67547;
    wire N__67544;
    wire N__67541;
    wire N__67538;
    wire N__67531;
    wire N__67530;
    wire N__67529;
    wire N__67528;
    wire N__67527;
    wire N__67526;
    wire N__67523;
    wire N__67522;
    wire N__67519;
    wire N__67516;
    wire N__67511;
    wire N__67508;
    wire N__67505;
    wire N__67504;
    wire N__67501;
    wire N__67498;
    wire N__67495;
    wire N__67492;
    wire N__67489;
    wire N__67486;
    wire N__67483;
    wire N__67478;
    wire N__67475;
    wire N__67472;
    wire N__67467;
    wire N__67462;
    wire N__67459;
    wire N__67456;
    wire N__67453;
    wire N__67450;
    wire N__67447;
    wire N__67438;
    wire N__67435;
    wire N__67434;
    wire N__67431;
    wire N__67428;
    wire N__67427;
    wire N__67424;
    wire N__67421;
    wire N__67418;
    wire N__67413;
    wire N__67408;
    wire N__67405;
    wire N__67404;
    wire N__67401;
    wire N__67398;
    wire N__67393;
    wire N__67390;
    wire N__67387;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67379;
    wire N__67378;
    wire N__67373;
    wire N__67368;
    wire N__67365;
    wire N__67360;
    wire N__67357;
    wire N__67354;
    wire N__67351;
    wire N__67348;
    wire N__67345;
    wire N__67342;
    wire N__67339;
    wire N__67336;
    wire N__67333;
    wire N__67330;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67318;
    wire N__67315;
    wire N__67312;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67302;
    wire N__67299;
    wire N__67296;
    wire N__67293;
    wire N__67290;
    wire N__67289;
    wire N__67288;
    wire N__67285;
    wire N__67282;
    wire N__67277;
    wire N__67270;
    wire N__67267;
    wire N__67266;
    wire N__67265;
    wire N__67264;
    wire N__67263;
    wire N__67260;
    wire N__67255;
    wire N__67250;
    wire N__67243;
    wire N__67242;
    wire N__67241;
    wire N__67234;
    wire N__67231;
    wire N__67228;
    wire N__67227;
    wire N__67226;
    wire N__67225;
    wire N__67224;
    wire N__67223;
    wire N__67222;
    wire N__67221;
    wire N__67220;
    wire N__67219;
    wire N__67218;
    wire N__67213;
    wire N__67204;
    wire N__67201;
    wire N__67200;
    wire N__67199;
    wire N__67198;
    wire N__67197;
    wire N__67196;
    wire N__67191;
    wire N__67188;
    wire N__67187;
    wire N__67184;
    wire N__67179;
    wire N__67178;
    wire N__67173;
    wire N__67170;
    wire N__67167;
    wire N__67166;
    wire N__67163;
    wire N__67160;
    wire N__67157;
    wire N__67154;
    wire N__67151;
    wire N__67148;
    wire N__67145;
    wire N__67144;
    wire N__67141;
    wire N__67138;
    wire N__67135;
    wire N__67132;
    wire N__67131;
    wire N__67130;
    wire N__67127;
    wire N__67122;
    wire N__67119;
    wire N__67118;
    wire N__67113;
    wire N__67108;
    wire N__67105;
    wire N__67102;
    wire N__67095;
    wire N__67092;
    wire N__67089;
    wire N__67086;
    wire N__67081;
    wire N__67078;
    wire N__67075;
    wire N__67072;
    wire N__67065;
    wire N__67062;
    wire N__67057;
    wire N__67054;
    wire N__67051;
    wire N__67044;
    wire N__67041;
    wire N__67038;
    wire N__67035;
    wire N__67030;
    wire N__67021;
    wire N__67020;
    wire N__67017;
    wire N__67014;
    wire N__67011;
    wire N__67008;
    wire N__67005;
    wire N__67002;
    wire N__66999;
    wire N__66994;
    wire N__66991;
    wire N__66988;
    wire N__66987;
    wire N__66984;
    wire N__66981;
    wire N__66980;
    wire N__66979;
    wire N__66978;
    wire N__66977;
    wire N__66976;
    wire N__66975;
    wire N__66974;
    wire N__66973;
    wire N__66972;
    wire N__66963;
    wire N__66962;
    wire N__66959;
    wire N__66958;
    wire N__66957;
    wire N__66956;
    wire N__66955;
    wire N__66954;
    wire N__66953;
    wire N__66952;
    wire N__66949;
    wire N__66948;
    wire N__66947;
    wire N__66944;
    wire N__66943;
    wire N__66942;
    wire N__66941;
    wire N__66938;
    wire N__66935;
    wire N__66934;
    wire N__66933;
    wire N__66928;
    wire N__66925;
    wire N__66924;
    wire N__66923;
    wire N__66918;
    wire N__66917;
    wire N__66916;
    wire N__66913;
    wire N__66912;
    wire N__66909;
    wire N__66900;
    wire N__66899;
    wire N__66898;
    wire N__66897;
    wire N__66896;
    wire N__66889;
    wire N__66882;
    wire N__66881;
    wire N__66880;
    wire N__66879;
    wire N__66868;
    wire N__66865;
    wire N__66860;
    wire N__66857;
    wire N__66854;
    wire N__66851;
    wire N__66850;
    wire N__66849;
    wire N__66846;
    wire N__66841;
    wire N__66838;
    wire N__66835;
    wire N__66832;
    wire N__66829;
    wire N__66826;
    wire N__66821;
    wire N__66816;
    wire N__66809;
    wire N__66806;
    wire N__66799;
    wire N__66794;
    wire N__66791;
    wire N__66788;
    wire N__66785;
    wire N__66782;
    wire N__66777;
    wire N__66774;
    wire N__66771;
    wire N__66768;
    wire N__66761;
    wire N__66758;
    wire N__66755;
    wire N__66754;
    wire N__66751;
    wire N__66748;
    wire N__66739;
    wire N__66732;
    wire N__66729;
    wire N__66724;
    wire N__66721;
    wire N__66718;
    wire N__66711;
    wire N__66708;
    wire N__66705;
    wire N__66694;
    wire N__66691;
    wire N__66690;
    wire N__66687;
    wire N__66684;
    wire N__66681;
    wire N__66676;
    wire N__66673;
    wire N__66670;
    wire N__66667;
    wire N__66664;
    wire N__66661;
    wire N__66658;
    wire N__66655;
    wire N__66652;
    wire N__66649;
    wire N__66648;
    wire N__66647;
    wire N__66644;
    wire N__66641;
    wire N__66636;
    wire N__66633;
    wire N__66632;
    wire N__66631;
    wire N__66628;
    wire N__66625;
    wire N__66622;
    wire N__66619;
    wire N__66616;
    wire N__66613;
    wire N__66604;
    wire N__66601;
    wire N__66598;
    wire N__66595;
    wire N__66592;
    wire N__66589;
    wire N__66586;
    wire N__66583;
    wire N__66582;
    wire N__66579;
    wire N__66576;
    wire N__66571;
    wire N__66570;
    wire N__66567;
    wire N__66564;
    wire N__66559;
    wire N__66556;
    wire N__66553;
    wire N__66550;
    wire N__66547;
    wire N__66546;
    wire N__66545;
    wire N__66542;
    wire N__66537;
    wire N__66532;
    wire N__66529;
    wire N__66526;
    wire N__66523;
    wire N__66520;
    wire N__66517;
    wire N__66514;
    wire N__66511;
    wire N__66510;
    wire N__66507;
    wire N__66504;
    wire N__66501;
    wire N__66500;
    wire N__66497;
    wire N__66496;
    wire N__66493;
    wire N__66490;
    wire N__66487;
    wire N__66484;
    wire N__66481;
    wire N__66476;
    wire N__66469;
    wire N__66466;
    wire N__66465;
    wire N__66464;
    wire N__66461;
    wire N__66458;
    wire N__66455;
    wire N__66454;
    wire N__66453;
    wire N__66448;
    wire N__66445;
    wire N__66440;
    wire N__66437;
    wire N__66434;
    wire N__66427;
    wire N__66424;
    wire N__66421;
    wire N__66418;
    wire N__66417;
    wire N__66416;
    wire N__66411;
    wire N__66408;
    wire N__66405;
    wire N__66402;
    wire N__66397;
    wire N__66396;
    wire N__66395;
    wire N__66392;
    wire N__66387;
    wire N__66382;
    wire N__66381;
    wire N__66378;
    wire N__66375;
    wire N__66370;
    wire N__66367;
    wire N__66364;
    wire N__66361;
    wire N__66358;
    wire N__66355;
    wire N__66354;
    wire N__66351;
    wire N__66348;
    wire N__66345;
    wire N__66342;
    wire N__66337;
    wire N__66336;
    wire N__66333;
    wire N__66330;
    wire N__66327;
    wire N__66326;
    wire N__66323;
    wire N__66320;
    wire N__66317;
    wire N__66310;
    wire N__66307;
    wire N__66304;
    wire N__66301;
    wire N__66298;
    wire N__66295;
    wire N__66294;
    wire N__66291;
    wire N__66288;
    wire N__66287;
    wire N__66286;
    wire N__66281;
    wire N__66278;
    wire N__66275;
    wire N__66272;
    wire N__66269;
    wire N__66266;
    wire N__66261;
    wire N__66256;
    wire N__66253;
    wire N__66250;
    wire N__66247;
    wire N__66244;
    wire N__66243;
    wire N__66240;
    wire N__66239;
    wire N__66236;
    wire N__66233;
    wire N__66230;
    wire N__66227;
    wire N__66224;
    wire N__66221;
    wire N__66216;
    wire N__66211;
    wire N__66210;
    wire N__66209;
    wire N__66206;
    wire N__66205;
    wire N__66204;
    wire N__66203;
    wire N__66198;
    wire N__66195;
    wire N__66194;
    wire N__66193;
    wire N__66190;
    wire N__66189;
    wire N__66188;
    wire N__66187;
    wire N__66186;
    wire N__66185;
    wire N__66184;
    wire N__66181;
    wire N__66178;
    wire N__66177;
    wire N__66172;
    wire N__66169;
    wire N__66166;
    wire N__66163;
    wire N__66162;
    wire N__66159;
    wire N__66158;
    wire N__66157;
    wire N__66156;
    wire N__66155;
    wire N__66154;
    wire N__66153;
    wire N__66150;
    wire N__66147;
    wire N__66146;
    wire N__66145;
    wire N__66144;
    wire N__66141;
    wire N__66140;
    wire N__66139;
    wire N__66136;
    wire N__66133;
    wire N__66126;
    wire N__66125;
    wire N__66122;
    wire N__66121;
    wire N__66120;
    wire N__66117;
    wire N__66114;
    wire N__66111;
    wire N__66102;
    wire N__66099;
    wire N__66096;
    wire N__66093;
    wire N__66084;
    wire N__66081;
    wire N__66078;
    wire N__66071;
    wire N__66068;
    wire N__66067;
    wire N__66066;
    wire N__66061;
    wire N__66060;
    wire N__66057;
    wire N__66054;
    wire N__66051;
    wire N__66050;
    wire N__66047;
    wire N__66046;
    wire N__66045;
    wire N__66040;
    wire N__66039;
    wire N__66038;
    wire N__66033;
    wire N__66026;
    wire N__66023;
    wire N__66020;
    wire N__66013;
    wire N__66012;
    wire N__66011;
    wire N__66008;
    wire N__66007;
    wire N__66004;
    wire N__66001;
    wire N__65998;
    wire N__65995;
    wire N__65992;
    wire N__65989;
    wire N__65986;
    wire N__65979;
    wire N__65976;
    wire N__65971;
    wire N__65968;
    wire N__65965;
    wire N__65958;
    wire N__65955;
    wire N__65952;
    wire N__65949;
    wire N__65944;
    wire N__65941;
    wire N__65936;
    wire N__65933;
    wire N__65930;
    wire N__65921;
    wire N__65918;
    wire N__65913;
    wire N__65904;
    wire N__65901;
    wire N__65894;
    wire N__65891;
    wire N__65888;
    wire N__65885;
    wire N__65878;
    wire N__65869;
    wire N__65868;
    wire N__65865;
    wire N__65864;
    wire N__65863;
    wire N__65860;
    wire N__65857;
    wire N__65854;
    wire N__65853;
    wire N__65850;
    wire N__65849;
    wire N__65846;
    wire N__65843;
    wire N__65840;
    wire N__65837;
    wire N__65834;
    wire N__65831;
    wire N__65828;
    wire N__65823;
    wire N__65818;
    wire N__65815;
    wire N__65812;
    wire N__65809;
    wire N__65806;
    wire N__65797;
    wire N__65796;
    wire N__65795;
    wire N__65792;
    wire N__65789;
    wire N__65786;
    wire N__65783;
    wire N__65782;
    wire N__65781;
    wire N__65780;
    wire N__65775;
    wire N__65772;
    wire N__65769;
    wire N__65766;
    wire N__65763;
    wire N__65762;
    wire N__65759;
    wire N__65752;
    wire N__65749;
    wire N__65746;
    wire N__65743;
    wire N__65738;
    wire N__65735;
    wire N__65732;
    wire N__65729;
    wire N__65722;
    wire N__65719;
    wire N__65716;
    wire N__65715;
    wire N__65712;
    wire N__65711;
    wire N__65708;
    wire N__65705;
    wire N__65702;
    wire N__65695;
    wire N__65694;
    wire N__65693;
    wire N__65690;
    wire N__65687;
    wire N__65684;
    wire N__65681;
    wire N__65680;
    wire N__65675;
    wire N__65674;
    wire N__65671;
    wire N__65668;
    wire N__65665;
    wire N__65662;
    wire N__65661;
    wire N__65658;
    wire N__65655;
    wire N__65652;
    wire N__65649;
    wire N__65646;
    wire N__65643;
    wire N__65638;
    wire N__65635;
    wire N__65626;
    wire N__65623;
    wire N__65620;
    wire N__65619;
    wire N__65618;
    wire N__65615;
    wire N__65610;
    wire N__65605;
    wire N__65602;
    wire N__65599;
    wire N__65598;
    wire N__65597;
    wire N__65596;
    wire N__65595;
    wire N__65594;
    wire N__65591;
    wire N__65590;
    wire N__65587;
    wire N__65584;
    wire N__65581;
    wire N__65580;
    wire N__65575;
    wire N__65572;
    wire N__65569;
    wire N__65566;
    wire N__65563;
    wire N__65560;
    wire N__65557;
    wire N__65554;
    wire N__65551;
    wire N__65544;
    wire N__65541;
    wire N__65532;
    wire N__65527;
    wire N__65526;
    wire N__65525;
    wire N__65522;
    wire N__65521;
    wire N__65520;
    wire N__65519;
    wire N__65516;
    wire N__65515;
    wire N__65512;
    wire N__65509;
    wire N__65504;
    wire N__65499;
    wire N__65496;
    wire N__65495;
    wire N__65494;
    wire N__65493;
    wire N__65490;
    wire N__65485;
    wire N__65482;
    wire N__65479;
    wire N__65474;
    wire N__65471;
    wire N__65466;
    wire N__65459;
    wire N__65452;
    wire N__65449;
    wire N__65448;
    wire N__65445;
    wire N__65442;
    wire N__65439;
    wire N__65434;
    wire N__65433;
    wire N__65430;
    wire N__65429;
    wire N__65426;
    wire N__65423;
    wire N__65420;
    wire N__65417;
    wire N__65412;
    wire N__65407;
    wire N__65406;
    wire N__65403;
    wire N__65400;
    wire N__65399;
    wire N__65398;
    wire N__65397;
    wire N__65394;
    wire N__65391;
    wire N__65388;
    wire N__65385;
    wire N__65382;
    wire N__65379;
    wire N__65374;
    wire N__65371;
    wire N__65368;
    wire N__65365;
    wire N__65362;
    wire N__65359;
    wire N__65350;
    wire N__65347;
    wire N__65344;
    wire N__65343;
    wire N__65340;
    wire N__65337;
    wire N__65334;
    wire N__65331;
    wire N__65326;
    wire N__65325;
    wire N__65322;
    wire N__65321;
    wire N__65320;
    wire N__65317;
    wire N__65314;
    wire N__65309;
    wire N__65306;
    wire N__65299;
    wire N__65298;
    wire N__65293;
    wire N__65292;
    wire N__65289;
    wire N__65286;
    wire N__65281;
    wire N__65278;
    wire N__65275;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65263;
    wire N__65262;
    wire N__65261;
    wire N__65260;
    wire N__65259;
    wire N__65258;
    wire N__65253;
    wire N__65250;
    wire N__65249;
    wire N__65248;
    wire N__65247;
    wire N__65246;
    wire N__65243;
    wire N__65242;
    wire N__65241;
    wire N__65240;
    wire N__65239;
    wire N__65238;
    wire N__65235;
    wire N__65234;
    wire N__65231;
    wire N__65230;
    wire N__65227;
    wire N__65226;
    wire N__65223;
    wire N__65218;
    wire N__65217;
    wire N__65212;
    wire N__65209;
    wire N__65206;
    wire N__65203;
    wire N__65202;
    wire N__65199;
    wire N__65198;
    wire N__65195;
    wire N__65192;
    wire N__65191;
    wire N__65190;
    wire N__65189;
    wire N__65186;
    wire N__65179;
    wire N__65176;
    wire N__65173;
    wire N__65172;
    wire N__65169;
    wire N__65166;
    wire N__65163;
    wire N__65160;
    wire N__65155;
    wire N__65152;
    wire N__65149;
    wire N__65148;
    wire N__65147;
    wire N__65144;
    wire N__65141;
    wire N__65136;
    wire N__65129;
    wire N__65124;
    wire N__65119;
    wire N__65118;
    wire N__65117;
    wire N__65114;
    wire N__65109;
    wire N__65104;
    wire N__65101;
    wire N__65098;
    wire N__65095;
    wire N__65094;
    wire N__65091;
    wire N__65088;
    wire N__65085;
    wire N__65082;
    wire N__65079;
    wire N__65074;
    wire N__65071;
    wire N__65070;
    wire N__65069;
    wire N__65064;
    wire N__65057;
    wire N__65052;
    wire N__65049;
    wire N__65046;
    wire N__65037;
    wire N__65034;
    wire N__65031;
    wire N__65028;
    wire N__65025;
    wire N__65022;
    wire N__65019;
    wire N__65014;
    wire N__65011;
    wire N__65000;
    wire N__64991;
    wire N__64984;
    wire N__64983;
    wire N__64980;
    wire N__64979;
    wire N__64976;
    wire N__64973;
    wire N__64972;
    wire N__64969;
    wire N__64966;
    wire N__64963;
    wire N__64960;
    wire N__64951;
    wire N__64950;
    wire N__64949;
    wire N__64946;
    wire N__64943;
    wire N__64942;
    wire N__64939;
    wire N__64936;
    wire N__64933;
    wire N__64930;
    wire N__64927;
    wire N__64924;
    wire N__64921;
    wire N__64920;
    wire N__64917;
    wire N__64910;
    wire N__64907;
    wire N__64900;
    wire N__64899;
    wire N__64896;
    wire N__64893;
    wire N__64892;
    wire N__64889;
    wire N__64888;
    wire N__64887;
    wire N__64886;
    wire N__64883;
    wire N__64880;
    wire N__64877;
    wire N__64874;
    wire N__64871;
    wire N__64868;
    wire N__64865;
    wire N__64860;
    wire N__64857;
    wire N__64854;
    wire N__64849;
    wire N__64846;
    wire N__64843;
    wire N__64834;
    wire N__64833;
    wire N__64832;
    wire N__64831;
    wire N__64830;
    wire N__64827;
    wire N__64822;
    wire N__64821;
    wire N__64818;
    wire N__64815;
    wire N__64812;
    wire N__64809;
    wire N__64806;
    wire N__64803;
    wire N__64800;
    wire N__64795;
    wire N__64792;
    wire N__64789;
    wire N__64786;
    wire N__64781;
    wire N__64776;
    wire N__64771;
    wire N__64770;
    wire N__64769;
    wire N__64764;
    wire N__64761;
    wire N__64760;
    wire N__64757;
    wire N__64754;
    wire N__64751;
    wire N__64748;
    wire N__64745;
    wire N__64742;
    wire N__64739;
    wire N__64736;
    wire N__64731;
    wire N__64728;
    wire N__64723;
    wire N__64720;
    wire N__64717;
    wire N__64714;
    wire N__64711;
    wire N__64708;
    wire N__64707;
    wire N__64704;
    wire N__64703;
    wire N__64700;
    wire N__64699;
    wire N__64696;
    wire N__64693;
    wire N__64690;
    wire N__64687;
    wire N__64684;
    wire N__64683;
    wire N__64680;
    wire N__64675;
    wire N__64672;
    wire N__64669;
    wire N__64666;
    wire N__64661;
    wire N__64658;
    wire N__64655;
    wire N__64652;
    wire N__64645;
    wire N__64642;
    wire N__64639;
    wire N__64636;
    wire N__64633;
    wire N__64632;
    wire N__64629;
    wire N__64628;
    wire N__64625;
    wire N__64624;
    wire N__64623;
    wire N__64620;
    wire N__64617;
    wire N__64614;
    wire N__64609;
    wire N__64608;
    wire N__64603;
    wire N__64598;
    wire N__64595;
    wire N__64590;
    wire N__64585;
    wire N__64584;
    wire N__64583;
    wire N__64582;
    wire N__64579;
    wire N__64578;
    wire N__64577;
    wire N__64574;
    wire N__64569;
    wire N__64566;
    wire N__64565;
    wire N__64564;
    wire N__64561;
    wire N__64558;
    wire N__64555;
    wire N__64552;
    wire N__64551;
    wire N__64550;
    wire N__64549;
    wire N__64548;
    wire N__64547;
    wire N__64546;
    wire N__64543;
    wire N__64542;
    wire N__64535;
    wire N__64530;
    wire N__64527;
    wire N__64524;
    wire N__64519;
    wire N__64512;
    wire N__64509;
    wire N__64506;
    wire N__64503;
    wire N__64502;
    wire N__64499;
    wire N__64496;
    wire N__64493;
    wire N__64486;
    wire N__64481;
    wire N__64478;
    wire N__64475;
    wire N__64472;
    wire N__64467;
    wire N__64464;
    wire N__64453;
    wire N__64450;
    wire N__64449;
    wire N__64446;
    wire N__64443;
    wire N__64442;
    wire N__64439;
    wire N__64438;
    wire N__64435;
    wire N__64432;
    wire N__64429;
    wire N__64426;
    wire N__64423;
    wire N__64414;
    wire N__64413;
    wire N__64412;
    wire N__64411;
    wire N__64410;
    wire N__64409;
    wire N__64406;
    wire N__64401;
    wire N__64398;
    wire N__64397;
    wire N__64394;
    wire N__64393;
    wire N__64390;
    wire N__64389;
    wire N__64388;
    wire N__64387;
    wire N__64386;
    wire N__64379;
    wire N__64376;
    wire N__64373;
    wire N__64370;
    wire N__64367;
    wire N__64366;
    wire N__64363;
    wire N__64362;
    wire N__64355;
    wire N__64352;
    wire N__64349;
    wire N__64346;
    wire N__64345;
    wire N__64344;
    wire N__64341;
    wire N__64340;
    wire N__64337;
    wire N__64330;
    wire N__64327;
    wire N__64322;
    wire N__64319;
    wire N__64314;
    wire N__64311;
    wire N__64308;
    wire N__64305;
    wire N__64302;
    wire N__64299;
    wire N__64296;
    wire N__64293;
    wire N__64290;
    wire N__64287;
    wire N__64284;
    wire N__64279;
    wire N__64272;
    wire N__64267;
    wire N__64264;
    wire N__64255;
    wire N__64254;
    wire N__64253;
    wire N__64252;
    wire N__64251;
    wire N__64250;
    wire N__64249;
    wire N__64248;
    wire N__64247;
    wire N__64246;
    wire N__64245;
    wire N__64244;
    wire N__64243;
    wire N__64242;
    wire N__64239;
    wire N__64238;
    wire N__64237;
    wire N__64228;
    wire N__64225;
    wire N__64222;
    wire N__64221;
    wire N__64220;
    wire N__64217;
    wire N__64210;
    wire N__64203;
    wire N__64200;
    wire N__64199;
    wire N__64198;
    wire N__64193;
    wire N__64188;
    wire N__64185;
    wire N__64184;
    wire N__64183;
    wire N__64180;
    wire N__64177;
    wire N__64174;
    wire N__64167;
    wire N__64164;
    wire N__64161;
    wire N__64158;
    wire N__64153;
    wire N__64148;
    wire N__64145;
    wire N__64140;
    wire N__64137;
    wire N__64136;
    wire N__64133;
    wire N__64130;
    wire N__64127;
    wire N__64124;
    wire N__64121;
    wire N__64114;
    wire N__64113;
    wire N__64110;
    wire N__64107;
    wire N__64104;
    wire N__64101;
    wire N__64096;
    wire N__64093;
    wire N__64090;
    wire N__64087;
    wire N__64084;
    wire N__64081;
    wire N__64078;
    wire N__64075;
    wire N__64072;
    wire N__64057;
    wire N__64056;
    wire N__64053;
    wire N__64050;
    wire N__64049;
    wire N__64046;
    wire N__64043;
    wire N__64040;
    wire N__64039;
    wire N__64036;
    wire N__64033;
    wire N__64028;
    wire N__64021;
    wire N__64018;
    wire N__64015;
    wire N__64014;
    wire N__64013;
    wire N__64010;
    wire N__64007;
    wire N__64004;
    wire N__64003;
    wire N__64002;
    wire N__63999;
    wire N__63996;
    wire N__63995;
    wire N__63994;
    wire N__63991;
    wire N__63988;
    wire N__63985;
    wire N__63982;
    wire N__63979;
    wire N__63974;
    wire N__63971;
    wire N__63968;
    wire N__63955;
    wire N__63952;
    wire N__63949;
    wire N__63948;
    wire N__63945;
    wire N__63944;
    wire N__63943;
    wire N__63940;
    wire N__63939;
    wire N__63938;
    wire N__63937;
    wire N__63934;
    wire N__63931;
    wire N__63928;
    wire N__63925;
    wire N__63922;
    wire N__63919;
    wire N__63916;
    wire N__63915;
    wire N__63910;
    wire N__63907;
    wire N__63900;
    wire N__63897;
    wire N__63894;
    wire N__63891;
    wire N__63888;
    wire N__63885;
    wire N__63880;
    wire N__63871;
    wire N__63870;
    wire N__63865;
    wire N__63862;
    wire N__63861;
    wire N__63858;
    wire N__63855;
    wire N__63854;
    wire N__63853;
    wire N__63850;
    wire N__63847;
    wire N__63844;
    wire N__63843;
    wire N__63840;
    wire N__63837;
    wire N__63834;
    wire N__63831;
    wire N__63828;
    wire N__63825;
    wire N__63822;
    wire N__63819;
    wire N__63814;
    wire N__63805;
    wire N__63802;
    wire N__63799;
    wire N__63796;
    wire N__63795;
    wire N__63794;
    wire N__63791;
    wire N__63786;
    wire N__63781;
    wire N__63778;
    wire N__63777;
    wire N__63776;
    wire N__63775;
    wire N__63774;
    wire N__63771;
    wire N__63768;
    wire N__63767;
    wire N__63766;
    wire N__63765;
    wire N__63762;
    wire N__63759;
    wire N__63756;
    wire N__63753;
    wire N__63748;
    wire N__63743;
    wire N__63742;
    wire N__63741;
    wire N__63736;
    wire N__63733;
    wire N__63728;
    wire N__63725;
    wire N__63720;
    wire N__63715;
    wire N__63712;
    wire N__63709;
    wire N__63700;
    wire N__63697;
    wire N__63694;
    wire N__63691;
    wire N__63688;
    wire N__63687;
    wire N__63684;
    wire N__63683;
    wire N__63680;
    wire N__63679;
    wire N__63678;
    wire N__63673;
    wire N__63670;
    wire N__63665;
    wire N__63658;
    wire N__63655;
    wire N__63652;
    wire N__63651;
    wire N__63648;
    wire N__63647;
    wire N__63646;
    wire N__63643;
    wire N__63640;
    wire N__63637;
    wire N__63634;
    wire N__63631;
    wire N__63630;
    wire N__63629;
    wire N__63628;
    wire N__63627;
    wire N__63622;
    wire N__63619;
    wire N__63616;
    wire N__63611;
    wire N__63608;
    wire N__63605;
    wire N__63602;
    wire N__63597;
    wire N__63590;
    wire N__63583;
    wire N__63580;
    wire N__63577;
    wire N__63576;
    wire N__63575;
    wire N__63574;
    wire N__63573;
    wire N__63570;
    wire N__63567;
    wire N__63564;
    wire N__63561;
    wire N__63560;
    wire N__63557;
    wire N__63552;
    wire N__63549;
    wire N__63546;
    wire N__63543;
    wire N__63540;
    wire N__63535;
    wire N__63534;
    wire N__63529;
    wire N__63526;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63512;
    wire N__63509;
    wire N__63506;
    wire N__63503;
    wire N__63496;
    wire N__63495;
    wire N__63494;
    wire N__63489;
    wire N__63486;
    wire N__63485;
    wire N__63482;
    wire N__63479;
    wire N__63476;
    wire N__63473;
    wire N__63468;
    wire N__63465;
    wire N__63462;
    wire N__63457;
    wire N__63456;
    wire N__63455;
    wire N__63452;
    wire N__63449;
    wire N__63446;
    wire N__63441;
    wire N__63438;
    wire N__63435;
    wire N__63432;
    wire N__63429;
    wire N__63426;
    wire N__63423;
    wire N__63418;
    wire N__63417;
    wire N__63416;
    wire N__63415;
    wire N__63414;
    wire N__63413;
    wire N__63412;
    wire N__63409;
    wire N__63404;
    wire N__63399;
    wire N__63396;
    wire N__63395;
    wire N__63394;
    wire N__63391;
    wire N__63390;
    wire N__63389;
    wire N__63386;
    wire N__63381;
    wire N__63380;
    wire N__63379;
    wire N__63378;
    wire N__63377;
    wire N__63374;
    wire N__63371;
    wire N__63368;
    wire N__63365;
    wire N__63362;
    wire N__63359;
    wire N__63358;
    wire N__63357;
    wire N__63356;
    wire N__63355;
    wire N__63354;
    wire N__63353;
    wire N__63348;
    wire N__63343;
    wire N__63340;
    wire N__63337;
    wire N__63334;
    wire N__63331;
    wire N__63328;
    wire N__63325;
    wire N__63318;
    wire N__63315;
    wire N__63312;
    wire N__63305;
    wire N__63300;
    wire N__63295;
    wire N__63292;
    wire N__63287;
    wire N__63282;
    wire N__63281;
    wire N__63280;
    wire N__63273;
    wire N__63270;
    wire N__63265;
    wire N__63260;
    wire N__63257;
    wire N__63254;
    wire N__63251;
    wire N__63246;
    wire N__63243;
    wire N__63232;
    wire N__63231;
    wire N__63228;
    wire N__63225;
    wire N__63224;
    wire N__63219;
    wire N__63218;
    wire N__63215;
    wire N__63212;
    wire N__63209;
    wire N__63202;
    wire N__63201;
    wire N__63198;
    wire N__63197;
    wire N__63194;
    wire N__63191;
    wire N__63188;
    wire N__63181;
    wire N__63180;
    wire N__63175;
    wire N__63172;
    wire N__63169;
    wire N__63166;
    wire N__63163;
    wire N__63162;
    wire N__63159;
    wire N__63156;
    wire N__63155;
    wire N__63150;
    wire N__63149;
    wire N__63148;
    wire N__63145;
    wire N__63142;
    wire N__63139;
    wire N__63136;
    wire N__63135;
    wire N__63132;
    wire N__63129;
    wire N__63124;
    wire N__63121;
    wire N__63118;
    wire N__63109;
    wire N__63106;
    wire N__63105;
    wire N__63104;
    wire N__63101;
    wire N__63100;
    wire N__63099;
    wire N__63096;
    wire N__63093;
    wire N__63090;
    wire N__63087;
    wire N__63084;
    wire N__63081;
    wire N__63070;
    wire N__63067;
    wire N__63066;
    wire N__63065;
    wire N__63062;
    wire N__63057;
    wire N__63054;
    wire N__63049;
    wire N__63048;
    wire N__63045;
    wire N__63044;
    wire N__63041;
    wire N__63038;
    wire N__63035;
    wire N__63034;
    wire N__63031;
    wire N__63028;
    wire N__63025;
    wire N__63022;
    wire N__63013;
    wire N__63010;
    wire N__63007;
    wire N__63004;
    wire N__63001;
    wire N__62998;
    wire N__62995;
    wire N__62992;
    wire N__62989;
    wire N__62988;
    wire N__62985;
    wire N__62982;
    wire N__62981;
    wire N__62976;
    wire N__62973;
    wire N__62970;
    wire N__62969;
    wire N__62968;
    wire N__62965;
    wire N__62962;
    wire N__62957;
    wire N__62950;
    wire N__62947;
    wire N__62944;
    wire N__62941;
    wire N__62938;
    wire N__62935;
    wire N__62934;
    wire N__62931;
    wire N__62928;
    wire N__62927;
    wire N__62926;
    wire N__62923;
    wire N__62916;
    wire N__62911;
    wire N__62908;
    wire N__62905;
    wire N__62904;
    wire N__62901;
    wire N__62898;
    wire N__62895;
    wire N__62890;
    wire N__62889;
    wire N__62886;
    wire N__62885;
    wire N__62882;
    wire N__62879;
    wire N__62878;
    wire N__62875;
    wire N__62872;
    wire N__62869;
    wire N__62866;
    wire N__62863;
    wire N__62858;
    wire N__62855;
    wire N__62848;
    wire N__62847;
    wire N__62846;
    wire N__62845;
    wire N__62844;
    wire N__62839;
    wire N__62838;
    wire N__62837;
    wire N__62834;
    wire N__62831;
    wire N__62830;
    wire N__62827;
    wire N__62824;
    wire N__62819;
    wire N__62816;
    wire N__62813;
    wire N__62812;
    wire N__62811;
    wire N__62810;
    wire N__62807;
    wire N__62804;
    wire N__62803;
    wire N__62802;
    wire N__62801;
    wire N__62798;
    wire N__62795;
    wire N__62794;
    wire N__62793;
    wire N__62788;
    wire N__62785;
    wire N__62782;
    wire N__62779;
    wire N__62774;
    wire N__62771;
    wire N__62766;
    wire N__62763;
    wire N__62760;
    wire N__62755;
    wire N__62752;
    wire N__62743;
    wire N__62734;
    wire N__62725;
    wire N__62724;
    wire N__62721;
    wire N__62720;
    wire N__62717;
    wire N__62716;
    wire N__62713;
    wire N__62710;
    wire N__62705;
    wire N__62698;
    wire N__62695;
    wire N__62692;
    wire N__62689;
    wire N__62686;
    wire N__62683;
    wire N__62682;
    wire N__62681;
    wire N__62680;
    wire N__62679;
    wire N__62676;
    wire N__62673;
    wire N__62670;
    wire N__62667;
    wire N__62664;
    wire N__62659;
    wire N__62658;
    wire N__62655;
    wire N__62650;
    wire N__62647;
    wire N__62644;
    wire N__62635;
    wire N__62632;
    wire N__62629;
    wire N__62626;
    wire N__62625;
    wire N__62624;
    wire N__62621;
    wire N__62620;
    wire N__62619;
    wire N__62618;
    wire N__62615;
    wire N__62612;
    wire N__62609;
    wire N__62606;
    wire N__62601;
    wire N__62596;
    wire N__62587;
    wire N__62584;
    wire N__62583;
    wire N__62582;
    wire N__62579;
    wire N__62576;
    wire N__62573;
    wire N__62570;
    wire N__62567;
    wire N__62564;
    wire N__62561;
    wire N__62556;
    wire N__62551;
    wire N__62548;
    wire N__62545;
    wire N__62544;
    wire N__62541;
    wire N__62538;
    wire N__62535;
    wire N__62532;
    wire N__62527;
    wire N__62524;
    wire N__62523;
    wire N__62522;
    wire N__62519;
    wire N__62516;
    wire N__62513;
    wire N__62512;
    wire N__62507;
    wire N__62502;
    wire N__62497;
    wire N__62496;
    wire N__62495;
    wire N__62492;
    wire N__62489;
    wire N__62486;
    wire N__62483;
    wire N__62480;
    wire N__62477;
    wire N__62474;
    wire N__62467;
    wire N__62466;
    wire N__62465;
    wire N__62464;
    wire N__62461;
    wire N__62456;
    wire N__62453;
    wire N__62448;
    wire N__62447;
    wire N__62444;
    wire N__62441;
    wire N__62440;
    wire N__62437;
    wire N__62434;
    wire N__62431;
    wire N__62428;
    wire N__62419;
    wire N__62418;
    wire N__62415;
    wire N__62412;
    wire N__62411;
    wire N__62410;
    wire N__62409;
    wire N__62406;
    wire N__62403;
    wire N__62400;
    wire N__62399;
    wire N__62396;
    wire N__62393;
    wire N__62386;
    wire N__62383;
    wire N__62382;
    wire N__62379;
    wire N__62374;
    wire N__62371;
    wire N__62368;
    wire N__62359;
    wire N__62356;
    wire N__62355;
    wire N__62354;
    wire N__62353;
    wire N__62350;
    wire N__62347;
    wire N__62344;
    wire N__62343;
    wire N__62340;
    wire N__62335;
    wire N__62332;
    wire N__62329;
    wire N__62320;
    wire N__62317;
    wire N__62314;
    wire N__62313;
    wire N__62310;
    wire N__62309;
    wire N__62308;
    wire N__62307;
    wire N__62304;
    wire N__62301;
    wire N__62298;
    wire N__62293;
    wire N__62290;
    wire N__62287;
    wire N__62284;
    wire N__62281;
    wire N__62278;
    wire N__62275;
    wire N__62270;
    wire N__62267;
    wire N__62264;
    wire N__62257;
    wire N__62256;
    wire N__62255;
    wire N__62254;
    wire N__62251;
    wire N__62250;
    wire N__62247;
    wire N__62244;
    wire N__62241;
    wire N__62238;
    wire N__62235;
    wire N__62232;
    wire N__62229;
    wire N__62226;
    wire N__62223;
    wire N__62218;
    wire N__62215;
    wire N__62206;
    wire N__62203;
    wire N__62200;
    wire N__62199;
    wire N__62198;
    wire N__62197;
    wire N__62194;
    wire N__62187;
    wire N__62182;
    wire N__62181;
    wire N__62180;
    wire N__62177;
    wire N__62176;
    wire N__62173;
    wire N__62172;
    wire N__62169;
    wire N__62166;
    wire N__62165;
    wire N__62164;
    wire N__62163;
    wire N__62160;
    wire N__62157;
    wire N__62156;
    wire N__62153;
    wire N__62148;
    wire N__62145;
    wire N__62140;
    wire N__62135;
    wire N__62132;
    wire N__62131;
    wire N__62130;
    wire N__62129;
    wire N__62128;
    wire N__62127;
    wire N__62126;
    wire N__62123;
    wire N__62118;
    wire N__62111;
    wire N__62108;
    wire N__62105;
    wire N__62100;
    wire N__62095;
    wire N__62080;
    wire N__62077;
    wire N__62076;
    wire N__62073;
    wire N__62070;
    wire N__62067;
    wire N__62062;
    wire N__62059;
    wire N__62058;
    wire N__62053;
    wire N__62050;
    wire N__62049;
    wire N__62048;
    wire N__62045;
    wire N__62042;
    wire N__62041;
    wire N__62040;
    wire N__62039;
    wire N__62036;
    wire N__62035;
    wire N__62034;
    wire N__62031;
    wire N__62030;
    wire N__62027;
    wire N__62024;
    wire N__62019;
    wire N__62018;
    wire N__62013;
    wire N__62010;
    wire N__62009;
    wire N__62006;
    wire N__62003;
    wire N__62002;
    wire N__61997;
    wire N__61994;
    wire N__61991;
    wire N__61988;
    wire N__61987;
    wire N__61984;
    wire N__61981;
    wire N__61976;
    wire N__61973;
    wire N__61968;
    wire N__61965;
    wire N__61962;
    wire N__61959;
    wire N__61956;
    wire N__61955;
    wire N__61954;
    wire N__61951;
    wire N__61948;
    wire N__61945;
    wire N__61942;
    wire N__61937;
    wire N__61934;
    wire N__61931;
    wire N__61928;
    wire N__61927;
    wire N__61924;
    wire N__61921;
    wire N__61916;
    wire N__61911;
    wire N__61904;
    wire N__61901;
    wire N__61898;
    wire N__61893;
    wire N__61888;
    wire N__61879;
    wire N__61878;
    wire N__61875;
    wire N__61874;
    wire N__61873;
    wire N__61872;
    wire N__61871;
    wire N__61868;
    wire N__61865;
    wire N__61862;
    wire N__61861;
    wire N__61860;
    wire N__61857;
    wire N__61852;
    wire N__61847;
    wire N__61844;
    wire N__61841;
    wire N__61838;
    wire N__61833;
    wire N__61830;
    wire N__61827;
    wire N__61826;
    wire N__61823;
    wire N__61820;
    wire N__61813;
    wire N__61810;
    wire N__61801;
    wire N__61798;
    wire N__61797;
    wire N__61796;
    wire N__61795;
    wire N__61794;
    wire N__61791;
    wire N__61786;
    wire N__61781;
    wire N__61780;
    wire N__61779;
    wire N__61778;
    wire N__61777;
    wire N__61774;
    wire N__61769;
    wire N__61768;
    wire N__61767;
    wire N__61766;
    wire N__61761;
    wire N__61760;
    wire N__61759;
    wire N__61758;
    wire N__61757;
    wire N__61756;
    wire N__61755;
    wire N__61754;
    wire N__61753;
    wire N__61752;
    wire N__61749;
    wire N__61746;
    wire N__61745;
    wire N__61744;
    wire N__61739;
    wire N__61732;
    wire N__61731;
    wire N__61730;
    wire N__61727;
    wire N__61726;
    wire N__61725;
    wire N__61724;
    wire N__61723;
    wire N__61716;
    wire N__61713;
    wire N__61702;
    wire N__61693;
    wire N__61692;
    wire N__61691;
    wire N__61690;
    wire N__61689;
    wire N__61688;
    wire N__61687;
    wire N__61686;
    wire N__61685;
    wire N__61684;
    wire N__61683;
    wire N__61678;
    wire N__61677;
    wire N__61674;
    wire N__61673;
    wire N__61672;
    wire N__61671;
    wire N__61670;
    wire N__61667;
    wire N__61664;
    wire N__61659;
    wire N__61654;
    wire N__61651;
    wire N__61644;
    wire N__61635;
    wire N__61632;
    wire N__61627;
    wire N__61624;
    wire N__61619;
    wire N__61616;
    wire N__61615;
    wire N__61612;
    wire N__61609;
    wire N__61600;
    wire N__61599;
    wire N__61598;
    wire N__61597;
    wire N__61596;
    wire N__61595;
    wire N__61594;
    wire N__61593;
    wire N__61584;
    wire N__61577;
    wire N__61572;
    wire N__61567;
    wire N__61564;
    wire N__61561;
    wire N__61560;
    wire N__61553;
    wire N__61552;
    wire N__61551;
    wire N__61550;
    wire N__61549;
    wire N__61546;
    wire N__61543;
    wire N__61538;
    wire N__61531;
    wire N__61522;
    wire N__61519;
    wire N__61516;
    wire N__61513;
    wire N__61510;
    wire N__61501;
    wire N__61498;
    wire N__61485;
    wire N__61478;
    wire N__61475;
    wire N__61472;
    wire N__61469;
    wire N__61466;
    wire N__61461;
    wire N__61456;
    wire N__61455;
    wire N__61454;
    wire N__61453;
    wire N__61450;
    wire N__61449;
    wire N__61448;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61434;
    wire N__61431;
    wire N__61430;
    wire N__61425;
    wire N__61424;
    wire N__61421;
    wire N__61418;
    wire N__61415;
    wire N__61412;
    wire N__61409;
    wire N__61408;
    wire N__61407;
    wire N__61404;
    wire N__61401;
    wire N__61398;
    wire N__61395;
    wire N__61392;
    wire N__61389;
    wire N__61384;
    wire N__61381;
    wire N__61378;
    wire N__61373;
    wire N__61368;
    wire N__61361;
    wire N__61354;
    wire N__61351;
    wire N__61348;
    wire N__61347;
    wire N__61346;
    wire N__61345;
    wire N__61342;
    wire N__61337;
    wire N__61334;
    wire N__61331;
    wire N__61328;
    wire N__61327;
    wire N__61326;
    wire N__61323;
    wire N__61318;
    wire N__61313;
    wire N__61306;
    wire N__61303;
    wire N__61300;
    wire N__61297;
    wire N__61294;
    wire N__61291;
    wire N__61288;
    wire N__61285;
    wire N__61284;
    wire N__61281;
    wire N__61278;
    wire N__61275;
    wire N__61272;
    wire N__61269;
    wire N__61266;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61254;
    wire N__61251;
    wire N__61248;
    wire N__61247;
    wire N__61246;
    wire N__61241;
    wire N__61236;
    wire N__61231;
    wire N__61228;
    wire N__61227;
    wire N__61226;
    wire N__61225;
    wire N__61222;
    wire N__61219;
    wire N__61216;
    wire N__61213;
    wire N__61212;
    wire N__61209;
    wire N__61206;
    wire N__61205;
    wire N__61202;
    wire N__61199;
    wire N__61198;
    wire N__61197;
    wire N__61196;
    wire N__61195;
    wire N__61194;
    wire N__61193;
    wire N__61190;
    wire N__61187;
    wire N__61184;
    wire N__61181;
    wire N__61176;
    wire N__61173;
    wire N__61170;
    wire N__61163;
    wire N__61160;
    wire N__61141;
    wire N__61138;
    wire N__61135;
    wire N__61132;
    wire N__61131;
    wire N__61128;
    wire N__61127;
    wire N__61126;
    wire N__61123;
    wire N__61122;
    wire N__61119;
    wire N__61118;
    wire N__61117;
    wire N__61112;
    wire N__61109;
    wire N__61106;
    wire N__61103;
    wire N__61100;
    wire N__61099;
    wire N__61096;
    wire N__61093;
    wire N__61092;
    wire N__61087;
    wire N__61082;
    wire N__61081;
    wire N__61080;
    wire N__61079;
    wire N__61078;
    wire N__61077;
    wire N__61074;
    wire N__61073;
    wire N__61070;
    wire N__61067;
    wire N__61064;
    wire N__61061;
    wire N__61058;
    wire N__61055;
    wire N__61048;
    wire N__61045;
    wire N__61040;
    wire N__61033;
    wire N__61018;
    wire N__61015;
    wire N__61012;
    wire N__61011;
    wire N__61008;
    wire N__61005;
    wire N__61002;
    wire N__60999;
    wire N__60994;
    wire N__60991;
    wire N__60988;
    wire N__60987;
    wire N__60984;
    wire N__60983;
    wire N__60980;
    wire N__60977;
    wire N__60976;
    wire N__60973;
    wire N__60970;
    wire N__60967;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60957;
    wire N__60956;
    wire N__60953;
    wire N__60950;
    wire N__60945;
    wire N__60940;
    wire N__60931;
    wire N__60928;
    wire N__60927;
    wire N__60926;
    wire N__60923;
    wire N__60922;
    wire N__60917;
    wire N__60916;
    wire N__60913;
    wire N__60910;
    wire N__60909;
    wire N__60908;
    wire N__60907;
    wire N__60906;
    wire N__60905;
    wire N__60902;
    wire N__60901;
    wire N__60900;
    wire N__60899;
    wire N__60896;
    wire N__60893;
    wire N__60890;
    wire N__60887;
    wire N__60884;
    wire N__60881;
    wire N__60876;
    wire N__60873;
    wire N__60868;
    wire N__60865;
    wire N__60844;
    wire N__60843;
    wire N__60842;
    wire N__60839;
    wire N__60836;
    wire N__60833;
    wire N__60830;
    wire N__60829;
    wire N__60826;
    wire N__60823;
    wire N__60820;
    wire N__60817;
    wire N__60814;
    wire N__60811;
    wire N__60808;
    wire N__60805;
    wire N__60802;
    wire N__60793;
    wire N__60792;
    wire N__60791;
    wire N__60788;
    wire N__60785;
    wire N__60782;
    wire N__60779;
    wire N__60778;
    wire N__60775;
    wire N__60772;
    wire N__60771;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60756;
    wire N__60745;
    wire N__60742;
    wire N__60739;
    wire N__60736;
    wire N__60733;
    wire N__60730;
    wire N__60729;
    wire N__60726;
    wire N__60723;
    wire N__60718;
    wire N__60717;
    wire N__60714;
    wire N__60711;
    wire N__60710;
    wire N__60709;
    wire N__60704;
    wire N__60699;
    wire N__60696;
    wire N__60695;
    wire N__60694;
    wire N__60693;
    wire N__60692;
    wire N__60691;
    wire N__60690;
    wire N__60689;
    wire N__60688;
    wire N__60687;
    wire N__60686;
    wire N__60683;
    wire N__60680;
    wire N__60677;
    wire N__60668;
    wire N__60663;
    wire N__60660;
    wire N__60655;
    wire N__60654;
    wire N__60653;
    wire N__60652;
    wire N__60651;
    wire N__60650;
    wire N__60647;
    wire N__60644;
    wire N__60641;
    wire N__60636;
    wire N__60635;
    wire N__60634;
    wire N__60633;
    wire N__60632;
    wire N__60629;
    wire N__60626;
    wire N__60621;
    wire N__60620;
    wire N__60619;
    wire N__60618;
    wire N__60617;
    wire N__60612;
    wire N__60609;
    wire N__60606;
    wire N__60603;
    wire N__60600;
    wire N__60597;
    wire N__60592;
    wire N__60589;
    wire N__60586;
    wire N__60585;
    wire N__60584;
    wire N__60583;
    wire N__60576;
    wire N__60567;
    wire N__60560;
    wire N__60555;
    wire N__60552;
    wire N__60549;
    wire N__60546;
    wire N__60543;
    wire N__60538;
    wire N__60535;
    wire N__60528;
    wire N__60511;
    wire N__60508;
    wire N__60505;
    wire N__60502;
    wire N__60499;
    wire N__60496;
    wire N__60493;
    wire N__60492;
    wire N__60489;
    wire N__60488;
    wire N__60487;
    wire N__60482;
    wire N__60479;
    wire N__60478;
    wire N__60475;
    wire N__60472;
    wire N__60469;
    wire N__60466;
    wire N__60461;
    wire N__60458;
    wire N__60451;
    wire N__60450;
    wire N__60449;
    wire N__60448;
    wire N__60445;
    wire N__60442;
    wire N__60439;
    wire N__60436;
    wire N__60433;
    wire N__60430;
    wire N__60427;
    wire N__60422;
    wire N__60419;
    wire N__60412;
    wire N__60411;
    wire N__60408;
    wire N__60405;
    wire N__60402;
    wire N__60399;
    wire N__60398;
    wire N__60395;
    wire N__60392;
    wire N__60391;
    wire N__60390;
    wire N__60389;
    wire N__60388;
    wire N__60385;
    wire N__60382;
    wire N__60379;
    wire N__60372;
    wire N__60369;
    wire N__60358;
    wire N__60355;
    wire N__60354;
    wire N__60353;
    wire N__60352;
    wire N__60347;
    wire N__60346;
    wire N__60343;
    wire N__60340;
    wire N__60337;
    wire N__60336;
    wire N__60333;
    wire N__60330;
    wire N__60329;
    wire N__60326;
    wire N__60323;
    wire N__60320;
    wire N__60319;
    wire N__60316;
    wire N__60313;
    wire N__60310;
    wire N__60309;
    wire N__60302;
    wire N__60299;
    wire N__60296;
    wire N__60293;
    wire N__60288;
    wire N__60281;
    wire N__60274;
    wire N__60273;
    wire N__60272;
    wire N__60269;
    wire N__60268;
    wire N__60265;
    wire N__60264;
    wire N__60263;
    wire N__60260;
    wire N__60257;
    wire N__60256;
    wire N__60253;
    wire N__60252;
    wire N__60249;
    wire N__60246;
    wire N__60243;
    wire N__60242;
    wire N__60239;
    wire N__60236;
    wire N__60235;
    wire N__60232;
    wire N__60229;
    wire N__60226;
    wire N__60223;
    wire N__60220;
    wire N__60215;
    wire N__60212;
    wire N__60209;
    wire N__60208;
    wire N__60205;
    wire N__60204;
    wire N__60201;
    wire N__60198;
    wire N__60195;
    wire N__60192;
    wire N__60189;
    wire N__60186;
    wire N__60183;
    wire N__60180;
    wire N__60177;
    wire N__60174;
    wire N__60171;
    wire N__60168;
    wire N__60163;
    wire N__60154;
    wire N__60151;
    wire N__60148;
    wire N__60133;
    wire N__60132;
    wire N__60129;
    wire N__60128;
    wire N__60125;
    wire N__60122;
    wire N__60121;
    wire N__60118;
    wire N__60117;
    wire N__60116;
    wire N__60115;
    wire N__60112;
    wire N__60109;
    wire N__60108;
    wire N__60105;
    wire N__60104;
    wire N__60101;
    wire N__60098;
    wire N__60095;
    wire N__60092;
    wire N__60089;
    wire N__60086;
    wire N__60083;
    wire N__60080;
    wire N__60077;
    wire N__60072;
    wire N__60069;
    wire N__60064;
    wire N__60061;
    wire N__60058;
    wire N__60053;
    wire N__60050;
    wire N__60049;
    wire N__60048;
    wire N__60047;
    wire N__60042;
    wire N__60041;
    wire N__60038;
    wire N__60035;
    wire N__60032;
    wire N__60029;
    wire N__60022;
    wire N__60019;
    wire N__60016;
    wire N__60001;
    wire N__60000;
    wire N__59997;
    wire N__59996;
    wire N__59993;
    wire N__59992;
    wire N__59989;
    wire N__59986;
    wire N__59985;
    wire N__59982;
    wire N__59979;
    wire N__59978;
    wire N__59977;
    wire N__59972;
    wire N__59969;
    wire N__59966;
    wire N__59965;
    wire N__59962;
    wire N__59959;
    wire N__59956;
    wire N__59951;
    wire N__59948;
    wire N__59945;
    wire N__59944;
    wire N__59939;
    wire N__59934;
    wire N__59931;
    wire N__59928;
    wire N__59927;
    wire N__59924;
    wire N__59923;
    wire N__59922;
    wire N__59921;
    wire N__59914;
    wire N__59911;
    wire N__59908;
    wire N__59899;
    wire N__59896;
    wire N__59893;
    wire N__59884;
    wire N__59883;
    wire N__59880;
    wire N__59877;
    wire N__59876;
    wire N__59875;
    wire N__59870;
    wire N__59869;
    wire N__59868;
    wire N__59867;
    wire N__59866;
    wire N__59861;
    wire N__59858;
    wire N__59855;
    wire N__59848;
    wire N__59845;
    wire N__59842;
    wire N__59833;
    wire N__59832;
    wire N__59829;
    wire N__59828;
    wire N__59825;
    wire N__59822;
    wire N__59819;
    wire N__59812;
    wire N__59809;
    wire N__59806;
    wire N__59803;
    wire N__59800;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59784;
    wire N__59783;
    wire N__59780;
    wire N__59779;
    wire N__59776;
    wire N__59775;
    wire N__59772;
    wire N__59769;
    wire N__59766;
    wire N__59763;
    wire N__59760;
    wire N__59757;
    wire N__59748;
    wire N__59743;
    wire N__59742;
    wire N__59739;
    wire N__59738;
    wire N__59735;
    wire N__59732;
    wire N__59729;
    wire N__59726;
    wire N__59723;
    wire N__59720;
    wire N__59719;
    wire N__59712;
    wire N__59709;
    wire N__59706;
    wire N__59701;
    wire N__59700;
    wire N__59699;
    wire N__59696;
    wire N__59693;
    wire N__59692;
    wire N__59689;
    wire N__59688;
    wire N__59685;
    wire N__59682;
    wire N__59679;
    wire N__59676;
    wire N__59673;
    wire N__59670;
    wire N__59669;
    wire N__59666;
    wire N__59663;
    wire N__59660;
    wire N__59657;
    wire N__59654;
    wire N__59651;
    wire N__59644;
    wire N__59639;
    wire N__59636;
    wire N__59633;
    wire N__59630;
    wire N__59623;
    wire N__59620;
    wire N__59617;
    wire N__59616;
    wire N__59613;
    wire N__59612;
    wire N__59609;
    wire N__59606;
    wire N__59603;
    wire N__59596;
    wire N__59595;
    wire N__59592;
    wire N__59589;
    wire N__59588;
    wire N__59585;
    wire N__59582;
    wire N__59579;
    wire N__59576;
    wire N__59571;
    wire N__59568;
    wire N__59565;
    wire N__59560;
    wire N__59557;
    wire N__59556;
    wire N__59553;
    wire N__59550;
    wire N__59549;
    wire N__59548;
    wire N__59545;
    wire N__59540;
    wire N__59537;
    wire N__59530;
    wire N__59527;
    wire N__59524;
    wire N__59521;
    wire N__59518;
    wire N__59515;
    wire N__59512;
    wire N__59511;
    wire N__59508;
    wire N__59505;
    wire N__59504;
    wire N__59501;
    wire N__59498;
    wire N__59495;
    wire N__59488;
    wire N__59485;
    wire N__59482;
    wire N__59481;
    wire N__59480;
    wire N__59479;
    wire N__59478;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59466;
    wire N__59463;
    wire N__59460;
    wire N__59459;
    wire N__59456;
    wire N__59455;
    wire N__59452;
    wire N__59449;
    wire N__59448;
    wire N__59443;
    wire N__59440;
    wire N__59439;
    wire N__59436;
    wire N__59433;
    wire N__59432;
    wire N__59429;
    wire N__59426;
    wire N__59423;
    wire N__59418;
    wire N__59415;
    wire N__59412;
    wire N__59409;
    wire N__59406;
    wire N__59403;
    wire N__59396;
    wire N__59393;
    wire N__59380;
    wire N__59377;
    wire N__59374;
    wire N__59371;
    wire N__59368;
    wire N__59365;
    wire N__59362;
    wire N__59359;
    wire N__59358;
    wire N__59355;
    wire N__59352;
    wire N__59349;
    wire N__59346;
    wire N__59345;
    wire N__59340;
    wire N__59337;
    wire N__59332;
    wire N__59329;
    wire N__59326;
    wire N__59325;
    wire N__59324;
    wire N__59321;
    wire N__59318;
    wire N__59315;
    wire N__59312;
    wire N__59307;
    wire N__59302;
    wire N__59301;
    wire N__59300;
    wire N__59297;
    wire N__59294;
    wire N__59291;
    wire N__59288;
    wire N__59285;
    wire N__59282;
    wire N__59279;
    wire N__59276;
    wire N__59275;
    wire N__59274;
    wire N__59269;
    wire N__59266;
    wire N__59261;
    wire N__59254;
    wire N__59251;
    wire N__59250;
    wire N__59247;
    wire N__59244;
    wire N__59241;
    wire N__59238;
    wire N__59237;
    wire N__59232;
    wire N__59231;
    wire N__59230;
    wire N__59227;
    wire N__59224;
    wire N__59219;
    wire N__59212;
    wire N__59211;
    wire N__59208;
    wire N__59205;
    wire N__59202;
    wire N__59199;
    wire N__59196;
    wire N__59191;
    wire N__59190;
    wire N__59187;
    wire N__59184;
    wire N__59179;
    wire N__59178;
    wire N__59175;
    wire N__59172;
    wire N__59169;
    wire N__59166;
    wire N__59165;
    wire N__59162;
    wire N__59159;
    wire N__59156;
    wire N__59149;
    wire N__59146;
    wire N__59143;
    wire N__59140;
    wire N__59137;
    wire N__59134;
    wire N__59133;
    wire N__59130;
    wire N__59127;
    wire N__59126;
    wire N__59123;
    wire N__59120;
    wire N__59117;
    wire N__59116;
    wire N__59115;
    wire N__59112;
    wire N__59107;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59086;
    wire N__59085;
    wire N__59082;
    wire N__59079;
    wire N__59076;
    wire N__59075;
    wire N__59074;
    wire N__59073;
    wire N__59072;
    wire N__59069;
    wire N__59066;
    wire N__59061;
    wire N__59056;
    wire N__59047;
    wire N__59046;
    wire N__59043;
    wire N__59040;
    wire N__59039;
    wire N__59036;
    wire N__59033;
    wire N__59032;
    wire N__59029;
    wire N__59024;
    wire N__59021;
    wire N__59014;
    wire N__59011;
    wire N__59010;
    wire N__59009;
    wire N__59006;
    wire N__59005;
    wire N__59004;
    wire N__59003;
    wire N__59002;
    wire N__58999;
    wire N__58998;
    wire N__58995;
    wire N__58992;
    wire N__58985;
    wire N__58982;
    wire N__58979;
    wire N__58976;
    wire N__58967;
    wire N__58962;
    wire N__58959;
    wire N__58954;
    wire N__58951;
    wire N__58948;
    wire N__58945;
    wire N__58942;
    wire N__58941;
    wire N__58940;
    wire N__58937;
    wire N__58932;
    wire N__58931;
    wire N__58926;
    wire N__58923;
    wire N__58920;
    wire N__58917;
    wire N__58912;
    wire N__58909;
    wire N__58906;
    wire N__58903;
    wire N__58900;
    wire N__58899;
    wire N__58896;
    wire N__58895;
    wire N__58892;
    wire N__58889;
    wire N__58886;
    wire N__58883;
    wire N__58878;
    wire N__58875;
    wire N__58872;
    wire N__58871;
    wire N__58868;
    wire N__58865;
    wire N__58862;
    wire N__58859;
    wire N__58856;
    wire N__58849;
    wire N__58846;
    wire N__58843;
    wire N__58840;
    wire N__58839;
    wire N__58836;
    wire N__58833;
    wire N__58832;
    wire N__58829;
    wire N__58826;
    wire N__58823;
    wire N__58822;
    wire N__58819;
    wire N__58814;
    wire N__58811;
    wire N__58808;
    wire N__58805;
    wire N__58798;
    wire N__58795;
    wire N__58794;
    wire N__58791;
    wire N__58790;
    wire N__58787;
    wire N__58784;
    wire N__58781;
    wire N__58778;
    wire N__58775;
    wire N__58768;
    wire N__58765;
    wire N__58762;
    wire N__58761;
    wire N__58760;
    wire N__58757;
    wire N__58756;
    wire N__58753;
    wire N__58750;
    wire N__58747;
    wire N__58744;
    wire N__58741;
    wire N__58738;
    wire N__58735;
    wire N__58726;
    wire N__58725;
    wire N__58724;
    wire N__58719;
    wire N__58716;
    wire N__58715;
    wire N__58712;
    wire N__58709;
    wire N__58708;
    wire N__58705;
    wire N__58700;
    wire N__58697;
    wire N__58694;
    wire N__58691;
    wire N__58688;
    wire N__58685;
    wire N__58682;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58668;
    wire N__58667;
    wire N__58664;
    wire N__58661;
    wire N__58658;
    wire N__58655;
    wire N__58650;
    wire N__58649;
    wire N__58646;
    wire N__58643;
    wire N__58640;
    wire N__58633;
    wire N__58630;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58620;
    wire N__58617;
    wire N__58612;
    wire N__58609;
    wire N__58606;
    wire N__58603;
    wire N__58600;
    wire N__58599;
    wire N__58598;
    wire N__58595;
    wire N__58592;
    wire N__58589;
    wire N__58582;
    wire N__58579;
    wire N__58576;
    wire N__58573;
    wire N__58570;
    wire N__58567;
    wire N__58564;
    wire N__58561;
    wire N__58558;
    wire N__58555;
    wire N__58552;
    wire N__58551;
    wire N__58550;
    wire N__58547;
    wire N__58544;
    wire N__58541;
    wire N__58538;
    wire N__58535;
    wire N__58532;
    wire N__58529;
    wire N__58526;
    wire N__58523;
    wire N__58518;
    wire N__58515;
    wire N__58510;
    wire N__58507;
    wire N__58506;
    wire N__58503;
    wire N__58500;
    wire N__58495;
    wire N__58492;
    wire N__58491;
    wire N__58488;
    wire N__58485;
    wire N__58482;
    wire N__58479;
    wire N__58476;
    wire N__58473;
    wire N__58468;
    wire N__58467;
    wire N__58466;
    wire N__58463;
    wire N__58462;
    wire N__58461;
    wire N__58458;
    wire N__58455;
    wire N__58452;
    wire N__58449;
    wire N__58446;
    wire N__58443;
    wire N__58440;
    wire N__58433;
    wire N__58432;
    wire N__58431;
    wire N__58428;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58408;
    wire N__58405;
    wire N__58404;
    wire N__58401;
    wire N__58398;
    wire N__58395;
    wire N__58392;
    wire N__58387;
    wire N__58384;
    wire N__58381;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58369;
    wire N__58368;
    wire N__58365;
    wire N__58362;
    wire N__58359;
    wire N__58354;
    wire N__58353;
    wire N__58350;
    wire N__58347;
    wire N__58342;
    wire N__58339;
    wire N__58336;
    wire N__58335;
    wire N__58330;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58309;
    wire N__58306;
    wire N__58305;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58287;
    wire N__58284;
    wire N__58281;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58255;
    wire N__58252;
    wire N__58249;
    wire N__58248;
    wire N__58247;
    wire N__58244;
    wire N__58239;
    wire N__58236;
    wire N__58233;
    wire N__58228;
    wire N__58227;
    wire N__58224;
    wire N__58221;
    wire N__58218;
    wire N__58217;
    wire N__58212;
    wire N__58209;
    wire N__58204;
    wire N__58201;
    wire N__58200;
    wire N__58199;
    wire N__58194;
    wire N__58191;
    wire N__58186;
    wire N__58183;
    wire N__58180;
    wire N__58177;
    wire N__58174;
    wire N__58171;
    wire N__58168;
    wire N__58165;
    wire N__58162;
    wire N__58159;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58147;
    wire N__58144;
    wire N__58141;
    wire N__58138;
    wire N__58135;
    wire N__58132;
    wire N__58131;
    wire N__58130;
    wire N__58127;
    wire N__58124;
    wire N__58121;
    wire N__58114;
    wire N__58111;
    wire N__58108;
    wire N__58105;
    wire N__58102;
    wire N__58099;
    wire N__58098;
    wire N__58097;
    wire N__58094;
    wire N__58089;
    wire N__58084;
    wire N__58081;
    wire N__58078;
    wire N__58075;
    wire N__58072;
    wire N__58069;
    wire N__58068;
    wire N__58067;
    wire N__58064;
    wire N__58059;
    wire N__58054;
    wire N__58053;
    wire N__58050;
    wire N__58047;
    wire N__58042;
    wire N__58041;
    wire N__58038;
    wire N__58037;
    wire N__58034;
    wire N__58031;
    wire N__58028;
    wire N__58025;
    wire N__58024;
    wire N__58017;
    wire N__58014;
    wire N__58009;
    wire N__58006;
    wire N__58003;
    wire N__58000;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57987;
    wire N__57982;
    wire N__57979;
    wire N__57976;
    wire N__57973;
    wire N__57970;
    wire N__57969;
    wire N__57966;
    wire N__57963;
    wire N__57960;
    wire N__57957;
    wire N__57952;
    wire N__57951;
    wire N__57948;
    wire N__57945;
    wire N__57940;
    wire N__57937;
    wire N__57934;
    wire N__57931;
    wire N__57928;
    wire N__57925;
    wire N__57922;
    wire N__57921;
    wire N__57916;
    wire N__57913;
    wire N__57910;
    wire N__57909;
    wire N__57906;
    wire N__57903;
    wire N__57900;
    wire N__57897;
    wire N__57894;
    wire N__57889;
    wire N__57886;
    wire N__57883;
    wire N__57882;
    wire N__57879;
    wire N__57876;
    wire N__57871;
    wire N__57868;
    wire N__57865;
    wire N__57862;
    wire N__57859;
    wire N__57858;
    wire N__57857;
    wire N__57854;
    wire N__57849;
    wire N__57846;
    wire N__57841;
    wire N__57838;
    wire N__57837;
    wire N__57834;
    wire N__57831;
    wire N__57828;
    wire N__57825;
    wire N__57820;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57802;
    wire N__57799;
    wire N__57796;
    wire N__57793;
    wire N__57790;
    wire N__57789;
    wire N__57786;
    wire N__57783;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57766;
    wire N__57763;
    wire N__57760;
    wire N__57757;
    wire N__57754;
    wire N__57751;
    wire N__57748;
    wire N__57747;
    wire N__57744;
    wire N__57741;
    wire N__57736;
    wire N__57733;
    wire N__57732;
    wire N__57729;
    wire N__57726;
    wire N__57725;
    wire N__57724;
    wire N__57723;
    wire N__57720;
    wire N__57717;
    wire N__57714;
    wire N__57713;
    wire N__57710;
    wire N__57709;
    wire N__57706;
    wire N__57701;
    wire N__57698;
    wire N__57693;
    wire N__57692;
    wire N__57689;
    wire N__57682;
    wire N__57679;
    wire N__57676;
    wire N__57673;
    wire N__57670;
    wire N__57667;
    wire N__57658;
    wire N__57657;
    wire N__57656;
    wire N__57655;
    wire N__57652;
    wire N__57647;
    wire N__57646;
    wire N__57645;
    wire N__57642;
    wire N__57637;
    wire N__57634;
    wire N__57633;
    wire N__57632;
    wire N__57629;
    wire N__57626;
    wire N__57623;
    wire N__57620;
    wire N__57617;
    wire N__57614;
    wire N__57611;
    wire N__57606;
    wire N__57603;
    wire N__57600;
    wire N__57589;
    wire N__57586;
    wire N__57583;
    wire N__57582;
    wire N__57581;
    wire N__57578;
    wire N__57573;
    wire N__57572;
    wire N__57571;
    wire N__57568;
    wire N__57565;
    wire N__57562;
    wire N__57559;
    wire N__57552;
    wire N__57547;
    wire N__57544;
    wire N__57541;
    wire N__57538;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57525;
    wire N__57522;
    wire N__57519;
    wire N__57514;
    wire N__57511;
    wire N__57508;
    wire N__57505;
    wire N__57502;
    wire N__57501;
    wire N__57500;
    wire N__57499;
    wire N__57496;
    wire N__57493;
    wire N__57490;
    wire N__57487;
    wire N__57484;
    wire N__57481;
    wire N__57478;
    wire N__57475;
    wire N__57472;
    wire N__57467;
    wire N__57460;
    wire N__57457;
    wire N__57456;
    wire N__57455;
    wire N__57454;
    wire N__57447;
    wire N__57444;
    wire N__57443;
    wire N__57438;
    wire N__57435;
    wire N__57434;
    wire N__57429;
    wire N__57426;
    wire N__57423;
    wire N__57420;
    wire N__57417;
    wire N__57412;
    wire N__57409;
    wire N__57408;
    wire N__57405;
    wire N__57402;
    wire N__57401;
    wire N__57398;
    wire N__57395;
    wire N__57392;
    wire N__57389;
    wire N__57384;
    wire N__57379;
    wire N__57376;
    wire N__57373;
    wire N__57372;
    wire N__57371;
    wire N__57368;
    wire N__57365;
    wire N__57362;
    wire N__57361;
    wire N__57358;
    wire N__57355;
    wire N__57352;
    wire N__57349;
    wire N__57346;
    wire N__57343;
    wire N__57340;
    wire N__57331;
    wire N__57330;
    wire N__57329;
    wire N__57328;
    wire N__57325;
    wire N__57322;
    wire N__57317;
    wire N__57314;
    wire N__57309;
    wire N__57308;
    wire N__57307;
    wire N__57302;
    wire N__57299;
    wire N__57296;
    wire N__57289;
    wire N__57286;
    wire N__57283;
    wire N__57280;
    wire N__57277;
    wire N__57274;
    wire N__57271;
    wire N__57268;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57256;
    wire N__57255;
    wire N__57252;
    wire N__57251;
    wire N__57248;
    wire N__57245;
    wire N__57242;
    wire N__57239;
    wire N__57236;
    wire N__57235;
    wire N__57232;
    wire N__57229;
    wire N__57226;
    wire N__57225;
    wire N__57222;
    wire N__57219;
    wire N__57216;
    wire N__57213;
    wire N__57208;
    wire N__57205;
    wire N__57196;
    wire N__57195;
    wire N__57192;
    wire N__57191;
    wire N__57188;
    wire N__57187;
    wire N__57184;
    wire N__57181;
    wire N__57178;
    wire N__57175;
    wire N__57170;
    wire N__57165;
    wire N__57162;
    wire N__57157;
    wire N__57154;
    wire N__57153;
    wire N__57152;
    wire N__57149;
    wire N__57144;
    wire N__57143;
    wire N__57142;
    wire N__57139;
    wire N__57136;
    wire N__57133;
    wire N__57130;
    wire N__57121;
    wire N__57118;
    wire N__57115;
    wire N__57114;
    wire N__57111;
    wire N__57108;
    wire N__57107;
    wire N__57104;
    wire N__57103;
    wire N__57098;
    wire N__57095;
    wire N__57092;
    wire N__57091;
    wire N__57084;
    wire N__57081;
    wire N__57076;
    wire N__57075;
    wire N__57072;
    wire N__57071;
    wire N__57068;
    wire N__57065;
    wire N__57062;
    wire N__57059;
    wire N__57056;
    wire N__57051;
    wire N__57046;
    wire N__57045;
    wire N__57044;
    wire N__57043;
    wire N__57040;
    wire N__57037;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57025;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57013;
    wire N__57010;
    wire N__57007;
    wire N__57006;
    wire N__57005;
    wire N__57004;
    wire N__57001;
    wire N__56998;
    wire N__56993;
    wire N__56988;
    wire N__56985;
    wire N__56974;
    wire N__56971;
    wire N__56970;
    wire N__56967;
    wire N__56964;
    wire N__56961;
    wire N__56958;
    wire N__56957;
    wire N__56954;
    wire N__56951;
    wire N__56948;
    wire N__56941;
    wire N__56940;
    wire N__56939;
    wire N__56938;
    wire N__56933;
    wire N__56930;
    wire N__56927;
    wire N__56922;
    wire N__56917;
    wire N__56914;
    wire N__56911;
    wire N__56908;
    wire N__56905;
    wire N__56904;
    wire N__56903;
    wire N__56902;
    wire N__56899;
    wire N__56896;
    wire N__56891;
    wire N__56888;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56869;
    wire N__56866;
    wire N__56863;
    wire N__56860;
    wire N__56857;
    wire N__56854;
    wire N__56853;
    wire N__56852;
    wire N__56849;
    wire N__56848;
    wire N__56847;
    wire N__56846;
    wire N__56843;
    wire N__56840;
    wire N__56837;
    wire N__56834;
    wire N__56831;
    wire N__56830;
    wire N__56829;
    wire N__56826;
    wire N__56825;
    wire N__56824;
    wire N__56823;
    wire N__56818;
    wire N__56811;
    wire N__56810;
    wire N__56807;
    wire N__56804;
    wire N__56803;
    wire N__56802;
    wire N__56801;
    wire N__56800;
    wire N__56797;
    wire N__56794;
    wire N__56791;
    wire N__56788;
    wire N__56783;
    wire N__56776;
    wire N__56771;
    wire N__56768;
    wire N__56765;
    wire N__56758;
    wire N__56743;
    wire N__56740;
    wire N__56737;
    wire N__56734;
    wire N__56731;
    wire N__56728;
    wire N__56727;
    wire N__56726;
    wire N__56723;
    wire N__56720;
    wire N__56719;
    wire N__56716;
    wire N__56711;
    wire N__56708;
    wire N__56707;
    wire N__56704;
    wire N__56703;
    wire N__56700;
    wire N__56697;
    wire N__56694;
    wire N__56691;
    wire N__56688;
    wire N__56685;
    wire N__56682;
    wire N__56671;
    wire N__56668;
    wire N__56665;
    wire N__56662;
    wire N__56659;
    wire N__56656;
    wire N__56653;
    wire N__56652;
    wire N__56651;
    wire N__56650;
    wire N__56647;
    wire N__56646;
    wire N__56643;
    wire N__56642;
    wire N__56637;
    wire N__56634;
    wire N__56631;
    wire N__56630;
    wire N__56629;
    wire N__56626;
    wire N__56623;
    wire N__56620;
    wire N__56617;
    wire N__56614;
    wire N__56611;
    wire N__56608;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56594;
    wire N__56591;
    wire N__56578;
    wire N__56575;
    wire N__56572;
    wire N__56569;
    wire N__56566;
    wire N__56563;
    wire N__56562;
    wire N__56561;
    wire N__56560;
    wire N__56557;
    wire N__56552;
    wire N__56549;
    wire N__56546;
    wire N__56543;
    wire N__56540;
    wire N__56533;
    wire N__56530;
    wire N__56529;
    wire N__56528;
    wire N__56525;
    wire N__56524;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56512;
    wire N__56509;
    wire N__56504;
    wire N__56501;
    wire N__56498;
    wire N__56495;
    wire N__56488;
    wire N__56485;
    wire N__56484;
    wire N__56481;
    wire N__56478;
    wire N__56475;
    wire N__56470;
    wire N__56467;
    wire N__56464;
    wire N__56461;
    wire N__56458;
    wire N__56455;
    wire N__56452;
    wire N__56451;
    wire N__56450;
    wire N__56447;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56437;
    wire N__56434;
    wire N__56429;
    wire N__56426;
    wire N__56421;
    wire N__56418;
    wire N__56413;
    wire N__56410;
    wire N__56409;
    wire N__56406;
    wire N__56403;
    wire N__56400;
    wire N__56399;
    wire N__56398;
    wire N__56393;
    wire N__56390;
    wire N__56387;
    wire N__56384;
    wire N__56379;
    wire N__56378;
    wire N__56373;
    wire N__56370;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56356;
    wire N__56353;
    wire N__56352;
    wire N__56351;
    wire N__56348;
    wire N__56345;
    wire N__56342;
    wire N__56341;
    wire N__56338;
    wire N__56335;
    wire N__56332;
    wire N__56329;
    wire N__56326;
    wire N__56323;
    wire N__56314;
    wire N__56313;
    wire N__56308;
    wire N__56305;
    wire N__56302;
    wire N__56299;
    wire N__56296;
    wire N__56295;
    wire N__56292;
    wire N__56291;
    wire N__56290;
    wire N__56287;
    wire N__56284;
    wire N__56279;
    wire N__56272;
    wire N__56269;
    wire N__56266;
    wire N__56263;
    wire N__56260;
    wire N__56259;
    wire N__56256;
    wire N__56253;
    wire N__56248;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56238;
    wire N__56237;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56226;
    wire N__56225;
    wire N__56224;
    wire N__56221;
    wire N__56214;
    wire N__56213;
    wire N__56210;
    wire N__56207;
    wire N__56204;
    wire N__56201;
    wire N__56200;
    wire N__56197;
    wire N__56194;
    wire N__56193;
    wire N__56188;
    wire N__56185;
    wire N__56182;
    wire N__56179;
    wire N__56176;
    wire N__56173;
    wire N__56170;
    wire N__56167;
    wire N__56164;
    wire N__56161;
    wire N__56158;
    wire N__56155;
    wire N__56154;
    wire N__56149;
    wire N__56146;
    wire N__56143;
    wire N__56140;
    wire N__56135;
    wire N__56132;
    wire N__56127;
    wire N__56126;
    wire N__56123;
    wire N__56120;
    wire N__56117;
    wire N__56114;
    wire N__56111;
    wire N__56108;
    wire N__56103;
    wire N__56098;
    wire N__56093;
    wire N__56086;
    wire N__56085;
    wire N__56084;
    wire N__56081;
    wire N__56080;
    wire N__56077;
    wire N__56074;
    wire N__56071;
    wire N__56068;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56056;
    wire N__56053;
    wire N__56048;
    wire N__56043;
    wire N__56040;
    wire N__56035;
    wire N__56032;
    wire N__56029;
    wire N__56028;
    wire N__56027;
    wire N__56024;
    wire N__56021;
    wire N__56018;
    wire N__56017;
    wire N__56014;
    wire N__56011;
    wire N__56008;
    wire N__56005;
    wire N__56002;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55988;
    wire N__55985;
    wire N__55978;
    wire N__55975;
    wire N__55972;
    wire N__55969;
    wire N__55966;
    wire N__55963;
    wire N__55960;
    wire N__55959;
    wire N__55956;
    wire N__55953;
    wire N__55952;
    wire N__55951;
    wire N__55948;
    wire N__55945;
    wire N__55942;
    wire N__55939;
    wire N__55932;
    wire N__55929;
    wire N__55926;
    wire N__55921;
    wire N__55920;
    wire N__55919;
    wire N__55916;
    wire N__55913;
    wire N__55910;
    wire N__55907;
    wire N__55904;
    wire N__55901;
    wire N__55898;
    wire N__55893;
    wire N__55888;
    wire N__55887;
    wire N__55886;
    wire N__55885;
    wire N__55884;
    wire N__55883;
    wire N__55880;
    wire N__55877;
    wire N__55876;
    wire N__55875;
    wire N__55874;
    wire N__55873;
    wire N__55872;
    wire N__55869;
    wire N__55868;
    wire N__55867;
    wire N__55862;
    wire N__55859;
    wire N__55854;
    wire N__55849;
    wire N__55842;
    wire N__55839;
    wire N__55836;
    wire N__55833;
    wire N__55828;
    wire N__55825;
    wire N__55820;
    wire N__55819;
    wire N__55816;
    wire N__55813;
    wire N__55812;
    wire N__55809;
    wire N__55806;
    wire N__55801;
    wire N__55800;
    wire N__55797;
    wire N__55796;
    wire N__55795;
    wire N__55792;
    wire N__55789;
    wire N__55786;
    wire N__55783;
    wire N__55778;
    wire N__55775;
    wire N__55768;
    wire N__55765;
    wire N__55762;
    wire N__55757;
    wire N__55754;
    wire N__55747;
    wire N__55742;
    wire N__55737;
    wire N__55732;
    wire N__55729;
    wire N__55726;
    wire N__55725;
    wire N__55724;
    wire N__55721;
    wire N__55718;
    wire N__55715;
    wire N__55708;
    wire N__55705;
    wire N__55704;
    wire N__55701;
    wire N__55698;
    wire N__55697;
    wire N__55696;
    wire N__55693;
    wire N__55690;
    wire N__55685;
    wire N__55678;
    wire N__55675;
    wire N__55672;
    wire N__55671;
    wire N__55670;
    wire N__55669;
    wire N__55668;
    wire N__55665;
    wire N__55662;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55642;
    wire N__55639;
    wire N__55636;
    wire N__55631;
    wire N__55628;
    wire N__55623;
    wire N__55618;
    wire N__55615;
    wire N__55614;
    wire N__55611;
    wire N__55610;
    wire N__55607;
    wire N__55604;
    wire N__55601;
    wire N__55598;
    wire N__55593;
    wire N__55588;
    wire N__55587;
    wire N__55586;
    wire N__55585;
    wire N__55584;
    wire N__55583;
    wire N__55580;
    wire N__55575;
    wire N__55572;
    wire N__55569;
    wire N__55566;
    wire N__55559;
    wire N__55556;
    wire N__55549;
    wire N__55548;
    wire N__55545;
    wire N__55544;
    wire N__55541;
    wire N__55540;
    wire N__55537;
    wire N__55532;
    wire N__55529;
    wire N__55526;
    wire N__55523;
    wire N__55516;
    wire N__55515;
    wire N__55512;
    wire N__55511;
    wire N__55510;
    wire N__55509;
    wire N__55506;
    wire N__55505;
    wire N__55502;
    wire N__55499;
    wire N__55496;
    wire N__55493;
    wire N__55490;
    wire N__55487;
    wire N__55484;
    wire N__55477;
    wire N__55468;
    wire N__55467;
    wire N__55466;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55454;
    wire N__55451;
    wire N__55448;
    wire N__55445;
    wire N__55442;
    wire N__55439;
    wire N__55436;
    wire N__55433;
    wire N__55430;
    wire N__55425;
    wire N__55420;
    wire N__55417;
    wire N__55414;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55390;
    wire N__55387;
    wire N__55384;
    wire N__55383;
    wire N__55382;
    wire N__55379;
    wire N__55378;
    wire N__55377;
    wire N__55374;
    wire N__55371;
    wire N__55368;
    wire N__55365;
    wire N__55364;
    wire N__55361;
    wire N__55358;
    wire N__55355;
    wire N__55350;
    wire N__55349;
    wire N__55346;
    wire N__55345;
    wire N__55344;
    wire N__55341;
    wire N__55338;
    wire N__55333;
    wire N__55330;
    wire N__55327;
    wire N__55322;
    wire N__55309;
    wire N__55308;
    wire N__55305;
    wire N__55300;
    wire N__55297;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55285;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55277;
    wire N__55272;
    wire N__55269;
    wire N__55264;
    wire N__55263;
    wire N__55260;
    wire N__55257;
    wire N__55254;
    wire N__55251;
    wire N__55248;
    wire N__55245;
    wire N__55240;
    wire N__55239;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55231;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55219;
    wire N__55214;
    wire N__55213;
    wire N__55212;
    wire N__55209;
    wire N__55206;
    wire N__55203;
    wire N__55200;
    wire N__55197;
    wire N__55186;
    wire N__55185;
    wire N__55184;
    wire N__55183;
    wire N__55182;
    wire N__55181;
    wire N__55180;
    wire N__55179;
    wire N__55178;
    wire N__55175;
    wire N__55172;
    wire N__55169;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55163;
    wire N__55162;
    wire N__55157;
    wire N__55154;
    wire N__55151;
    wire N__55148;
    wire N__55147;
    wire N__55144;
    wire N__55137;
    wire N__55130;
    wire N__55129;
    wire N__55128;
    wire N__55127;
    wire N__55124;
    wire N__55121;
    wire N__55118;
    wire N__55115;
    wire N__55110;
    wire N__55109;
    wire N__55108;
    wire N__55105;
    wire N__55100;
    wire N__55095;
    wire N__55092;
    wire N__55089;
    wire N__55080;
    wire N__55077;
    wire N__55074;
    wire N__55069;
    wire N__55054;
    wire N__55053;
    wire N__55052;
    wire N__55049;
    wire N__55046;
    wire N__55043;
    wire N__55040;
    wire N__55035;
    wire N__55034;
    wire N__55033;
    wire N__55032;
    wire N__55031;
    wire N__55028;
    wire N__55025;
    wire N__55022;
    wire N__55017;
    wire N__55016;
    wire N__55015;
    wire N__55014;
    wire N__55011;
    wire N__55010;
    wire N__55007;
    wire N__55000;
    wire N__54995;
    wire N__54992;
    wire N__54987;
    wire N__54976;
    wire N__54973;
    wire N__54970;
    wire N__54967;
    wire N__54966;
    wire N__54965;
    wire N__54962;
    wire N__54957;
    wire N__54952;
    wire N__54949;
    wire N__54946;
    wire N__54943;
    wire N__54940;
    wire N__54937;
    wire N__54934;
    wire N__54931;
    wire N__54928;
    wire N__54925;
    wire N__54922;
    wire N__54919;
    wire N__54916;
    wire N__54913;
    wire N__54910;
    wire N__54907;
    wire N__54904;
    wire N__54901;
    wire N__54898;
    wire N__54895;
    wire N__54894;
    wire N__54893;
    wire N__54892;
    wire N__54889;
    wire N__54888;
    wire N__54887;
    wire N__54884;
    wire N__54881;
    wire N__54880;
    wire N__54877;
    wire N__54876;
    wire N__54873;
    wire N__54868;
    wire N__54865;
    wire N__54862;
    wire N__54859;
    wire N__54858;
    wire N__54855;
    wire N__54852;
    wire N__54851;
    wire N__54846;
    wire N__54843;
    wire N__54842;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54834;
    wire N__54831;
    wire N__54828;
    wire N__54825;
    wire N__54822;
    wire N__54819;
    wire N__54816;
    wire N__54813;
    wire N__54810;
    wire N__54807;
    wire N__54800;
    wire N__54781;
    wire N__54778;
    wire N__54775;
    wire N__54772;
    wire N__54771;
    wire N__54770;
    wire N__54767;
    wire N__54762;
    wire N__54757;
    wire N__54754;
    wire N__54751;
    wire N__54750;
    wire N__54747;
    wire N__54744;
    wire N__54741;
    wire N__54738;
    wire N__54733;
    wire N__54732;
    wire N__54731;
    wire N__54728;
    wire N__54727;
    wire N__54722;
    wire N__54719;
    wire N__54716;
    wire N__54713;
    wire N__54706;
    wire N__54703;
    wire N__54700;
    wire N__54697;
    wire N__54694;
    wire N__54691;
    wire N__54688;
    wire N__54685;
    wire N__54684;
    wire N__54681;
    wire N__54680;
    wire N__54677;
    wire N__54676;
    wire N__54675;
    wire N__54674;
    wire N__54673;
    wire N__54672;
    wire N__54671;
    wire N__54668;
    wire N__54665;
    wire N__54658;
    wire N__54655;
    wire N__54652;
    wire N__54647;
    wire N__54634;
    wire N__54631;
    wire N__54628;
    wire N__54627;
    wire N__54624;
    wire N__54623;
    wire N__54620;
    wire N__54617;
    wire N__54614;
    wire N__54613;
    wire N__54612;
    wire N__54609;
    wire N__54606;
    wire N__54603;
    wire N__54598;
    wire N__54589;
    wire N__54586;
    wire N__54583;
    wire N__54580;
    wire N__54579;
    wire N__54576;
    wire N__54571;
    wire N__54568;
    wire N__54567;
    wire N__54564;
    wire N__54561;
    wire N__54560;
    wire N__54557;
    wire N__54556;
    wire N__54553;
    wire N__54550;
    wire N__54547;
    wire N__54544;
    wire N__54541;
    wire N__54532;
    wire N__54531;
    wire N__54530;
    wire N__54525;
    wire N__54522;
    wire N__54519;
    wire N__54518;
    wire N__54515;
    wire N__54512;
    wire N__54509;
    wire N__54502;
    wire N__54499;
    wire N__54496;
    wire N__54493;
    wire N__54492;
    wire N__54489;
    wire N__54486;
    wire N__54481;
    wire N__54480;
    wire N__54479;
    wire N__54476;
    wire N__54473;
    wire N__54472;
    wire N__54469;
    wire N__54468;
    wire N__54467;
    wire N__54466;
    wire N__54463;
    wire N__54462;
    wire N__54461;
    wire N__54460;
    wire N__54459;
    wire N__54456;
    wire N__54453;
    wire N__54452;
    wire N__54449;
    wire N__54446;
    wire N__54443;
    wire N__54442;
    wire N__54439;
    wire N__54436;
    wire N__54431;
    wire N__54428;
    wire N__54427;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54421;
    wire N__54418;
    wire N__54415;
    wire N__54412;
    wire N__54411;
    wire N__54410;
    wire N__54405;
    wire N__54402;
    wire N__54399;
    wire N__54396;
    wire N__54395;
    wire N__54388;
    wire N__54385;
    wire N__54384;
    wire N__54383;
    wire N__54378;
    wire N__54373;
    wire N__54370;
    wire N__54365;
    wire N__54360;
    wire N__54351;
    wire N__54348;
    wire N__54343;
    wire N__54340;
    wire N__54337;
    wire N__54316;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54308;
    wire N__54305;
    wire N__54302;
    wire N__54299;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54291;
    wire N__54288;
    wire N__54285;
    wire N__54280;
    wire N__54271;
    wire N__54268;
    wire N__54267;
    wire N__54266;
    wire N__54263;
    wire N__54262;
    wire N__54261;
    wire N__54258;
    wire N__54255;
    wire N__54254;
    wire N__54251;
    wire N__54246;
    wire N__54243;
    wire N__54242;
    wire N__54239;
    wire N__54236;
    wire N__54233;
    wire N__54230;
    wire N__54227;
    wire N__54224;
    wire N__54211;
    wire N__54210;
    wire N__54205;
    wire N__54202;
    wire N__54199;
    wire N__54198;
    wire N__54195;
    wire N__54192;
    wire N__54187;
    wire N__54186;
    wire N__54185;
    wire N__54178;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54166;
    wire N__54163;
    wire N__54162;
    wire N__54159;
    wire N__54156;
    wire N__54155;
    wire N__54152;
    wire N__54149;
    wire N__54146;
    wire N__54143;
    wire N__54136;
    wire N__54135;
    wire N__54134;
    wire N__54131;
    wire N__54130;
    wire N__54127;
    wire N__54126;
    wire N__54123;
    wire N__54122;
    wire N__54119;
    wire N__54116;
    wire N__54115;
    wire N__54112;
    wire N__54109;
    wire N__54106;
    wire N__54103;
    wire N__54098;
    wire N__54097;
    wire N__54096;
    wire N__54095;
    wire N__54094;
    wire N__54091;
    wire N__54088;
    wire N__54079;
    wire N__54070;
    wire N__54067;
    wire N__54058;
    wire N__54055;
    wire N__54054;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54042;
    wire N__54039;
    wire N__54036;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54022;
    wire N__54021;
    wire N__54020;
    wire N__54017;
    wire N__54014;
    wire N__54011;
    wire N__54008;
    wire N__54005;
    wire N__54002;
    wire N__53999;
    wire N__53996;
    wire N__53993;
    wire N__53986;
    wire N__53983;
    wire N__53980;
    wire N__53977;
    wire N__53974;
    wire N__53973;
    wire N__53970;
    wire N__53967;
    wire N__53964;
    wire N__53963;
    wire N__53960;
    wire N__53957;
    wire N__53954;
    wire N__53947;
    wire N__53944;
    wire N__53943;
    wire N__53942;
    wire N__53939;
    wire N__53936;
    wire N__53933;
    wire N__53930;
    wire N__53927;
    wire N__53924;
    wire N__53921;
    wire N__53918;
    wire N__53911;
    wire N__53908;
    wire N__53907;
    wire N__53904;
    wire N__53901;
    wire N__53898;
    wire N__53895;
    wire N__53892;
    wire N__53889;
    wire N__53884;
    wire N__53881;
    wire N__53878;
    wire N__53875;
    wire N__53874;
    wire N__53871;
    wire N__53870;
    wire N__53869;
    wire N__53868;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53854;
    wire N__53851;
    wire N__53842;
    wire N__53839;
    wire N__53838;
    wire N__53837;
    wire N__53834;
    wire N__53829;
    wire N__53824;
    wire N__53821;
    wire N__53818;
    wire N__53815;
    wire N__53812;
    wire N__53809;
    wire N__53808;
    wire N__53805;
    wire N__53804;
    wire N__53801;
    wire N__53798;
    wire N__53795;
    wire N__53794;
    wire N__53791;
    wire N__53786;
    wire N__53783;
    wire N__53780;
    wire N__53777;
    wire N__53770;
    wire N__53769;
    wire N__53768;
    wire N__53765;
    wire N__53760;
    wire N__53755;
    wire N__53752;
    wire N__53751;
    wire N__53748;
    wire N__53745;
    wire N__53744;
    wire N__53741;
    wire N__53738;
    wire N__53735;
    wire N__53732;
    wire N__53729;
    wire N__53722;
    wire N__53721;
    wire N__53720;
    wire N__53715;
    wire N__53714;
    wire N__53711;
    wire N__53710;
    wire N__53709;
    wire N__53706;
    wire N__53703;
    wire N__53702;
    wire N__53699;
    wire N__53694;
    wire N__53693;
    wire N__53688;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53676;
    wire N__53671;
    wire N__53662;
    wire N__53659;
    wire N__53658;
    wire N__53657;
    wire N__53654;
    wire N__53651;
    wire N__53648;
    wire N__53645;
    wire N__53642;
    wire N__53639;
    wire N__53636;
    wire N__53633;
    wire N__53626;
    wire N__53623;
    wire N__53622;
    wire N__53619;
    wire N__53618;
    wire N__53615;
    wire N__53612;
    wire N__53609;
    wire N__53602;
    wire N__53601;
    wire N__53598;
    wire N__53595;
    wire N__53592;
    wire N__53587;
    wire N__53586;
    wire N__53585;
    wire N__53582;
    wire N__53579;
    wire N__53576;
    wire N__53573;
    wire N__53570;
    wire N__53563;
    wire N__53560;
    wire N__53557;
    wire N__53556;
    wire N__53553;
    wire N__53550;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53538;
    wire N__53537;
    wire N__53532;
    wire N__53529;
    wire N__53526;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53512;
    wire N__53511;
    wire N__53510;
    wire N__53507;
    wire N__53506;
    wire N__53501;
    wire N__53498;
    wire N__53495;
    wire N__53494;
    wire N__53491;
    wire N__53488;
    wire N__53485;
    wire N__53482;
    wire N__53473;
    wire N__53470;
    wire N__53469;
    wire N__53466;
    wire N__53463;
    wire N__53460;
    wire N__53459;
    wire N__53456;
    wire N__53453;
    wire N__53450;
    wire N__53443;
    wire N__53442;
    wire N__53439;
    wire N__53436;
    wire N__53433;
    wire N__53430;
    wire N__53425;
    wire N__53422;
    wire N__53421;
    wire N__53418;
    wire N__53415;
    wire N__53414;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53400;
    wire N__53395;
    wire N__53392;
    wire N__53391;
    wire N__53386;
    wire N__53383;
    wire N__53380;
    wire N__53379;
    wire N__53376;
    wire N__53375;
    wire N__53372;
    wire N__53369;
    wire N__53366;
    wire N__53363;
    wire N__53358;
    wire N__53353;
    wire N__53350;
    wire N__53347;
    wire N__53344;
    wire N__53343;
    wire N__53342;
    wire N__53339;
    wire N__53334;
    wire N__53333;
    wire N__53330;
    wire N__53327;
    wire N__53326;
    wire N__53325;
    wire N__53322;
    wire N__53319;
    wire N__53316;
    wire N__53311;
    wire N__53302;
    wire N__53299;
    wire N__53298;
    wire N__53297;
    wire N__53294;
    wire N__53289;
    wire N__53284;
    wire N__53281;
    wire N__53280;
    wire N__53275;
    wire N__53272;
    wire N__53271;
    wire N__53266;
    wire N__53263;
    wire N__53260;
    wire N__53259;
    wire N__53256;
    wire N__53255;
    wire N__53252;
    wire N__53249;
    wire N__53246;
    wire N__53243;
    wire N__53238;
    wire N__53235;
    wire N__53230;
    wire N__53229;
    wire N__53228;
    wire N__53227;
    wire N__53226;
    wire N__53225;
    wire N__53224;
    wire N__53223;
    wire N__53222;
    wire N__53221;
    wire N__53220;
    wire N__53219;
    wire N__53218;
    wire N__53217;
    wire N__53216;
    wire N__53215;
    wire N__53212;
    wire N__53211;
    wire N__53210;
    wire N__53209;
    wire N__53208;
    wire N__53205;
    wire N__53202;
    wire N__53199;
    wire N__53196;
    wire N__53195;
    wire N__53192;
    wire N__53189;
    wire N__53188;
    wire N__53187;
    wire N__53180;
    wire N__53179;
    wire N__53178;
    wire N__53177;
    wire N__53176;
    wire N__53175;
    wire N__53174;
    wire N__53173;
    wire N__53172;
    wire N__53165;
    wire N__53160;
    wire N__53157;
    wire N__53154;
    wire N__53145;
    wire N__53136;
    wire N__53135;
    wire N__53132;
    wire N__53129;
    wire N__53122;
    wire N__53119;
    wire N__53118;
    wire N__53115;
    wire N__53112;
    wire N__53109;
    wire N__53106;
    wire N__53103;
    wire N__53100;
    wire N__53095;
    wire N__53092;
    wire N__53087;
    wire N__53080;
    wire N__53079;
    wire N__53076;
    wire N__53071;
    wire N__53066;
    wire N__53063;
    wire N__53060;
    wire N__53055;
    wire N__53040;
    wire N__53037;
    wire N__53036;
    wire N__53033;
    wire N__53030;
    wire N__53027;
    wire N__53024;
    wire N__53015;
    wire N__53012;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53000;
    wire N__52997;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52978;
    wire N__52975;
    wire N__52960;
    wire N__52957;
    wire N__52956;
    wire N__52953;
    wire N__52950;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52942;
    wire N__52939;
    wire N__52936;
    wire N__52933;
    wire N__52930;
    wire N__52921;
    wire N__52920;
    wire N__52919;
    wire N__52916;
    wire N__52913;
    wire N__52910;
    wire N__52907;
    wire N__52904;
    wire N__52903;
    wire N__52900;
    wire N__52895;
    wire N__52892;
    wire N__52889;
    wire N__52886;
    wire N__52879;
    wire N__52876;
    wire N__52875;
    wire N__52872;
    wire N__52869;
    wire N__52864;
    wire N__52863;
    wire N__52862;
    wire N__52859;
    wire N__52854;
    wire N__52849;
    wire N__52846;
    wire N__52843;
    wire N__52840;
    wire N__52837;
    wire N__52834;
    wire N__52831;
    wire N__52828;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52818;
    wire N__52815;
    wire N__52812;
    wire N__52809;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52774;
    wire N__52771;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52759;
    wire N__52758;
    wire N__52755;
    wire N__52752;
    wire N__52749;
    wire N__52746;
    wire N__52743;
    wire N__52740;
    wire N__52735;
    wire N__52734;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52722;
    wire N__52719;
    wire N__52716;
    wire N__52711;
    wire N__52708;
    wire N__52707;
    wire N__52706;
    wire N__52703;
    wire N__52698;
    wire N__52693;
    wire N__52690;
    wire N__52689;
    wire N__52686;
    wire N__52683;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52671;
    wire N__52668;
    wire N__52665;
    wire N__52662;
    wire N__52657;
    wire N__52654;
    wire N__52651;
    wire N__52648;
    wire N__52647;
    wire N__52646;
    wire N__52645;
    wire N__52642;
    wire N__52637;
    wire N__52634;
    wire N__52629;
    wire N__52626;
    wire N__52623;
    wire N__52620;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52579;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52567;
    wire N__52564;
    wire N__52563;
    wire N__52560;
    wire N__52559;
    wire N__52556;
    wire N__52553;
    wire N__52550;
    wire N__52547;
    wire N__52544;
    wire N__52543;
    wire N__52540;
    wire N__52535;
    wire N__52532;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52510;
    wire N__52507;
    wire N__52506;
    wire N__52505;
    wire N__52500;
    wire N__52497;
    wire N__52492;
    wire N__52491;
    wire N__52490;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52482;
    wire N__52479;
    wire N__52476;
    wire N__52473;
    wire N__52470;
    wire N__52467;
    wire N__52462;
    wire N__52459;
    wire N__52454;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52435;
    wire N__52432;
    wire N__52423;
    wire N__52420;
    wire N__52417;
    wire N__52416;
    wire N__52413;
    wire N__52410;
    wire N__52405;
    wire N__52402;
    wire N__52399;
    wire N__52398;
    wire N__52397;
    wire N__52394;
    wire N__52391;
    wire N__52388;
    wire N__52385;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52351;
    wire N__52350;
    wire N__52347;
    wire N__52346;
    wire N__52345;
    wire N__52342;
    wire N__52339;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52331;
    wire N__52328;
    wire N__52325;
    wire N__52322;
    wire N__52319;
    wire N__52316;
    wire N__52313;
    wire N__52308;
    wire N__52305;
    wire N__52300;
    wire N__52297;
    wire N__52294;
    wire N__52289;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52275;
    wire N__52272;
    wire N__52269;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52210;
    wire N__52207;
    wire N__52206;
    wire N__52203;
    wire N__52200;
    wire N__52195;
    wire N__52192;
    wire N__52189;
    wire N__52186;
    wire N__52185;
    wire N__52184;
    wire N__52181;
    wire N__52176;
    wire N__52171;
    wire N__52168;
    wire N__52167;
    wire N__52166;
    wire N__52163;
    wire N__52160;
    wire N__52159;
    wire N__52158;
    wire N__52155;
    wire N__52152;
    wire N__52149;
    wire N__52144;
    wire N__52135;
    wire N__52134;
    wire N__52131;
    wire N__52130;
    wire N__52127;
    wire N__52124;
    wire N__52121;
    wire N__52118;
    wire N__52115;
    wire N__52108;
    wire N__52107;
    wire N__52104;
    wire N__52103;
    wire N__52100;
    wire N__52097;
    wire N__52094;
    wire N__52093;
    wire N__52092;
    wire N__52089;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52070;
    wire N__52067;
    wire N__52060;
    wire N__52057;
    wire N__52054;
    wire N__52053;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52041;
    wire N__52040;
    wire N__52037;
    wire N__52034;
    wire N__52031;
    wire N__52024;
    wire N__52021;
    wire N__52020;
    wire N__52019;
    wire N__52016;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51997;
    wire N__51992;
    wire N__51991;
    wire N__51986;
    wire N__51983;
    wire N__51980;
    wire N__51973;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51951;
    wire N__51946;
    wire N__51943;
    wire N__51942;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51927;
    wire N__51924;
    wire N__51919;
    wire N__51916;
    wire N__51913;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51903;
    wire N__51900;
    wire N__51895;
    wire N__51892;
    wire N__51889;
    wire N__51886;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51846;
    wire N__51843;
    wire N__51840;
    wire N__51837;
    wire N__51834;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51824;
    wire N__51821;
    wire N__51818;
    wire N__51811;
    wire N__51808;
    wire N__51807;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51792;
    wire N__51787;
    wire N__51786;
    wire N__51785;
    wire N__51782;
    wire N__51777;
    wire N__51776;
    wire N__51775;
    wire N__51770;
    wire N__51765;
    wire N__51760;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51744;
    wire N__51741;
    wire N__51736;
    wire N__51733;
    wire N__51730;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51718;
    wire N__51715;
    wire N__51712;
    wire N__51711;
    wire N__51708;
    wire N__51707;
    wire N__51706;
    wire N__51703;
    wire N__51700;
    wire N__51695;
    wire N__51688;
    wire N__51687;
    wire N__51686;
    wire N__51685;
    wire N__51682;
    wire N__51675;
    wire N__51674;
    wire N__51673;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51658;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51627;
    wire N__51624;
    wire N__51623;
    wire N__51618;
    wire N__51617;
    wire N__51614;
    wire N__51611;
    wire N__51608;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51588;
    wire N__51583;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51573;
    wire N__51570;
    wire N__51567;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51541;
    wire N__51540;
    wire N__51539;
    wire N__51538;
    wire N__51535;
    wire N__51532;
    wire N__51527;
    wire N__51520;
    wire N__51519;
    wire N__51518;
    wire N__51515;
    wire N__51514;
    wire N__51513;
    wire N__51510;
    wire N__51507;
    wire N__51504;
    wire N__51501;
    wire N__51498;
    wire N__51495;
    wire N__51492;
    wire N__51489;
    wire N__51484;
    wire N__51479;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51457;
    wire N__51456;
    wire N__51453;
    wire N__51450;
    wire N__51445;
    wire N__51442;
    wire N__51439;
    wire N__51436;
    wire N__51433;
    wire N__51432;
    wire N__51429;
    wire N__51426;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51414;
    wire N__51411;
    wire N__51410;
    wire N__51407;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51349;
    wire N__51346;
    wire N__51345;
    wire N__51342;
    wire N__51339;
    wire N__51338;
    wire N__51335;
    wire N__51332;
    wire N__51331;
    wire N__51330;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51312;
    wire N__51301;
    wire N__51298;
    wire N__51295;
    wire N__51292;
    wire N__51291;
    wire N__51288;
    wire N__51287;
    wire N__51284;
    wire N__51283;
    wire N__51282;
    wire N__51279;
    wire N__51276;
    wire N__51273;
    wire N__51270;
    wire N__51267;
    wire N__51266;
    wire N__51261;
    wire N__51260;
    wire N__51259;
    wire N__51258;
    wire N__51257;
    wire N__51256;
    wire N__51255;
    wire N__51252;
    wire N__51249;
    wire N__51244;
    wire N__51241;
    wire N__51234;
    wire N__51227;
    wire N__51214;
    wire N__51211;
    wire N__51208;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51171;
    wire N__51168;
    wire N__51165;
    wire N__51162;
    wire N__51157;
    wire N__51154;
    wire N__51153;
    wire N__51150;
    wire N__51147;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51114;
    wire N__51109;
    wire N__51108;
    wire N__51105;
    wire N__51104;
    wire N__51101;
    wire N__51098;
    wire N__51097;
    wire N__51094;
    wire N__51091;
    wire N__51090;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51078;
    wire N__51075;
    wire N__51070;
    wire N__51061;
    wire N__51058;
    wire N__51055;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51043;
    wire N__51040;
    wire N__51037;
    wire N__51034;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51015;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50997;
    wire N__50992;
    wire N__50989;
    wire N__50988;
    wire N__50985;
    wire N__50984;
    wire N__50981;
    wire N__50978;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50968;
    wire N__50965;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50953;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50937;
    wire N__50934;
    wire N__50933;
    wire N__50930;
    wire N__50927;
    wire N__50924;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50908;
    wire N__50905;
    wire N__50904;
    wire N__50903;
    wire N__50900;
    wire N__50897;
    wire N__50894;
    wire N__50891;
    wire N__50888;
    wire N__50885;
    wire N__50882;
    wire N__50879;
    wire N__50872;
    wire N__50869;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50853;
    wire N__50852;
    wire N__50849;
    wire N__50844;
    wire N__50839;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50797;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50785;
    wire N__50784;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50763;
    wire N__50760;
    wire N__50757;
    wire N__50754;
    wire N__50749;
    wire N__50746;
    wire N__50743;
    wire N__50740;
    wire N__50739;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50722;
    wire N__50719;
    wire N__50716;
    wire N__50713;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50695;
    wire N__50692;
    wire N__50691;
    wire N__50688;
    wire N__50685;
    wire N__50680;
    wire N__50679;
    wire N__50678;
    wire N__50675;
    wire N__50674;
    wire N__50673;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50659;
    wire N__50654;
    wire N__50651;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50641;
    wire N__50640;
    wire N__50639;
    wire N__50636;
    wire N__50633;
    wire N__50624;
    wire N__50621;
    wire N__50616;
    wire N__50605;
    wire N__50604;
    wire N__50603;
    wire N__50602;
    wire N__50601;
    wire N__50600;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50583;
    wire N__50582;
    wire N__50579;
    wire N__50576;
    wire N__50573;
    wire N__50570;
    wire N__50567;
    wire N__50566;
    wire N__50563;
    wire N__50558;
    wire N__50555;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50551;
    wire N__50550;
    wire N__50545;
    wire N__50538;
    wire N__50535;
    wire N__50530;
    wire N__50525;
    wire N__50518;
    wire N__50515;
    wire N__50500;
    wire N__50497;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50486;
    wire N__50485;
    wire N__50482;
    wire N__50479;
    wire N__50474;
    wire N__50467;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50457;
    wire N__50456;
    wire N__50453;
    wire N__50450;
    wire N__50447;
    wire N__50442;
    wire N__50439;
    wire N__50434;
    wire N__50433;
    wire N__50432;
    wire N__50429;
    wire N__50426;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50412;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50379;
    wire N__50376;
    wire N__50371;
    wire N__50362;
    wire N__50361;
    wire N__50360;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50350;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50346;
    wire N__50343;
    wire N__50340;
    wire N__50339;
    wire N__50336;
    wire N__50333;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50321;
    wire N__50318;
    wire N__50317;
    wire N__50314;
    wire N__50313;
    wire N__50310;
    wire N__50305;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50297;
    wire N__50290;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50282;
    wire N__50279;
    wire N__50272;
    wire N__50267;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50226;
    wire N__50223;
    wire N__50220;
    wire N__50217;
    wire N__50214;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50150;
    wire N__50149;
    wire N__50146;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50129;
    wire N__50126;
    wire N__50123;
    wire N__50120;
    wire N__50113;
    wire N__50110;
    wire N__50109;
    wire N__50108;
    wire N__50105;
    wire N__50102;
    wire N__50099;
    wire N__50092;
    wire N__50089;
    wire N__50086;
    wire N__50083;
    wire N__50082;
    wire N__50081;
    wire N__50078;
    wire N__50077;
    wire N__50076;
    wire N__50073;
    wire N__50070;
    wire N__50067;
    wire N__50064;
    wire N__50063;
    wire N__50060;
    wire N__50057;
    wire N__50054;
    wire N__50049;
    wire N__50046;
    wire N__50043;
    wire N__50038;
    wire N__50033;
    wire N__50026;
    wire N__50023;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50005;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49995;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49976;
    wire N__49975;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49965;
    wire N__49960;
    wire N__49951;
    wire N__49948;
    wire N__49945;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49927;
    wire N__49924;
    wire N__49921;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49907;
    wire N__49906;
    wire N__49903;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49886;
    wire N__49879;
    wire N__49876;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49858;
    wire N__49855;
    wire N__49852;
    wire N__49851;
    wire N__49848;
    wire N__49847;
    wire N__49844;
    wire N__49841;
    wire N__49838;
    wire N__49835;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49816;
    wire N__49813;
    wire N__49810;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49802;
    wire N__49799;
    wire N__49794;
    wire N__49789;
    wire N__49786;
    wire N__49785;
    wire N__49782;
    wire N__49781;
    wire N__49778;
    wire N__49775;
    wire N__49770;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49751;
    wire N__49748;
    wire N__49745;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49734;
    wire N__49731;
    wire N__49730;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49706;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49688;
    wire N__49683;
    wire N__49678;
    wire N__49677;
    wire N__49676;
    wire N__49673;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49665;
    wire N__49662;
    wire N__49659;
    wire N__49656;
    wire N__49655;
    wire N__49652;
    wire N__49649;
    wire N__49644;
    wire N__49641;
    wire N__49638;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49619;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49606;
    wire N__49597;
    wire N__49594;
    wire N__49591;
    wire N__49588;
    wire N__49585;
    wire N__49582;
    wire N__49581;
    wire N__49578;
    wire N__49577;
    wire N__49574;
    wire N__49571;
    wire N__49566;
    wire N__49563;
    wire N__49560;
    wire N__49559;
    wire N__49558;
    wire N__49553;
    wire N__49548;
    wire N__49543;
    wire N__49540;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49532;
    wire N__49527;
    wire N__49522;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49510;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49502;
    wire N__49499;
    wire N__49498;
    wire N__49495;
    wire N__49492;
    wire N__49491;
    wire N__49488;
    wire N__49487;
    wire N__49484;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49459;
    wire N__49458;
    wire N__49455;
    wire N__49454;
    wire N__49451;
    wire N__49448;
    wire N__49445;
    wire N__49444;
    wire N__49441;
    wire N__49436;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49423;
    wire N__49414;
    wire N__49411;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49401;
    wire N__49398;
    wire N__49397;
    wire N__49396;
    wire N__49393;
    wire N__49390;
    wire N__49387;
    wire N__49384;
    wire N__49375;
    wire N__49372;
    wire N__49371;
    wire N__49368;
    wire N__49365;
    wire N__49362;
    wire N__49357;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49347;
    wire N__49346;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49334;
    wire N__49329;
    wire N__49328;
    wire N__49327;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49312;
    wire N__49303;
    wire N__49302;
    wire N__49301;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49269;
    wire N__49266;
    wire N__49261;
    wire N__49260;
    wire N__49259;
    wire N__49258;
    wire N__49257;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49231;
    wire N__49230;
    wire N__49229;
    wire N__49228;
    wire N__49227;
    wire N__49222;
    wire N__49219;
    wire N__49214;
    wire N__49213;
    wire N__49210;
    wire N__49205;
    wire N__49202;
    wire N__49199;
    wire N__49196;
    wire N__49193;
    wire N__49188;
    wire N__49183;
    wire N__49182;
    wire N__49179;
    wire N__49178;
    wire N__49175;
    wire N__49172;
    wire N__49169;
    wire N__49166;
    wire N__49161;
    wire N__49160;
    wire N__49155;
    wire N__49152;
    wire N__49147;
    wire N__49144;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49124;
    wire N__49121;
    wire N__49118;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49098;
    wire N__49095;
    wire N__49092;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49076;
    wire N__49073;
    wire N__49070;
    wire N__49069;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49045;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49031;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49017;
    wire N__49014;
    wire N__49011;
    wire N__49006;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48960;
    wire N__48957;
    wire N__48954;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48933;
    wire N__48932;
    wire N__48931;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48921;
    wire N__48916;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48880;
    wire N__48877;
    wire N__48876;
    wire N__48873;
    wire N__48870;
    wire N__48869;
    wire N__48864;
    wire N__48861;
    wire N__48860;
    wire N__48855;
    wire N__48852;
    wire N__48849;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48837;
    wire N__48834;
    wire N__48831;
    wire N__48830;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48790;
    wire N__48789;
    wire N__48786;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48778;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48743;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48721;
    wire N__48716;
    wire N__48711;
    wire N__48708;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48666;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48654;
    wire N__48651;
    wire N__48650;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48618;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48605;
    wire N__48602;
    wire N__48599;
    wire N__48596;
    wire N__48595;
    wire N__48592;
    wire N__48587;
    wire N__48584;
    wire N__48581;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48534;
    wire N__48531;
    wire N__48528;
    wire N__48527;
    wire N__48524;
    wire N__48521;
    wire N__48518;
    wire N__48511;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48441;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48381;
    wire N__48378;
    wire N__48377;
    wire N__48374;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48366;
    wire N__48363;
    wire N__48360;
    wire N__48355;
    wire N__48352;
    wire N__48345;
    wire N__48342;
    wire N__48339;
    wire N__48334;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48314;
    wire N__48311;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48265;
    wire N__48262;
    wire N__48261;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48243;
    wire N__48240;
    wire N__48237;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48225;
    wire N__48220;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48192;
    wire N__48187;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48177;
    wire N__48174;
    wire N__48171;
    wire N__48168;
    wire N__48163;
    wire N__48162;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48127;
    wire N__48120;
    wire N__48117;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48103;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48085;
    wire N__48082;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48068;
    wire N__48065;
    wire N__48062;
    wire N__48059;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48033;
    wire N__48032;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48012;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47977;
    wire N__47976;
    wire N__47975;
    wire N__47972;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47944;
    wire N__47941;
    wire N__47938;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47925;
    wire N__47922;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47911;
    wire N__47908;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47850;
    wire N__47845;
    wire N__47842;
    wire N__47839;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47831;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47799;
    wire N__47794;
    wire N__47789;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47772;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47734;
    wire N__47731;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47689;
    wire N__47688;
    wire N__47685;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47670;
    wire N__47667;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47646;
    wire N__47643;
    wire N__47640;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47623;
    wire N__47620;
    wire N__47619;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47599;
    wire N__47598;
    wire N__47597;
    wire N__47596;
    wire N__47593;
    wire N__47588;
    wire N__47585;
    wire N__47582;
    wire N__47577;
    wire N__47572;
    wire N__47569;
    wire N__47560;
    wire N__47559;
    wire N__47556;
    wire N__47555;
    wire N__47552;
    wire N__47549;
    wire N__47548;
    wire N__47547;
    wire N__47546;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47531;
    wire N__47526;
    wire N__47521;
    wire N__47512;
    wire N__47509;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47491;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47479;
    wire N__47476;
    wire N__47473;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47374;
    wire N__47371;
    wire N__47370;
    wire N__47369;
    wire N__47366;
    wire N__47361;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47340;
    wire N__47337;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47322;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47298;
    wire N__47297;
    wire N__47296;
    wire N__47289;
    wire N__47286;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47274;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47259;
    wire N__47256;
    wire N__47255;
    wire N__47252;
    wire N__47247;
    wire N__47244;
    wire N__47239;
    wire N__47236;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47217;
    wire N__47216;
    wire N__47213;
    wire N__47210;
    wire N__47207;
    wire N__47206;
    wire N__47205;
    wire N__47200;
    wire N__47197;
    wire N__47192;
    wire N__47189;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47161;
    wire N__47158;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47145;
    wire N__47142;
    wire N__47139;
    wire N__47136;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47082;
    wire N__47079;
    wire N__47076;
    wire N__47071;
    wire N__47068;
    wire N__47065;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47034;
    wire N__47033;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47021;
    wire N__47014;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46993;
    wire N__46992;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46881;
    wire N__46878;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46864;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46848;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46830;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46821;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46803;
    wire N__46800;
    wire N__46799;
    wire N__46798;
    wire N__46797;
    wire N__46796;
    wire N__46795;
    wire N__46788;
    wire N__46781;
    wire N__46780;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46761;
    wire N__46756;
    wire N__46749;
    wire N__46744;
    wire N__46739;
    wire N__46738;
    wire N__46737;
    wire N__46736;
    wire N__46735;
    wire N__46734;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46730;
    wire N__46729;
    wire N__46728;
    wire N__46727;
    wire N__46726;
    wire N__46725;
    wire N__46724;
    wire N__46723;
    wire N__46714;
    wire N__46709;
    wire N__46704;
    wire N__46699;
    wire N__46696;
    wire N__46693;
    wire N__46692;
    wire N__46691;
    wire N__46688;
    wire N__46683;
    wire N__46678;
    wire N__46673;
    wire N__46668;
    wire N__46665;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46651;
    wire N__46650;
    wire N__46649;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46636;
    wire N__46627;
    wire N__46624;
    wire N__46623;
    wire N__46622;
    wire N__46619;
    wire N__46610;
    wire N__46603;
    wire N__46600;
    wire N__46593;
    wire N__46588;
    wire N__46585;
    wire N__46582;
    wire N__46577;
    wire N__46572;
    wire N__46569;
    wire N__46564;
    wire N__46549;
    wire N__46542;
    wire N__46531;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46513;
    wire N__46510;
    wire N__46505;
    wire N__46498;
    wire N__46495;
    wire N__46490;
    wire N__46485;
    wire N__46478;
    wire N__46473;
    wire N__46468;
    wire N__46463;
    wire N__46458;
    wire N__46455;
    wire N__46450;
    wire N__46443;
    wire N__46438;
    wire N__46431;
    wire N__46420;
    wire N__46417;
    wire N__46416;
    wire N__46415;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46393;
    wire N__46392;
    wire N__46391;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46369;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46334;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46303;
    wire N__46302;
    wire N__46301;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46288;
    wire N__46287;
    wire N__46284;
    wire N__46283;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46273;
    wire N__46270;
    wire N__46269;
    wire N__46266;
    wire N__46265;
    wire N__46262;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46230;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46153;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46139;
    wire N__46138;
    wire N__46137;
    wire N__46136;
    wire N__46135;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46116;
    wire N__46113;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46095;
    wire N__46094;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46053;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46035;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46003;
    wire N__46000;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45955;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45937;
    wire N__45936;
    wire N__45935;
    wire N__45932;
    wire N__45931;
    wire N__45930;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45876;
    wire N__45871;
    wire N__45870;
    wire N__45869;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45836;
    wire N__45829;
    wire N__45826;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45814;
    wire N__45811;
    wire N__45810;
    wire N__45805;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45766;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45748;
    wire N__45745;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45713;
    wire N__45710;
    wire N__45705;
    wire N__45704;
    wire N__45703;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45680;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45639;
    wire N__45638;
    wire N__45637;
    wire N__45634;
    wire N__45633;
    wire N__45630;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45613;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45586;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45564;
    wire N__45561;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45546;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45510;
    wire N__45509;
    wire N__45506;
    wire N__45501;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45453;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45422;
    wire N__45417;
    wire N__45412;
    wire N__45409;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45394;
    wire N__45391;
    wire N__45390;
    wire N__45385;
    wire N__45382;
    wire N__45379;
    wire N__45376;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45366;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45345;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45335;
    wire N__45334;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45316;
    wire N__45315;
    wire N__45310;
    wire N__45307;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45274;
    wire N__45271;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45189;
    wire N__45188;
    wire N__45183;
    wire N__45182;
    wire N__45181;
    wire N__45180;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45163;
    wire N__45154;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45141;
    wire N__45138;
    wire N__45137;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45107;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45070;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45052;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45038;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45022;
    wire N__45021;
    wire N__45020;
    wire N__45017;
    wire N__45016;
    wire N__45015;
    wire N__45014;
    wire N__45009;
    wire N__45006;
    wire N__44999;
    wire N__44996;
    wire N__44991;
    wire N__44986;
    wire N__44985;
    wire N__44980;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44969;
    wire N__44964;
    wire N__44957;
    wire N__44954;
    wire N__44947;
    wire N__44946;
    wire N__44945;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44929;
    wire N__44920;
    wire N__44917;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44897;
    wire N__44894;
    wire N__44893;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44860;
    wire N__44855;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44805;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44731;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44716;
    wire N__44713;
    wire N__44712;
    wire N__44707;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44676;
    wire N__44671;
    wire N__44668;
    wire N__44665;
    wire N__44662;
    wire N__44659;
    wire N__44658;
    wire N__44655;
    wire N__44654;
    wire N__44651;
    wire N__44646;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44634;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44624;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44602;
    wire N__44597;
    wire N__44594;
    wire N__44589;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44559;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44481;
    wire N__44480;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44424;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44413;
    wire N__44410;
    wire N__44403;
    wire N__44398;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44383;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44368;
    wire N__44359;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44328;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44310;
    wire N__44305;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44293;
    wire N__44292;
    wire N__44287;
    wire N__44284;
    wire N__44281;
    wire N__44280;
    wire N__44275;
    wire N__44272;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44253;
    wire N__44252;
    wire N__44249;
    wire N__44248;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44220;
    wire N__44217;
    wire N__44216;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44188;
    wire N__44185;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44158;
    wire N__44157;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44151;
    wire N__44148;
    wire N__44143;
    wire N__44140;
    wire N__44137;
    wire N__44128;
    wire N__44127;
    wire N__44126;
    wire N__44125;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44119;
    wire N__44118;
    wire N__44117;
    wire N__44114;
    wire N__44109;
    wire N__44102;
    wire N__44099;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44058;
    wire N__44053;
    wire N__44050;
    wire N__44049;
    wire N__44048;
    wire N__44047;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44031;
    wire N__44030;
    wire N__44029;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44014;
    wire N__44005;
    wire N__44002;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43974;
    wire N__43973;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43961;
    wire N__43954;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43942;
    wire N__43941;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43924;
    wire N__43923;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43908;
    wire N__43907;
    wire N__43906;
    wire N__43903;
    wire N__43898;
    wire N__43895;
    wire N__43888;
    wire N__43887;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43877;
    wire N__43870;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43849;
    wire N__43846;
    wire N__43841;
    wire N__43840;
    wire N__43839;
    wire N__43836;
    wire N__43831;
    wire N__43826;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43802;
    wire N__43801;
    wire N__43800;
    wire N__43799;
    wire N__43794;
    wire N__43791;
    wire N__43790;
    wire N__43783;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43744;
    wire N__43743;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43695;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43677;
    wire N__43674;
    wire N__43669;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43618;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43521;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43506;
    wire N__43503;
    wire N__43498;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43455;
    wire N__43454;
    wire N__43451;
    wire N__43446;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43420;
    wire N__43419;
    wire N__43416;
    wire N__43411;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43389;
    wire N__43386;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43282;
    wire N__43279;
    wire N__43278;
    wire N__43277;
    wire N__43276;
    wire N__43275;
    wire N__43274;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43262;
    wire N__43257;
    wire N__43254;
    wire N__43247;
    wire N__43240;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43089;
    wire N__43088;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43070;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43034;
    wire N__43027;
    wire N__43024;
    wire N__43023;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42969;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42909;
    wire N__42904;
    wire N__42901;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42792;
    wire N__42787;
    wire N__42784;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42717;
    wire N__42714;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42676;
    wire N__42673;
    wire N__42672;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42662;
    wire N__42659;
    wire N__42654;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42632;
    wire N__42629;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42599;
    wire N__42594;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42576;
    wire N__42575;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42555;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42541;
    wire N__42540;
    wire N__42537;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42527;
    wire N__42520;
    wire N__42519;
    wire N__42518;
    wire N__42517;
    wire N__42516;
    wire N__42513;
    wire N__42512;
    wire N__42509;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42505;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42497;
    wire N__42496;
    wire N__42495;
    wire N__42488;
    wire N__42483;
    wire N__42480;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42448;
    wire N__42443;
    wire N__42438;
    wire N__42435;
    wire N__42430;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42426;
    wire N__42423;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42403;
    wire N__42400;
    wire N__42393;
    wire N__42390;
    wire N__42385;
    wire N__42370;
    wire N__42369;
    wire N__42368;
    wire N__42365;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42343;
    wire N__42338;
    wire N__42331;
    wire N__42330;
    wire N__42329;
    wire N__42328;
    wire N__42325;
    wire N__42324;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42310;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42294;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42280;
    wire N__42277;
    wire N__42268;
    wire N__42267;
    wire N__42266;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42251;
    wire N__42250;
    wire N__42249;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42227;
    wire N__42226;
    wire N__42225;
    wire N__42224;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42204;
    wire N__42201;
    wire N__42200;
    wire N__42199;
    wire N__42198;
    wire N__42197;
    wire N__42196;
    wire N__42195;
    wire N__42184;
    wire N__42181;
    wire N__42178;
    wire N__42175;
    wire N__42172;
    wire N__42171;
    wire N__42170;
    wire N__42169;
    wire N__42164;
    wire N__42153;
    wire N__42146;
    wire N__42145;
    wire N__42144;
    wire N__42143;
    wire N__42142;
    wire N__42141;
    wire N__42140;
    wire N__42133;
    wire N__42132;
    wire N__42131;
    wire N__42128;
    wire N__42127;
    wire N__42126;
    wire N__42125;
    wire N__42122;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42082;
    wire N__42075;
    wire N__42072;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42057;
    wire N__42048;
    wire N__42043;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42026;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__41999;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41987;
    wire N__41982;
    wire N__41977;
    wire N__41974;
    wire N__41973;
    wire N__41972;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41960;
    wire N__41955;
    wire N__41950;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41942;
    wire N__41939;
    wire N__41934;
    wire N__41929;
    wire N__41928;
    wire N__41927;
    wire N__41926;
    wire N__41923;
    wire N__41918;
    wire N__41915;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41884;
    wire N__41881;
    wire N__41878;
    wire N__41877;
    wire N__41876;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41854;
    wire N__41853;
    wire N__41852;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41840;
    wire N__41833;
    wire N__41830;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41800;
    wire N__41799;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41721;
    wire N__41718;
    wire N__41715;
    wire N__41710;
    wire N__41707;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41695;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41624;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41612;
    wire N__41605;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41578;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41533;
    wire N__41530;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41505;
    wire N__41500;
    wire N__41497;
    wire N__41496;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41476;
    wire N__41473;
    wire N__41472;
    wire N__41471;
    wire N__41470;
    wire N__41469;
    wire N__41468;
    wire N__41467;
    wire N__41466;
    wire N__41465;
    wire N__41464;
    wire N__41463;
    wire N__41462;
    wire N__41461;
    wire N__41460;
    wire N__41459;
    wire N__41458;
    wire N__41457;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41449;
    wire N__41444;
    wire N__41441;
    wire N__41436;
    wire N__41435;
    wire N__41434;
    wire N__41433;
    wire N__41430;
    wire N__41429;
    wire N__41428;
    wire N__41423;
    wire N__41414;
    wire N__41405;
    wire N__41404;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41365;
    wire N__41358;
    wire N__41355;
    wire N__41352;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41330;
    wire N__41327;
    wire N__41320;
    wire N__41317;
    wire N__41310;
    wire N__41305;
    wire N__41298;
    wire N__41291;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41232;
    wire N__41229;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41217;
    wire N__41216;
    wire N__41213;
    wire N__41208;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41190;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41142;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41113;
    wire N__41110;
    wire N__41101;
    wire N__41098;
    wire N__41097;
    wire N__41096;
    wire N__41095;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41087;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41068;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41028;
    wire N__41027;
    wire N__41024;
    wire N__41019;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__41001;
    wire N__40996;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40938;
    wire N__40937;
    wire N__40936;
    wire N__40935;
    wire N__40932;
    wire N__40927;
    wire N__40926;
    wire N__40925;
    wire N__40924;
    wire N__40923;
    wire N__40920;
    wire N__40919;
    wire N__40916;
    wire N__40915;
    wire N__40914;
    wire N__40909;
    wire N__40908;
    wire N__40907;
    wire N__40906;
    wire N__40905;
    wire N__40904;
    wire N__40901;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40893;
    wire N__40892;
    wire N__40887;
    wire N__40886;
    wire N__40885;
    wire N__40884;
    wire N__40883;
    wire N__40882;
    wire N__40881;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40869;
    wire N__40866;
    wire N__40861;
    wire N__40858;
    wire N__40857;
    wire N__40856;
    wire N__40855;
    wire N__40854;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40846;
    wire N__40845;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40826;
    wire N__40825;
    wire N__40824;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40806;
    wire N__40801;
    wire N__40794;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40761;
    wire N__40754;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40739;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40716;
    wire N__40707;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40679;
    wire N__40674;
    wire N__40669;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40579;
    wire N__40576;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40562;
    wire N__40555;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40551;
    wire N__40550;
    wire N__40549;
    wire N__40548;
    wire N__40547;
    wire N__40546;
    wire N__40545;
    wire N__40544;
    wire N__40543;
    wire N__40542;
    wire N__40541;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40533;
    wire N__40530;
    wire N__40529;
    wire N__40528;
    wire N__40527;
    wire N__40526;
    wire N__40525;
    wire N__40524;
    wire N__40523;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40423;
    wire N__40420;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40404;
    wire N__40401;
    wire N__40396;
    wire N__40393;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40353;
    wire N__40346;
    wire N__40337;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40317;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40287;
    wire N__40286;
    wire N__40285;
    wire N__40284;
    wire N__40281;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40267;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40232;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40201;
    wire N__40200;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40186;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40170;
    wire N__40165;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40111;
    wire N__40110;
    wire N__40107;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40092;
    wire N__40085;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40071;
    wire N__40068;
    wire N__40063;
    wire N__40062;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40032;
    wire N__40027;
    wire N__40026;
    wire N__40025;
    wire N__40022;
    wire N__40017;
    wire N__40012;
    wire N__40009;
    wire N__40008;
    wire N__40005;
    wire N__40004;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39982;
    wire N__39981;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39961;
    wire N__39960;
    wire N__39955;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39924;
    wire N__39919;
    wire N__39916;
    wire N__39915;
    wire N__39914;
    wire N__39913;
    wire N__39910;
    wire N__39905;
    wire N__39900;
    wire N__39895;
    wire N__39892;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39880;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39868;
    wire N__39867;
    wire N__39866;
    wire N__39865;
    wire N__39862;
    wire N__39857;
    wire N__39854;
    wire N__39847;
    wire N__39846;
    wire N__39845;
    wire N__39844;
    wire N__39839;
    wire N__39834;
    wire N__39829;
    wire N__39828;
    wire N__39825;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39813;
    wire N__39808;
    wire N__39807;
    wire N__39806;
    wire N__39803;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39782;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39765;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39744;
    wire N__39743;
    wire N__39740;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39717;
    wire N__39712;
    wire N__39711;
    wire N__39706;
    wire N__39703;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39666;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39597;
    wire N__39596;
    wire N__39595;
    wire N__39594;
    wire N__39591;
    wire N__39590;
    wire N__39587;
    wire N__39582;
    wire N__39577;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39569;
    wire N__39568;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39515;
    wire N__39512;
    wire N__39493;
    wire N__39492;
    wire N__39491;
    wire N__39490;
    wire N__39487;
    wire N__39486;
    wire N__39483;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39433;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39402;
    wire N__39401;
    wire N__39398;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39375;
    wire N__39374;
    wire N__39371;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39345;
    wire N__39344;
    wire N__39343;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39335;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39314;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39291;
    wire N__39290;
    wire N__39289;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39264;
    wire N__39261;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39232;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39221;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39205;
    wire N__39204;
    wire N__39199;
    wire N__39196;
    wire N__39195;
    wire N__39194;
    wire N__39193;
    wire N__39192;
    wire N__39191;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39177;
    wire N__39172;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39143;
    wire N__39142;
    wire N__39137;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39076;
    wire N__39075;
    wire N__39072;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39064;
    wire N__39061;
    wire N__39060;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39004;
    wire N__39003;
    wire N__38998;
    wire N__38997;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38989;
    wire N__38986;
    wire N__38985;
    wire N__38984;
    wire N__38979;
    wire N__38978;
    wire N__38977;
    wire N__38976;
    wire N__38973;
    wire N__38972;
    wire N__38969;
    wire N__38968;
    wire N__38965;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38926;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38905;
    wire N__38902;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38880;
    wire N__38875;
    wire N__38870;
    wire N__38865;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38841;
    wire N__38838;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38752;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38674;
    wire N__38671;
    wire N__38670;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38643;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38620;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38608;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38600;
    wire N__38593;
    wire N__38590;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38520;
    wire N__38519;
    wire N__38516;
    wire N__38515;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38494;
    wire N__38493;
    wire N__38492;
    wire N__38491;
    wire N__38486;
    wire N__38481;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38458;
    wire N__38457;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38436;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38424;
    wire N__38419;
    wire N__38416;
    wire N__38415;
    wire N__38414;
    wire N__38413;
    wire N__38408;
    wire N__38403;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38362;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38354;
    wire N__38349;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38331;
    wire N__38326;
    wire N__38325;
    wire N__38322;
    wire N__38321;
    wire N__38318;
    wire N__38317;
    wire N__38314;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38293;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38266;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38248;
    wire N__38247;
    wire N__38246;
    wire N__38245;
    wire N__38238;
    wire N__38235;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38212;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38186;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38136;
    wire N__38135;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38107;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38083;
    wire N__38082;
    wire N__38081;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38068;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38046;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38019;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37929;
    wire N__37928;
    wire N__37927;
    wire N__37924;
    wire N__37923;
    wire N__37922;
    wire N__37921;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37913;
    wire N__37912;
    wire N__37907;
    wire N__37900;
    wire N__37895;
    wire N__37892;
    wire N__37887;
    wire N__37884;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37863;
    wire N__37862;
    wire N__37859;
    wire N__37858;
    wire N__37857;
    wire N__37854;
    wire N__37853;
    wire N__37852;
    wire N__37851;
    wire N__37850;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37838;
    wire N__37835;
    wire N__37828;
    wire N__37823;
    wire N__37810;
    wire N__37807;
    wire N__37806;
    wire N__37805;
    wire N__37802;
    wire N__37801;
    wire N__37800;
    wire N__37799;
    wire N__37798;
    wire N__37797;
    wire N__37796;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37780;
    wire N__37777;
    wire N__37772;
    wire N__37769;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37749;
    wire N__37748;
    wire N__37745;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37723;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37715;
    wire N__37714;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37699;
    wire N__37690;
    wire N__37687;
    wire N__37684;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37680;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37663;
    wire N__37654;
    wire N__37653;
    wire N__37652;
    wire N__37649;
    wire N__37648;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37633;
    wire N__37630;
    wire N__37621;
    wire N__37618;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37610;
    wire N__37609;
    wire N__37608;
    wire N__37603;
    wire N__37600;
    wire N__37595;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37548;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37511;
    wire N__37506;
    wire N__37503;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37467;
    wire N__37466;
    wire N__37465;
    wire N__37464;
    wire N__37463;
    wire N__37462;
    wire N__37461;
    wire N__37460;
    wire N__37455;
    wire N__37452;
    wire N__37451;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37443;
    wire N__37434;
    wire N__37429;
    wire N__37428;
    wire N__37425;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37412;
    wire N__37409;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37356;
    wire N__37345;
    wire N__37344;
    wire N__37343;
    wire N__37342;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37336;
    wire N__37335;
    wire N__37330;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37316;
    wire N__37313;
    wire N__37312;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37278;
    wire N__37275;
    wire N__37268;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37212;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37191;
    wire N__37188;
    wire N__37183;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37092;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37060;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37027;
    wire N__37024;
    wire N__37023;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37009;
    wire N__37006;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36987;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36969;
    wire N__36968;
    wire N__36967;
    wire N__36966;
    wire N__36965;
    wire N__36962;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36955;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36949;
    wire N__36944;
    wire N__36941;
    wire N__36940;
    wire N__36939;
    wire N__36932;
    wire N__36931;
    wire N__36930;
    wire N__36927;
    wire N__36926;
    wire N__36925;
    wire N__36922;
    wire N__36917;
    wire N__36912;
    wire N__36909;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36886;
    wire N__36885;
    wire N__36880;
    wire N__36877;
    wire N__36876;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36839;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36823;
    wire N__36820;
    wire N__36815;
    wire N__36810;
    wire N__36803;
    wire N__36800;
    wire N__36789;
    wire N__36778;
    wire N__36769;
    wire N__36766;
    wire N__36765;
    wire N__36764;
    wire N__36761;
    wire N__36760;
    wire N__36759;
    wire N__36758;
    wire N__36757;
    wire N__36756;
    wire N__36755;
    wire N__36750;
    wire N__36747;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36736;
    wire N__36735;
    wire N__36732;
    wire N__36731;
    wire N__36730;
    wire N__36729;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36716;
    wire N__36711;
    wire N__36708;
    wire N__36707;
    wire N__36704;
    wire N__36703;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36679;
    wire N__36670;
    wire N__36661;
    wire N__36656;
    wire N__36653;
    wire N__36648;
    wire N__36645;
    wire N__36642;
    wire N__36637;
    wire N__36634;
    wire N__36633;
    wire N__36628;
    wire N__36625;
    wire N__36624;
    wire N__36623;
    wire N__36622;
    wire N__36621;
    wire N__36618;
    wire N__36613;
    wire N__36608;
    wire N__36595;
    wire N__36590;
    wire N__36589;
    wire N__36588;
    wire N__36585;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36564;
    wire N__36561;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36538;
    wire N__36535;
    wire N__36526;
    wire N__36521;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36483;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36430;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36334;
    wire N__36331;
    wire N__36330;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36261;
    wire N__36260;
    wire N__36259;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36255;
    wire N__36254;
    wire N__36251;
    wire N__36250;
    wire N__36249;
    wire N__36248;
    wire N__36247;
    wire N__36246;
    wire N__36245;
    wire N__36240;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36196;
    wire N__36191;
    wire N__36184;
    wire N__36181;
    wire N__36180;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36169;
    wire N__36166;
    wire N__36159;
    wire N__36150;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36120;
    wire N__36117;
    wire N__36112;
    wire N__36107;
    wire N__36102;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36075;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36054;
    wire N__36049;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36037;
    wire N__36034;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36019;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__36000;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35872;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35860;
    wire N__35859;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35815;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35760;
    wire N__35757;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35719;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35706;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35688;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35663;
    wire N__35656;
    wire N__35645;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35639;
    wire N__35638;
    wire N__35637;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35621;
    wire N__35614;
    wire N__35609;
    wire N__35604;
    wire N__35587;
    wire N__35582;
    wire N__35577;
    wire N__35574;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35530;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35515;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35419;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35387;
    wire N__35380;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35292;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35247;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35134;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35111;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35079;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35059;
    wire N__35056;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34965;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34936;
    wire N__34933;
    wire N__34932;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34878;
    wire N__34873;
    wire N__34870;
    wire N__34869;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34849;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34758;
    wire N__34757;
    wire N__34754;
    wire N__34749;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34728;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34707;
    wire N__34704;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34650;
    wire N__34641;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34614;
    wire N__34611;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34594;
    wire N__34591;
    wire N__34590;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34557;
    wire N__34552;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34506;
    wire N__34501;
    wire N__34498;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34465;
    wire N__34464;
    wire N__34461;
    wire N__34456;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34441;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34386;
    wire N__34383;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34336;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34324;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34233;
    wire N__34230;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34226;
    wire N__34223;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34217;
    wire N__34212;
    wire N__34209;
    wire N__34204;
    wire N__34197;
    wire N__34194;
    wire N__34183;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34175;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34161;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34138;
    wire N__34135;
    wire N__34130;
    wire N__34127;
    wire N__34120;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34099;
    wire N__34098;
    wire N__34097;
    wire N__34096;
    wire N__34095;
    wire N__34094;
    wire N__34093;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34083;
    wire N__34078;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34021;
    wire N__34018;
    wire N__34011;
    wire N__34008;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33969;
    wire N__33966;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33931;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33916;
    wire N__33915;
    wire N__33910;
    wire N__33907;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33885;
    wire N__33882;
    wire N__33881;
    wire N__33880;
    wire N__33879;
    wire N__33878;
    wire N__33877;
    wire N__33874;
    wire N__33873;
    wire N__33870;
    wire N__33865;
    wire N__33862;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33848;
    wire N__33845;
    wire N__33840;
    wire N__33835;
    wire N__33832;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33805;
    wire N__33802;
    wire N__33801;
    wire N__33800;
    wire N__33799;
    wire N__33798;
    wire N__33797;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33785;
    wire N__33780;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33765;
    wire N__33762;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33675;
    wire N__33670;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33628;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33592;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33577;
    wire N__33574;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33526;
    wire N__33523;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33508;
    wire N__33507;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33462;
    wire N__33459;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33384;
    wire N__33383;
    wire N__33380;
    wire N__33375;
    wire N__33372;
    wire N__33367;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33330;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33270;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33127;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33088;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33004;
    wire N__33003;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32799;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32782;
    wire N__32781;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32724;
    wire N__32723;
    wire N__32722;
    wire N__32721;
    wire N__32720;
    wire N__32719;
    wire N__32718;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32705;
    wire N__32704;
    wire N__32703;
    wire N__32702;
    wire N__32701;
    wire N__32700;
    wire N__32699;
    wire N__32698;
    wire N__32697;
    wire N__32696;
    wire N__32695;
    wire N__32688;
    wire N__32679;
    wire N__32672;
    wire N__32663;
    wire N__32656;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32641;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32619;
    wire N__32618;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32605;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32581;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32567;
    wire N__32566;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32550;
    wire N__32543;
    wire N__32534;
    wire N__32527;
    wire N__32518;
    wire N__32511;
    wire N__32502;
    wire N__32495;
    wire N__32486;
    wire N__32485;
    wire N__32484;
    wire N__32483;
    wire N__32482;
    wire N__32481;
    wire N__32480;
    wire N__32479;
    wire N__32478;
    wire N__32477;
    wire N__32476;
    wire N__32475;
    wire N__32474;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32451;
    wire N__32436;
    wire N__32421;
    wire N__32420;
    wire N__32417;
    wire N__32416;
    wire N__32413;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32407;
    wire N__32404;
    wire N__32403;
    wire N__32400;
    wire N__32399;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32386;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32379;
    wire N__32378;
    wire N__32377;
    wire N__32376;
    wire N__32361;
    wire N__32360;
    wire N__32357;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32329;
    wire N__32322;
    wire N__32313;
    wire N__32306;
    wire N__32297;
    wire N__32290;
    wire N__32281;
    wire N__32274;
    wire N__32265;
    wire N__32264;
    wire N__32263;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32259;
    wire N__32258;
    wire N__32251;
    wire N__32236;
    wire N__32221;
    wire N__32206;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32193;
    wire N__32192;
    wire N__32189;
    wire N__32188;
    wire N__32185;
    wire N__32184;
    wire N__32181;
    wire N__32180;
    wire N__32177;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32154;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32129;
    wire N__32122;
    wire N__32113;
    wire N__32104;
    wire N__32089;
    wire N__32074;
    wire N__32073;
    wire N__32072;
    wire N__32071;
    wire N__32066;
    wire N__32059;
    wire N__32050;
    wire N__32043;
    wire N__32034;
    wire N__32027;
    wire N__32020;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32005;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31982;
    wire N__31977;
    wire N__31970;
    wire N__31961;
    wire N__31946;
    wire N__31939;
    wire N__31930;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31689;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31677;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31662;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31626;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31575;
    wire N__31572;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31506;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31488;
    wire N__31485;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31429;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31351;
    wire N__31350;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31295;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31273;
    wire N__31272;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31204;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31194;
    wire N__31191;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31167;
    wire N__31164;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31144;
    wire N__31141;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31127;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31090;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31060;
    wire N__31057;
    wire N__31056;
    wire N__31053;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31033;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31021;
    wire N__31018;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30973;
    wire N__30970;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30954;
    wire N__30953;
    wire N__30952;
    wire N__30949;
    wire N__30944;
    wire N__30943;
    wire N__30940;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30919;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30894;
    wire N__30889;
    wire N__30886;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30871;
    wire N__30870;
    wire N__30869;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30832;
    wire N__30829;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30814;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30786;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30768;
    wire N__30763;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30736;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30714;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30684;
    wire N__30681;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30642;
    wire N__30639;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30600;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30594;
    wire N__30593;
    wire N__30590;
    wire N__30589;
    wire N__30586;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30580;
    wire N__30579;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30575;
    wire N__30574;
    wire N__30573;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30567;
    wire N__30566;
    wire N__30565;
    wire N__30564;
    wire N__30561;
    wire N__30544;
    wire N__30535;
    wire N__30526;
    wire N__30517;
    wire N__30508;
    wire N__30507;
    wire N__30506;
    wire N__30505;
    wire N__30502;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30493;
    wire N__30484;
    wire N__30475;
    wire N__30466;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30411;
    wire N__30408;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30393;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30372;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30288;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30255;
    wire N__30252;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30219;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30033;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29884;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29874;
    wire N__29869;
    wire N__29868;
    wire N__29867;
    wire N__29866;
    wire N__29863;
    wire N__29858;
    wire N__29857;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29797;
    wire N__29796;
    wire N__29793;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29776;
    wire N__29775;
    wire N__29772;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29736;
    wire N__29735;
    wire N__29730;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29624;
    wire N__29619;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29604;
    wire N__29599;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29591;
    wire N__29590;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29569;
    wire N__29568;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29553;
    wire N__29550;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29540;
    wire N__29537;
    wire N__29532;
    wire N__29527;
    wire N__29524;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29496;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29452;
    wire N__29451;
    wire N__29450;
    wire N__29447;
    wire N__29442;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29424;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29328;
    wire N__29325;
    wire N__29324;
    wire N__29321;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29305;
    wire N__29304;
    wire N__29303;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29285;
    wire N__29284;
    wire N__29283;
    wire N__29282;
    wire N__29281;
    wire N__29280;
    wire N__29273;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29264;
    wire N__29261;
    wire N__29256;
    wire N__29253;
    wire N__29244;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29203;
    wire N__29200;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29170;
    wire N__29169;
    wire N__29168;
    wire N__29165;
    wire N__29164;
    wire N__29163;
    wire N__29162;
    wire N__29161;
    wire N__29160;
    wire N__29159;
    wire N__29158;
    wire N__29149;
    wire N__29146;
    wire N__29145;
    wire N__29144;
    wire N__29143;
    wire N__29142;
    wire N__29139;
    wire N__29134;
    wire N__29129;
    wire N__29126;
    wire N__29121;
    wire N__29118;
    wire N__29113;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29058;
    wire N__29057;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29043;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28992;
    wire N__28989;
    wire N__28988;
    wire N__28985;
    wire N__28980;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28894;
    wire N__28891;
    wire N__28890;
    wire N__28885;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28870;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28855;
    wire N__28854;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28819;
    wire N__28816;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28726;
    wire N__28725;
    wire N__28722;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28705;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28674;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28552;
    wire N__28549;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28492;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28474;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28459;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28447;
    wire N__28444;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28432;
    wire N__28429;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28417;
    wire N__28414;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28402;
    wire N__28399;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28387;
    wire N__28384;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28372;
    wire N__28369;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28354;
    wire N__28351;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28336;
    wire N__28333;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28321;
    wire N__28318;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28306;
    wire N__28303;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28245;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28231;
    wire N__28228;
    wire N__28223;
    wire N__28220;
    wire N__28213;
    wire N__28212;
    wire N__28207;
    wire N__28206;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28174;
    wire N__28171;
    wire N__28170;
    wire N__28169;
    wire N__28164;
    wire N__28161;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28131;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28105;
    wire N__28102;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28090;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28078;
    wire N__28075;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28045;
    wire N__28042;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28030;
    wire N__28027;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28015;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27985;
    wire N__27982;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27927;
    wire N__27926;
    wire N__27923;
    wire N__27918;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27889;
    wire N__27886;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27871;
    wire N__27868;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27856;
    wire N__27853;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27804;
    wire N__27799;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27756;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27738;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27723;
    wire N__27718;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27710;
    wire N__27707;
    wire N__27702;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27687;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27679;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27665;
    wire N__27662;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27633;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27592;
    wire N__27591;
    wire N__27590;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27531;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27503;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27435;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27417;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27402;
    wire N__27399;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27376;
    wire N__27375;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27331;
    wire N__27328;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27297;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27274;
    wire N__27273;
    wire N__27270;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27250;
    wire N__27249;
    wire N__27246;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27226;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27211;
    wire N__27208;
    wire N__27207;
    wire N__27204;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27189;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27154;
    wire N__27153;
    wire N__27150;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27130;
    wire N__27129;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27109;
    wire N__27108;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27085;
    wire N__27082;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27051;
    wire N__27048;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26937;
    wire N__26932;
    wire N__26929;
    wire N__26928;
    wire N__26927;
    wire N__26924;
    wire N__26919;
    wire N__26916;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26903;
    wire N__26900;
    wire N__26895;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26883;
    wire N__26882;
    wire N__26881;
    wire N__26880;
    wire N__26875;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26817;
    wire N__26816;
    wire N__26815;
    wire N__26810;
    wire N__26805;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26781;
    wire N__26780;
    wire N__26775;
    wire N__26772;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26716;
    wire N__26713;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26701;
    wire N__26698;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26686;
    wire N__26683;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26671;
    wire N__26668;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26656;
    wire N__26653;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26641;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26616;
    wire N__26615;
    wire N__26614;
    wire N__26613;
    wire N__26612;
    wire N__26611;
    wire N__26610;
    wire N__26609;
    wire N__26608;
    wire N__26607;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26603;
    wire N__26596;
    wire N__26595;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26581;
    wire N__26578;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26542;
    wire N__26541;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26504;
    wire N__26499;
    wire N__26494;
    wire N__26493;
    wire N__26492;
    wire N__26491;
    wire N__26490;
    wire N__26489;
    wire N__26488;
    wire N__26487;
    wire N__26486;
    wire N__26485;
    wire N__26484;
    wire N__26483;
    wire N__26482;
    wire N__26479;
    wire N__26478;
    wire N__26475;
    wire N__26474;
    wire N__26473;
    wire N__26472;
    wire N__26471;
    wire N__26466;
    wire N__26453;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26419;
    wire N__26416;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26400;
    wire N__26397;
    wire N__26392;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26366;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26313;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26295;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26239;
    wire N__26238;
    wire N__26237;
    wire N__26236;
    wire N__26235;
    wire N__26234;
    wire N__26233;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26229;
    wire N__26228;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26170;
    wire N__26161;
    wire N__26152;
    wire N__26143;
    wire N__26134;
    wire N__26133;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26047;
    wire N__26046;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26031;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25977;
    wire N__25974;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25968;
    wire N__25967;
    wire N__25966;
    wire N__25965;
    wire N__25964;
    wire N__25963;
    wire N__25960;
    wire N__25959;
    wire N__25958;
    wire N__25957;
    wire N__25956;
    wire N__25955;
    wire N__25954;
    wire N__25951;
    wire N__25942;
    wire N__25933;
    wire N__25922;
    wire N__25915;
    wire N__25914;
    wire N__25913;
    wire N__25912;
    wire N__25911;
    wire N__25910;
    wire N__25909;
    wire N__25908;
    wire N__25907;
    wire N__25906;
    wire N__25905;
    wire N__25902;
    wire N__25901;
    wire N__25900;
    wire N__25897;
    wire N__25896;
    wire N__25895;
    wire N__25884;
    wire N__25875;
    wire N__25866;
    wire N__25859;
    wire N__25848;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25791;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25698;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25617;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25600;
    wire N__25599;
    wire N__25598;
    wire N__25595;
    wire N__25594;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25566;
    wire N__25565;
    wire N__25558;
    wire N__25555;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25543;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25531;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25516;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25504;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25492;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25473;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25456;
    wire N__25453;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25441;
    wire N__25440;
    wire N__25435;
    wire N__25432;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25420;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25408;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25393;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25363;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25351;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25336;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25277;
    wire N__25272;
    wire N__25269;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25203;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25188;
    wire N__25185;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25172;
    wire N__25167;
    wire N__25164;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25152;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25118;
    wire N__25113;
    wire N__25110;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25088;
    wire N__25083;
    wire N__25080;
    wire N__25075;
    wire N__25072;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25064;
    wire N__25059;
    wire N__25056;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25032;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25017;
    wire N__25014;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24984;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24891;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24855;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24843;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24831;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24814;
    wire N__24813;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire tx_enable;
    wire LED_c;
    wire \c0.n18673 ;
    wire \c0.n18661 ;
    wire n39;
    wire bfn_9_7_0_;
    wire \quad_counter0.n17222 ;
    wire \quad_counter0.n17223 ;
    wire \quad_counter0.n17224 ;
    wire \quad_counter0.n17225 ;
    wire \quad_counter0.n17226 ;
    wire \quad_counter0.n17227 ;
    wire \quad_counter0.n17228 ;
    wire \quad_counter0.n17229 ;
    wire bfn_9_8_0_;
    wire \quad_counter0.n17230 ;
    wire \quad_counter0.n17231 ;
    wire \quad_counter0.n17232 ;
    wire \quad_counter0.n17233 ;
    wire \quad_counter0.n17234 ;
    wire \quad_counter0.n17235 ;
    wire \quad_counter0.n17236 ;
    wire data_out_frame_6_6;
    wire data_out_frame_5_1;
    wire data_out_frame_7_6;
    wire bfn_9_14_0_;
    wire \quad_counter0.b_delay_counter_1 ;
    wire \quad_counter0.n13182 ;
    wire \quad_counter0.n17207 ;
    wire \quad_counter0.n17208 ;
    wire \quad_counter0.n17209 ;
    wire \quad_counter0.b_delay_counter_4 ;
    wire \quad_counter0.n13197 ;
    wire \quad_counter0.n17210 ;
    wire \quad_counter0.n17211 ;
    wire \quad_counter0.n17212 ;
    wire \quad_counter0.b_delay_counter_7 ;
    wire \quad_counter0.n13214 ;
    wire \quad_counter0.n17213 ;
    wire \quad_counter0.n17214 ;
    wire bfn_9_15_0_;
    wire \quad_counter0.n17215 ;
    wire \quad_counter0.n17216 ;
    wire \quad_counter0.b_delay_counter_11 ;
    wire \quad_counter0.n13257 ;
    wire \quad_counter0.n17217 ;
    wire \quad_counter0.n17218 ;
    wire \quad_counter0.b_delay_counter_13 ;
    wire \quad_counter0.n13263 ;
    wire \quad_counter0.n17219 ;
    wire \quad_counter0.n17220 ;
    wire \quad_counter0.n17221 ;
    wire \quad_counter0.n13260 ;
    wire \quad_counter0.b_delay_counter_12 ;
    wire \quad_counter0.n13444 ;
    wire \quad_counter0.n13266 ;
    wire \quad_counter0.b_delay_counter_14 ;
    wire \quad_counter0.n13248 ;
    wire \quad_counter0.b_delay_counter_8 ;
    wire \quad_counter0.n13203 ;
    wire \quad_counter0.b_delay_counter_6 ;
    wire \quad_counter0.b_delay_counter_0 ;
    wire \quad_counter0.n13251 ;
    wire \quad_counter0.b_delay_counter_9 ;
    wire \quad_counter0.n13194 ;
    wire \quad_counter0.b_delay_counter_3 ;
    wire \quad_counter0.n13200 ;
    wire \quad_counter0.b_delay_counter_5 ;
    wire \c0.n18649 ;
    wire \c0.n18639 ;
    wire \c0.n18663 ;
    wire a_delay_counter_15__N_2916;
    wire n12447;
    wire PIN_7_c;
    wire quadA_delayed;
    wire \quad_counter0.a_delay_counter_15 ;
    wire \quad_counter0.a_delay_counter_8 ;
    wire \quad_counter0.a_delay_counter_1 ;
    wire \quad_counter0.a_delay_counter_6 ;
    wire \quad_counter0.a_delay_counter_9 ;
    wire \quad_counter0.a_delay_counter_7 ;
    wire \quad_counter0.n18_cascade_ ;
    wire a_delay_counter_0;
    wire \quad_counter0.n20_cascade_ ;
    wire \quad_counter0.a_delay_counter_2 ;
    wire n11349;
    wire \quad_counter0.a_delay_counter_5 ;
    wire \quad_counter0.a_delay_counter_10 ;
    wire \quad_counter0.a_delay_counter_12 ;
    wire \quad_counter0.a_delay_counter_3 ;
    wire \quad_counter0.n20954 ;
    wire \quad_counter0.a_delay_counter_4 ;
    wire \quad_counter0.a_delay_counter_11 ;
    wire \quad_counter0.a_delay_counter_14 ;
    wire \quad_counter0.a_delay_counter_13 ;
    wire \quad_counter0.n19 ;
    wire bfn_10_9_0_;
    wire \quad_counter0.count_direction ;
    wire n2279;
    wire \quad_counter0.n17282 ;
    wire n2278;
    wire \quad_counter0.n17283 ;
    wire encoder0_position_2;
    wire n2277;
    wire \quad_counter0.n17284 ;
    wire encoder0_position_3;
    wire n2276;
    wire \quad_counter0.n17285 ;
    wire \quad_counter0.n17286 ;
    wire \quad_counter0.n17287 ;
    wire \quad_counter0.n17288 ;
    wire \quad_counter0.n17289 ;
    wire bfn_10_10_0_;
    wire \quad_counter0.n17290 ;
    wire \quad_counter0.n17291 ;
    wire \quad_counter0.n17292 ;
    wire \quad_counter0.n17293 ;
    wire \quad_counter0.n17294 ;
    wire \quad_counter0.n17295 ;
    wire \quad_counter0.n17296 ;
    wire \quad_counter0.n17297 ;
    wire bfn_10_11_0_;
    wire \quad_counter0.n17298 ;
    wire \quad_counter0.n17299 ;
    wire n2261;
    wire \quad_counter0.n17300 ;
    wire n2260;
    wire \quad_counter0.n17301 ;
    wire n2259;
    wire \quad_counter0.n17302 ;
    wire n2258;
    wire \quad_counter0.n17303 ;
    wire encoder0_position_22;
    wire n2257;
    wire \quad_counter0.n17304 ;
    wire \quad_counter0.n17305 ;
    wire n2256;
    wire bfn_10_12_0_;
    wire n2255;
    wire \quad_counter0.n17306 ;
    wire n2254;
    wire \quad_counter0.n17307 ;
    wire \quad_counter0.n17308 ;
    wire \quad_counter0.n17309 ;
    wire \quad_counter0.n17310 ;
    wire \quad_counter0.n17311 ;
    wire \quad_counter0.n17312 ;
    wire \quad_counter0.n17313 ;
    wire \quad_counter0.n2228 ;
    wire bfn_10_13_0_;
    wire n2275;
    wire n2272;
    wire n2274;
    wire n2248;
    wire \c0.n5_adj_3471 ;
    wire encoder0_position_5;
    wire data_out_frame_9_6;
    wire \quad_counter0.n13254 ;
    wire \quad_counter0.b_delay_counter_10 ;
    wire \quad_counter0.n13269 ;
    wire \quad_counter0.b_delay_counter_15 ;
    wire \quad_counter0.n26_adj_2991 ;
    wire \quad_counter0.n27_adj_2992 ;
    wire \quad_counter0.n28_adj_2990 ;
    wire \quad_counter0.n25_adj_2993 ;
    wire n11347;
    wire n11347_cascade_;
    wire \quad_counter0.n21603 ;
    wire data_out_frame_10_6;
    wire \c0.n21629 ;
    wire PIN_8_c;
    wire quadB_delayed;
    wire \quad_counter0.n13187 ;
    wire \quad_counter0.b_delay_counter_2 ;
    wire \c0.n21331_cascade_ ;
    wire \c0.n17354_cascade_ ;
    wire \c0.n21521 ;
    wire \c0.tx.n6_cascade_ ;
    wire \c0.n15938_cascade_ ;
    wire \c0.tx.r_Clock_Count_0 ;
    wire bfn_10_18_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n17274 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n17275 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n17276 ;
    wire \c0.tx.r_Clock_Count_4 ;
    wire \c0.tx.n17277 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire \c0.tx.n17278 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.n17279 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.n17280 ;
    wire \c0.tx.n17281 ;
    wire bfn_10_19_0_;
    wire \c0.n18671 ;
    wire \c0.n18617 ;
    wire \quad_counter1.n25_adj_3577_cascade_ ;
    wire n11343_cascade_;
    wire n12417_cascade_;
    wire \quad_counter1.n28_adj_3574 ;
    wire PIN_13_c;
    wire n11343;
    wire quadB_delayed_adj_3585;
    wire \quad_counter1.n26_adj_3575 ;
    wire \quad_counter1.n27_adj_3576 ;
    wire \quad_counter1.n16_cascade_ ;
    wire \quad_counter1.n24_adj_3578_cascade_ ;
    wire n11351;
    wire B_filtered;
    wire \quad_counter0.B_delayed ;
    wire \quad_counter1.n6 ;
    wire A_filtered;
    wire \quad_counter0.A_delayed ;
    wire \quad_counter1.n22 ;
    wire n2269;
    wire n2268;
    wire n2267;
    wire n2266;
    wire n2265;
    wire n2264;
    wire encoder0_position_15;
    wire n2263;
    wire n2262;
    wire data_out_frame_6_4;
    wire encoder0_position_25;
    wire encoder0_position_10;
    wire encoder0_position_20;
    wire data_out_frame_7_4;
    wire n2253;
    wire n2249;
    wire encoder0_position_30;
    wire data_out_frame_6_1;
    wire encoder0_position_1;
    wire n2251;
    wire encoder0_position_28;
    wire encoder0_position_16;
    wire encoder0_position_14;
    wire data_out_frame_8_6;
    wire encoder0_position_4;
    wire \c0.n21632 ;
    wire \c0.n21299 ;
    wire data_out_frame_8_7;
    wire \c0.n21626_cascade_ ;
    wire encoder0_position_7;
    wire data_out_frame_9_7;
    wire \c0.n11_adj_3472 ;
    wire \c0.n11_adj_3479 ;
    wire \c0.n11_adj_3444_cascade_ ;
    wire \c0.n21289_cascade_ ;
    wire \c0.n55_cascade_ ;
    wire \c0.n14301_cascade_ ;
    wire \c0.n15942 ;
    wire n6866;
    wire data_out_frame_10_4;
    wire \c0.n21288 ;
    wire n2273;
    wire encoder0_position_6;
    wire \c0.n21517 ;
    wire \c0.n21506_cascade_ ;
    wire \c0.n55 ;
    wire \c0.r_Bit_Index_2 ;
    wire \c0.n21414_cascade_ ;
    wire \c0.n11 ;
    wire \c0.n15938 ;
    wire \c0.tx.n8 ;
    wire \c0.tx.n4 ;
    wire \c0.tx.n21179_cascade_ ;
    wire \c0.r_Clock_Count_8 ;
    wire \c0.tx.n12759 ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n18669 ;
    wire \c0.n18679 ;
    wire \c0.n18637 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n18635 ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n18623 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n18665 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.n18651 ;
    wire \c0.n18625 ;
    wire \c0.n18641 ;
    wire b_delay_counter_0;
    wire n187;
    wire bfn_12_5_0_;
    wire \quad_counter1.b_delay_counter_1 ;
    wire \quad_counter1.n17237 ;
    wire \quad_counter1.b_delay_counter_2 ;
    wire \quad_counter1.n17238 ;
    wire \quad_counter1.b_delay_counter_3 ;
    wire \quad_counter1.n17239 ;
    wire \quad_counter1.b_delay_counter_4 ;
    wire \quad_counter1.n17240 ;
    wire \quad_counter1.b_delay_counter_5 ;
    wire \quad_counter1.n17241 ;
    wire \quad_counter1.b_delay_counter_6 ;
    wire \quad_counter1.n17242 ;
    wire \quad_counter1.b_delay_counter_7 ;
    wire \quad_counter1.n17243 ;
    wire \quad_counter1.n17244 ;
    wire \quad_counter1.b_delay_counter_8 ;
    wire bfn_12_6_0_;
    wire \quad_counter1.b_delay_counter_9 ;
    wire \quad_counter1.n17245 ;
    wire \quad_counter1.b_delay_counter_10 ;
    wire \quad_counter1.n17246 ;
    wire \quad_counter1.b_delay_counter_11 ;
    wire \quad_counter1.n17247 ;
    wire \quad_counter1.b_delay_counter_12 ;
    wire \quad_counter1.n17248 ;
    wire \quad_counter1.b_delay_counter_13 ;
    wire \quad_counter1.n17249 ;
    wire \quad_counter1.b_delay_counter_14 ;
    wire \quad_counter1.n17250 ;
    wire \quad_counter1.n17251 ;
    wire \quad_counter1.b_delay_counter_15 ;
    wire n12417;
    wire b_delay_counter_15__N_2933;
    wire PIN_12_c;
    wire quadA_delayed_adj_3584;
    wire a_delay_counter_15__N_2916_adj_3589_cascade_;
    wire \quad_counter1.n20 ;
    wire a_delay_counter_0_adj_3583;
    wire n39_adj_3587;
    wire bfn_12_8_0_;
    wire \quad_counter1.a_delay_counter_1 ;
    wire \quad_counter1.n17252 ;
    wire \quad_counter1.a_delay_counter_2 ;
    wire \quad_counter1.n17253 ;
    wire \quad_counter1.a_delay_counter_3 ;
    wire \quad_counter1.n17254 ;
    wire \quad_counter1.a_delay_counter_4 ;
    wire \quad_counter1.n17255 ;
    wire \quad_counter1.a_delay_counter_5 ;
    wire \quad_counter1.n17256 ;
    wire \quad_counter1.a_delay_counter_6 ;
    wire \quad_counter1.n17257 ;
    wire \quad_counter1.a_delay_counter_7 ;
    wire \quad_counter1.n17258 ;
    wire \quad_counter1.n17259 ;
    wire \quad_counter1.a_delay_counter_8 ;
    wire bfn_12_9_0_;
    wire \quad_counter1.a_delay_counter_9 ;
    wire \quad_counter1.n17260 ;
    wire \quad_counter1.a_delay_counter_10 ;
    wire \quad_counter1.n17261 ;
    wire \quad_counter1.a_delay_counter_11 ;
    wire \quad_counter1.n17262 ;
    wire \quad_counter1.a_delay_counter_12 ;
    wire \quad_counter1.n17263 ;
    wire \quad_counter1.a_delay_counter_13 ;
    wire \quad_counter1.n17264 ;
    wire \quad_counter1.a_delay_counter_14 ;
    wire \quad_counter1.n17265 ;
    wire \quad_counter1.n17266 ;
    wire \quad_counter1.a_delay_counter_15 ;
    wire n12477;
    wire a_delay_counter_15__N_2916_adj_3589;
    wire data_out_frame_9_2;
    wire data_out_frame_8_2;
    wire \c0.n21650 ;
    wire \c0.n21564_cascade_ ;
    wire n2270;
    wire n2250;
    wire encoder0_position_13;
    wire data_out_frame_11_6;
    wire n2271;
    wire data_out_frame_11_4;
    wire \c0.n5_adj_3033 ;
    wire data_out_frame_12_6;
    wire encoder0_position_17;
    wire data_out_frame_7_1;
    wire \c0.n6_adj_3324 ;
    wire data_out_frame_13_3;
    wire data_out_frame_12_7;
    wire data_out_frame_11_3;
    wire data_out_frame_10_3;
    wire encoder0_position_12;
    wire data_out_frame_13_6;
    wire \c0.n21301 ;
    wire \c0.n21653 ;
    wire \c0.n21305 ;
    wire \c0.n21570 ;
    wire \c0.n21307_cascade_ ;
    wire \c0.n21577 ;
    wire n21578_cascade_;
    wire n21656;
    wire data_out_frame_13_7;
    wire \c0.n21467 ;
    wire \c0.tx.n21330 ;
    wire n9_adj_3588;
    wire r_Tx_Data_6;
    wire \c0.n9753_cascade_ ;
    wire data_out_frame_12_3;
    wire \c0.n21456 ;
    wire \c0.r_Bit_Index_1 ;
    wire \c0.n21614 ;
    wire \c0.n32 ;
    wire \c0.n2_adj_3556_cascade_ ;
    wire \c0.n7_adj_3557 ;
    wire \c0.n21329 ;
    wire \c0.n19001_cascade_ ;
    wire \c0.n30_adj_3559 ;
    wire \c0.n12498 ;
    wire \c0.n15920 ;
    wire r_SM_Main_1_adj_3592;
    wire n4_adj_3580;
    wire n9_adj_3591;
    wire r_Tx_Data_4;
    wire \c0.n12512 ;
    wire \c0.r_SM_Main_0 ;
    wire \c0.n19023 ;
    wire \c0.n18609 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n10_adj_3488 ;
    wire \c0.n15850_cascade_ ;
    wire \c0.n11427_cascade_ ;
    wire \c0.n16_adj_3484 ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n19045_cascade_ ;
    wire \c0.n4_adj_3046 ;
    wire \c0.n19045 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n10_adj_3438 ;
    wire \c0.n19050 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.n63 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n18659 ;
    wire \c0.n19146 ;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.n18633 ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n17_adj_3486 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n18677 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.n18601 ;
    wire \c0.n6_adj_3143_cascade_ ;
    wire \c0.n4_adj_3227 ;
    wire \quad_counter1.A_delayed ;
    wire B_filtered_adj_3582;
    wire \quad_counter1.B_delayed ;
    wire A_filtered_adj_3581;
    wire bfn_13_9_0_;
    wire \quad_counter1.count_direction ;
    wire \quad_counter1.n17314 ;
    wire \quad_counter1.n17315 ;
    wire n2343;
    wire \quad_counter1.n17316 ;
    wire \quad_counter1.n17317 ;
    wire n2341;
    wire \quad_counter1.n17318 ;
    wire \quad_counter1.n17319 ;
    wire encoder1_position_6;
    wire n2339;
    wire \quad_counter1.n17320 ;
    wire \quad_counter1.n17321 ;
    wire encoder1_position_7;
    wire n2338;
    wire bfn_13_10_0_;
    wire n2337;
    wire \quad_counter1.n17322 ;
    wire n2336;
    wire \quad_counter1.n17323 ;
    wire encoder1_position_10;
    wire n2335;
    wire \quad_counter1.n17324 ;
    wire encoder1_position_11;
    wire n2334;
    wire \quad_counter1.n17325 ;
    wire \quad_counter1.n17326 ;
    wire encoder1_position_13;
    wire n2332;
    wire \quad_counter1.n17327 ;
    wire encoder1_position_14;
    wire n2331;
    wire \quad_counter1.n17328 ;
    wire \quad_counter1.n17329 ;
    wire encoder1_position_15;
    wire n2330;
    wire bfn_13_11_0_;
    wire encoder1_position_16;
    wire n2329;
    wire \quad_counter1.n17330 ;
    wire n2328;
    wire \quad_counter1.n17331 ;
    wire n2327;
    wire \quad_counter1.n17332 ;
    wire encoder1_position_19;
    wire n2326;
    wire \quad_counter1.n17333 ;
    wire encoder1_position_20;
    wire n2325;
    wire \quad_counter1.n17334 ;
    wire \quad_counter1.n17335 ;
    wire encoder1_position_22;
    wire n2323;
    wire \quad_counter1.n17336 ;
    wire \quad_counter1.n17337 ;
    wire bfn_13_12_0_;
    wire n2321;
    wire \quad_counter1.n17338 ;
    wire \quad_counter1.n17339 ;
    wire n2319;
    wire \quad_counter1.n17340 ;
    wire encoder1_position_27;
    wire n2318;
    wire \quad_counter1.n17341 ;
    wire \quad_counter1.n17342 ;
    wire \quad_counter1.n17343 ;
    wire encoder1_position_30;
    wire n2315;
    wire \quad_counter1.n17344 ;
    wire \quad_counter1.n17345 ;
    wire \quad_counter1.n2301 ;
    wire bfn_13_13_0_;
    wire n2314;
    wire n2345;
    wire data_out_frame_12_5;
    wire encoder1_position_4;
    wire data_out_frame_13_4;
    wire encoder1_position_31;
    wire n2320;
    wire r_Tx_Data_5;
    wire data_out_frame_9_4;
    wire data_out_frame_8_4;
    wire \c0.n21287 ;
    wire encoder0_position_9;
    wire encoder1_position_24;
    wire \c0.data_out_frame_0_4 ;
    wire encoder0_position_8;
    wire encoder0_position_0;
    wire encoder1_position_25;
    wire encoder1_position_2;
    wire encoder1_position_17;
    wire data_out_frame_13_2;
    wire data_out_frame_12_2;
    wire \c0.n11_adj_3108 ;
    wire data_out_frame_10_1;
    wire data_out_frame_11_1;
    wire data_out_frame_13_5;
    wire \c0.r_SM_Main_2_N_2547_0 ;
    wire tx_active;
    wire \c0.n15842 ;
    wire \c0.n11_adj_3404 ;
    wire \c0.n7_adj_3333 ;
    wire data_out_frame_9_1;
    wire \c0.n21605 ;
    wire data_out_frame_8_1;
    wire \c0.n21608_cascade_ ;
    wire \c0.r_Tx_Data_0 ;
    wire \c0.n21466 ;
    wire encoder1_position_9;
    wire \c0.n21566 ;
    wire n10_cascade_;
    wire r_Tx_Data_3;
    wire data_out_frame_12_1;
    wire \c0.n11_adj_3104 ;
    wire n10_adj_3593;
    wire r_Tx_Data_2;
    wire bfn_13_18_0_;
    wire \c0.n17346 ;
    wire \c0.n17347 ;
    wire \c0.n17348 ;
    wire \c0.n17349 ;
    wire \c0.n17350 ;
    wire \c0.n17351 ;
    wire \c0.n17352 ;
    wire \c0.n19052 ;
    wire \c0.n6_adj_3338 ;
    wire \c0.n12326 ;
    wire \c0.n12326_cascade_ ;
    wire \c0.n12758 ;
    wire \c0.n4_adj_3263_cascade_ ;
    wire \c0.n936_cascade_ ;
    wire \c0.tx_transmit_N_2443 ;
    wire \c0.n21420 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n18627 ;
    wire \c0.n19650 ;
    wire \c0.n19638_cascade_ ;
    wire \c0.FRAME_MATCHER_state_31_N_1864_2 ;
    wire \c0.n6_adj_3521_cascade_ ;
    wire \c0.n936 ;
    wire \c0.n11_adj_3370 ;
    wire \c0.n19638 ;
    wire \c0.n6_adj_3515_cascade_ ;
    wire \c0.n5_adj_3516 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.n18681 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n18657 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n18629 ;
    wire bfn_14_5_0_;
    wire \c0.n17176 ;
    wire \c0.n2_adj_3144 ;
    wire \c0.n17177 ;
    wire \c0.n2_adj_3145 ;
    wire \c0.n17178 ;
    wire \c0.n17179 ;
    wire \c0.n17180 ;
    wire \c0.n17180_THRU_CRY_0_THRU_CO ;
    wire \c0.n17180_THRU_CRY_1_THRU_CO ;
    wire \c0.n17180_THRU_CRY_2_THRU_CO ;
    wire bfn_14_6_0_;
    wire \c0.n17181 ;
    wire \c0.n17181_THRU_CRY_0_THRU_CO ;
    wire \c0.n17181_THRU_CRY_1_THRU_CO ;
    wire \c0.n17181_THRU_CRY_2_THRU_CO ;
    wire \c0.n17181_THRU_CRY_3_THRU_CO ;
    wire \c0.n17181_THRU_CRY_4_THRU_CO ;
    wire \c0.n17181_THRU_CRY_5_THRU_CO ;
    wire \c0.n17181_THRU_CRY_6_THRU_CO ;
    wire bfn_14_7_0_;
    wire \c0.n17182 ;
    wire \c0.n17182_THRU_CRY_0_THRU_CO ;
    wire \c0.n17182_THRU_CRY_1_THRU_CO ;
    wire \c0.n17182_THRU_CRY_2_THRU_CO ;
    wire \c0.n17182_THRU_CRY_3_THRU_CO ;
    wire \c0.n17182_THRU_CRY_4_THRU_CO ;
    wire \c0.n17182_THRU_CRY_5_THRU_CO ;
    wire \c0.n17182_THRU_CRY_6_THRU_CO ;
    wire bfn_14_8_0_;
    wire \c0.n17183 ;
    wire \c0.n17183_THRU_CRY_0_THRU_CO ;
    wire \c0.n17183_THRU_CRY_1_THRU_CO ;
    wire \c0.n17183_THRU_CRY_2_THRU_CO ;
    wire \c0.n17183_THRU_CRY_3_THRU_CO ;
    wire \c0.n17183_THRU_CRY_4_THRU_CO ;
    wire \c0.n17183_THRU_CRY_5_THRU_CO ;
    wire \c0.n17183_THRU_CRY_6_THRU_CO ;
    wire bfn_14_9_0_;
    wire \c0.n17184 ;
    wire \c0.n17184_THRU_CRY_0_THRU_CO ;
    wire \c0.n17184_THRU_CRY_1_THRU_CO ;
    wire \c0.n17184_THRU_CRY_2_THRU_CO ;
    wire \c0.n17184_THRU_CRY_3_THRU_CO ;
    wire \c0.n17184_THRU_CRY_4_THRU_CO ;
    wire \c0.n17184_THRU_CRY_5_THRU_CO ;
    wire \c0.n17184_THRU_CRY_6_THRU_CO ;
    wire bfn_14_10_0_;
    wire \c0.n17185 ;
    wire \c0.n17185_THRU_CRY_0_THRU_CO ;
    wire \c0.n17185_THRU_CRY_1_THRU_CO ;
    wire \c0.n17185_THRU_CRY_2_THRU_CO ;
    wire \c0.n17185_THRU_CRY_3_THRU_CO ;
    wire \c0.n17185_THRU_CRY_4_THRU_CO ;
    wire \c0.n17185_THRU_CRY_5_THRU_CO ;
    wire \c0.n17185_THRU_CRY_6_THRU_CO ;
    wire bfn_14_11_0_;
    wire \c0.n17186 ;
    wire \c0.n17186_THRU_CRY_0_THRU_CO ;
    wire \c0.n17186_THRU_CRY_1_THRU_CO ;
    wire \c0.n17186_THRU_CRY_2_THRU_CO ;
    wire \c0.n17186_THRU_CRY_3_THRU_CO ;
    wire \c0.n17186_THRU_CRY_4_THRU_CO ;
    wire \c0.n17186_THRU_CRY_5_THRU_CO ;
    wire \c0.n17186_THRU_CRY_6_THRU_CO ;
    wire bfn_14_12_0_;
    wire \c0.n17187 ;
    wire \c0.n17187_THRU_CRY_0_THRU_CO ;
    wire \c0.n17187_THRU_CRY_1_THRU_CO ;
    wire \c0.n17187_THRU_CRY_2_THRU_CO ;
    wire \c0.n17187_THRU_CRY_3_THRU_CO ;
    wire \c0.n17187_THRU_CRY_4_THRU_CO ;
    wire \c0.n17187_THRU_CRY_5_THRU_CO ;
    wire \c0.n17187_THRU_CRY_6_THRU_CO ;
    wire bfn_14_13_0_;
    wire \c0.n17188 ;
    wire \c0.n17188_THRU_CRY_0_THRU_CO ;
    wire \c0.n17188_THRU_CRY_1_THRU_CO ;
    wire \c0.n17188_THRU_CRY_2_THRU_CO ;
    wire \c0.n17188_THRU_CRY_3_THRU_CO ;
    wire \c0.n17188_THRU_CRY_4_THRU_CO ;
    wire \c0.n17188_THRU_CRY_5_THRU_CO ;
    wire \c0.n17188_THRU_CRY_6_THRU_CO ;
    wire bfn_14_14_0_;
    wire \c0.n6_adj_3162 ;
    wire \c0.n17189 ;
    wire \c0.n17189_THRU_CRY_0_THRU_CO ;
    wire \c0.n17189_THRU_CRY_1_THRU_CO ;
    wire \c0.n17189_THRU_CRY_2_THRU_CO ;
    wire \c0.n17189_THRU_CRY_3_THRU_CO ;
    wire \c0.n17189_THRU_CRY_4_THRU_CO ;
    wire \c0.n17189_THRU_CRY_5_THRU_CO ;
    wire \c0.n17189_THRU_CRY_6_THRU_CO ;
    wire bfn_14_15_0_;
    wire \c0.n17190 ;
    wire \c0.n17190_THRU_CRY_0_THRU_CO ;
    wire \c0.n17190_THRU_CRY_1_THRU_CO ;
    wire \c0.n17190_THRU_CRY_2_THRU_CO ;
    wire \c0.n17190_THRU_CRY_3_THRU_CO ;
    wire \c0.n17190_THRU_CRY_4_THRU_CO ;
    wire \c0.n17190_THRU_CRY_5_THRU_CO ;
    wire \c0.n17190_THRU_CRY_6_THRU_CO ;
    wire bfn_14_16_0_;
    wire \c0.n17191 ;
    wire \c0.n17191_THRU_CRY_0_THRU_CO ;
    wire \c0.n17191_THRU_CRY_1_THRU_CO ;
    wire \c0.n17191_THRU_CRY_2_THRU_CO ;
    wire \c0.n17191_THRU_CRY_3_THRU_CO ;
    wire \c0.n17191_THRU_CRY_4_THRU_CO ;
    wire \c0.n17191_THRU_CRY_5_THRU_CO ;
    wire \c0.n17191_THRU_CRY_6_THRU_CO ;
    wire bfn_14_17_0_;
    wire \c0.n17192 ;
    wire \c0.n17192_THRU_CRY_0_THRU_CO ;
    wire \c0.n17192_THRU_CRY_1_THRU_CO ;
    wire \c0.n17192_THRU_CRY_2_THRU_CO ;
    wire \c0.n17192_THRU_CRY_3_THRU_CO ;
    wire \c0.n17192_THRU_CRY_4_THRU_CO ;
    wire \c0.n17192_THRU_CRY_5_THRU_CO ;
    wire \c0.n17192_THRU_CRY_6_THRU_CO ;
    wire bfn_14_18_0_;
    wire \c0.n6_adj_3188 ;
    wire \c0.n17193 ;
    wire \c0.n17193_THRU_CRY_0_THRU_CO ;
    wire \c0.n17193_THRU_CRY_1_THRU_CO ;
    wire \c0.n17193_THRU_CRY_2_THRU_CO ;
    wire \c0.n17193_THRU_CRY_3_THRU_CO ;
    wire \c0.n17193_THRU_CRY_4_THRU_CO ;
    wire \c0.n17193_THRU_CRY_5_THRU_CO ;
    wire \c0.n17193_THRU_CRY_6_THRU_CO ;
    wire bfn_14_19_0_;
    wire \c0.n6_adj_3186 ;
    wire \c0.n17194 ;
    wire \c0.n17194_THRU_CRY_0_THRU_CO ;
    wire \c0.n17194_THRU_CRY_1_THRU_CO ;
    wire \c0.n17194_THRU_CRY_2_THRU_CO ;
    wire \c0.n17194_THRU_CRY_3_THRU_CO ;
    wire \c0.n17194_THRU_CRY_4_THRU_CO ;
    wire \c0.n17194_THRU_CRY_5_THRU_CO ;
    wire \c0.n17194_THRU_CRY_6_THRU_CO ;
    wire bfn_14_20_0_;
    wire \c0.n6_adj_3184 ;
    wire \c0.n17195 ;
    wire \c0.n17195_THRU_CRY_0_THRU_CO ;
    wire \c0.n17195_THRU_CRY_1_THRU_CO ;
    wire \c0.n17195_THRU_CRY_2_THRU_CO ;
    wire \c0.n17195_THRU_CRY_3_THRU_CO ;
    wire \c0.n17195_THRU_CRY_4_THRU_CO ;
    wire \c0.n17195_THRU_CRY_5_THRU_CO ;
    wire \c0.n17195_THRU_CRY_6_THRU_CO ;
    wire bfn_14_21_0_;
    wire \c0.n6_adj_3182 ;
    wire \c0.n17196 ;
    wire \c0.n17196_THRU_CRY_0_THRU_CO ;
    wire \c0.n17196_THRU_CRY_1_THRU_CO ;
    wire \c0.n17196_THRU_CRY_2_THRU_CO ;
    wire \c0.n17196_THRU_CRY_3_THRU_CO ;
    wire \c0.n17196_THRU_CRY_4_THRU_CO ;
    wire \c0.n17196_THRU_CRY_5_THRU_CO ;
    wire \c0.n17196_THRU_CRY_6_THRU_CO ;
    wire bfn_14_22_0_;
    wire \c0.n6_adj_3180 ;
    wire \c0.n17197 ;
    wire \c0.n17197_THRU_CRY_0_THRU_CO ;
    wire \c0.n17197_THRU_CRY_1_THRU_CO ;
    wire \c0.n17197_THRU_CRY_2_THRU_CO ;
    wire \c0.n17197_THRU_CRY_3_THRU_CO ;
    wire \c0.n17197_THRU_CRY_4_THRU_CO ;
    wire \c0.n17197_THRU_CRY_5_THRU_CO ;
    wire \c0.n17197_THRU_CRY_6_THRU_CO ;
    wire bfn_14_23_0_;
    wire \c0.n6_adj_3178 ;
    wire \c0.n17198 ;
    wire \c0.n17198_THRU_CRY_0_THRU_CO ;
    wire \c0.n17198_THRU_CRY_1_THRU_CO ;
    wire \c0.n17198_THRU_CRY_2_THRU_CO ;
    wire \c0.n17198_THRU_CRY_3_THRU_CO ;
    wire \c0.n17198_THRU_CRY_4_THRU_CO ;
    wire \c0.n17198_THRU_CRY_5_THRU_CO ;
    wire \c0.n17198_THRU_CRY_6_THRU_CO ;
    wire bfn_14_24_0_;
    wire \c0.n17199 ;
    wire \c0.n17199_THRU_CRY_0_THRU_CO ;
    wire \c0.n17199_THRU_CRY_1_THRU_CO ;
    wire \c0.n17199_THRU_CRY_2_THRU_CO ;
    wire \c0.n17199_THRU_CRY_3_THRU_CO ;
    wire \c0.n17199_THRU_CRY_4_THRU_CO ;
    wire \c0.n17199_THRU_CRY_5_THRU_CO ;
    wire \c0.n17199_THRU_CRY_6_THRU_CO ;
    wire bfn_14_25_0_;
    wire \c0.n17200 ;
    wire \c0.n17200_THRU_CRY_0_THRU_CO ;
    wire \c0.n17200_THRU_CRY_1_THRU_CO ;
    wire \c0.n17200_THRU_CRY_2_THRU_CO ;
    wire \c0.n17200_THRU_CRY_3_THRU_CO ;
    wire \c0.n17200_THRU_CRY_4_THRU_CO ;
    wire \c0.n17200_THRU_CRY_5_THRU_CO ;
    wire \c0.n17200_THRU_CRY_6_THRU_CO ;
    wire bfn_14_26_0_;
    wire \c0.n17201 ;
    wire \c0.n17201_THRU_CRY_0_THRU_CO ;
    wire \c0.n17201_THRU_CRY_1_THRU_CO ;
    wire \c0.n17201_THRU_CRY_2_THRU_CO ;
    wire \c0.n17201_THRU_CRY_3_THRU_CO ;
    wire \c0.n17201_THRU_CRY_4_THRU_CO ;
    wire \c0.n17201_THRU_CRY_5_THRU_CO ;
    wire \c0.n17201_THRU_CRY_6_THRU_CO ;
    wire bfn_14_27_0_;
    wire \c0.n17202 ;
    wire \c0.n17202_THRU_CRY_0_THRU_CO ;
    wire \c0.n17202_THRU_CRY_1_THRU_CO ;
    wire \c0.n17202_THRU_CRY_2_THRU_CO ;
    wire \c0.n17202_THRU_CRY_3_THRU_CO ;
    wire \c0.n17202_THRU_CRY_4_THRU_CO ;
    wire \c0.n17202_THRU_CRY_5_THRU_CO ;
    wire \c0.n17202_THRU_CRY_6_THRU_CO ;
    wire bfn_14_28_0_;
    wire \c0.n17203 ;
    wire \c0.n17203_THRU_CRY_0_THRU_CO ;
    wire \c0.n17203_THRU_CRY_1_THRU_CO ;
    wire \c0.n17203_THRU_CRY_2_THRU_CO ;
    wire \c0.n17203_THRU_CRY_3_THRU_CO ;
    wire \c0.n17203_THRU_CRY_4_THRU_CO ;
    wire \c0.n17203_THRU_CRY_5_THRU_CO ;
    wire \c0.n17203_THRU_CRY_6_THRU_CO ;
    wire bfn_14_29_0_;
    wire \c0.n17204 ;
    wire \c0.n17204_THRU_CRY_0_THRU_CO ;
    wire \c0.n17204_THRU_CRY_1_THRU_CO ;
    wire \c0.n17204_THRU_CRY_2_THRU_CO ;
    wire \c0.n17204_THRU_CRY_3_THRU_CO ;
    wire \c0.n17204_THRU_CRY_4_THRU_CO ;
    wire \c0.n17204_THRU_CRY_5_THRU_CO ;
    wire \c0.n17204_THRU_CRY_6_THRU_CO ;
    wire bfn_14_30_0_;
    wire \c0.n17205 ;
    wire \c0.n17205_THRU_CRY_0_THRU_CO ;
    wire \c0.n17205_THRU_CRY_1_THRU_CO ;
    wire \c0.n17205_THRU_CRY_2_THRU_CO ;
    wire \c0.n17205_THRU_CRY_3_THRU_CO ;
    wire \c0.n17205_THRU_CRY_4_THRU_CO ;
    wire \c0.n17205_THRU_CRY_5_THRU_CO ;
    wire \c0.n17205_THRU_CRY_6_THRU_CO ;
    wire bfn_14_31_0_;
    wire \c0.n17206 ;
    wire \c0.n17206_THRU_CRY_0_THRU_CO ;
    wire \c0.n17206_THRU_CRY_1_THRU_CO ;
    wire \c0.n17206_THRU_CRY_2_THRU_CO ;
    wire \c0.n17206_THRU_CRY_3_THRU_CO ;
    wire \c0.n17206_THRU_CRY_4_THRU_CO ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \c0.n17206_THRU_CRY_5_THRU_CO ;
    wire \c0.n17206_THRU_CRY_6_THRU_CO ;
    wire bfn_14_32_0_;
    wire n20764;
    wire n16;
    wire \c0.n6_adj_3155 ;
    wire encoder0_position_24;
    wire n2340;
    wire encoder1_position_5;
    wire \c0.n21647 ;
    wire encoder1_position_26;
    wire data_out_frame_10_2;
    wire \c0.n6_adj_3154 ;
    wire data_out_frame_6_0;
    wire \c0.n6_adj_3321 ;
    wire n2344;
    wire data_out_frame_28_4;
    wire n2342;
    wire encoder1_position_3;
    wire encoder0_position_19;
    wire \c0.n6_adj_3379_cascade_ ;
    wire n2324;
    wire encoder1_position_21;
    wire \c0.n21559 ;
    wire \c0.n5_adj_3102 ;
    wire n2322;
    wire encoder0_position_11;
    wire data_out_frame_10_7;
    wire \c0.n21623 ;
    wire data_out_frame_9_3;
    wire \c0.n21641 ;
    wire data_out_frame_8_3;
    wire \c0.n21644 ;
    wire data_out_frame_11_5;
    wire data_out_frame_8_5;
    wire \c0.n21635_cascade_ ;
    wire data_out_frame_9_5;
    wire data_out_frame_5_3;
    wire \c0.n21470 ;
    wire \c0.n21542 ;
    wire n2316;
    wire \c0.n6_adj_3156 ;
    wire encoder1_position_29;
    wire data_out_frame_10_5;
    wire encoder0_position_29;
    wire \c0.data_out_frame_7_0 ;
    wire \c0.n17150 ;
    wire encoder1_position_18;
    wire data_out_frame_11_2;
    wire data_out_frame_10_0;
    wire data_out_frame_11_0;
    wire data_out_frame_8_0;
    wire \c0.n21617_cascade_ ;
    wire data_out_frame_9_0;
    wire \c0.n21620_cascade_ ;
    wire \c0.n21574 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n7235 ;
    wire \c0.n2_adj_3147 ;
    wire \c0.n6_adj_3151 ;
    wire encoder0_position_21;
    wire r_Tx_Data_7;
    wire data_out_frame_7_5;
    wire data_out_frame_6_5;
    wire \c0.n5_adj_3447 ;
    wire byte_transmit_counter_5;
    wire n9377;
    wire data_out_frame_5_5;
    wire \c0.n21546 ;
    wire \c0.n6_adj_3192 ;
    wire encoder1_position_1;
    wire data_out_frame_13_1;
    wire \c0.n6_adj_3190 ;
    wire \c0.rx.n14601_cascade_ ;
    wire n12301;
    wire \c0.n15685 ;
    wire \c0.rx.n6 ;
    wire n12492_cascade_;
    wire \c0.r_Bit_Index_0 ;
    wire tx_o;
    wire r_Tx_Data_1;
    wire \c0.r_SM_Main_2 ;
    wire \c0.n21611 ;
    wire encoder0_position_23;
    wire data_out_frame_7_7;
    wire n13179;
    wire bfn_15_19_0_;
    wire \c0.rx.n17267 ;
    wire n12908;
    wire \c0.rx.n17268 ;
    wire \c0.rx.n17269 ;
    wire \c0.rx.n17270 ;
    wire \c0.rx.n17271 ;
    wire \c0.rx.n17272 ;
    wire \c0.rx.n3 ;
    wire \c0.rx.n17273 ;
    wire \c0.rx.n7 ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire \c0.n6_adj_3161 ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire \c0.n6_adj_3172 ;
    wire \c0.n6_adj_3194 ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire \c0.n6_adj_3160 ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire \c0.n41_adj_3258_cascade_ ;
    wire \c0.n43_adj_3257 ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire \c0.n40_adj_3259 ;
    wire \c0.n45_adj_3262 ;
    wire \c0.n39_adj_3260_cascade_ ;
    wire \c0.n50_adj_3261 ;
    wire \c0.n11432 ;
    wire \c0.n14_adj_3080_cascade_ ;
    wire \c0.n10_adj_3081 ;
    wire \c0.n4812 ;
    wire \c0.n19119 ;
    wire \c0.n19119_cascade_ ;
    wire \c0.n21273 ;
    wire \c0.n5_adj_3306_cascade_ ;
    wire \c0.n2_adj_3302 ;
    wire \c0.n11433_cascade_ ;
    wire \c0.n8_adj_3228_cascade_ ;
    wire \c0.n2103 ;
    wire \c0.n2103_cascade_ ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n18653 ;
    wire \c0.FRAME_MATCHER_state_31_N_1736_2 ;
    wire \c0.FRAME_MATCHER_state_31_N_1736_1 ;
    wire \c0.n6_adj_3176 ;
    wire \c0.n11433 ;
    wire \c0.n700 ;
    wire \c0.n1 ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire \c0.n44_adj_3255 ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire \c0.n6_adj_3174 ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n18675 ;
    wire n11289;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire n2108_cascade_;
    wire \c0.n6_adj_3170 ;
    wire \c0.n6_adj_3165 ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire \c0.n6_adj_3168 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.n6_adj_3166 ;
    wire \c0.n6_adj_3159 ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire \c0.n6_adj_3164 ;
    wire \c0.n6_adj_3150 ;
    wire n2333;
    wire \c0.n21319 ;
    wire encoder0_position_18;
    wire \c0.n21317 ;
    wire count_enable;
    wire n2252;
    wire encoder0_position_27;
    wire data_out_frame_7_3;
    wire data_out_frame_6_3;
    wire \c0.n5_adj_3380 ;
    wire \c0.n21320 ;
    wire \c0.n21562 ;
    wire \c0.n21322_cascade_ ;
    wire n10_adj_3594;
    wire data_out_frame_7_2;
    wire \c0.n5_adj_3106 ;
    wire encoder0_position_26;
    wire data_out_frame_6_2;
    wire \c0.data_out_frame_0_2 ;
    wire \c0.n21473_cascade_ ;
    wire \c0.n6_adj_3105 ;
    wire data_out_frame_28_6;
    wire \c0.data_out_frame_0_3 ;
    wire \c0.n11_adj_3325 ;
    wire encoder1_position_8;
    wire data_out_frame_12_0;
    wire encoder1_position_23;
    wire data_out_frame_11_7;
    wire n2317;
    wire count_enable_adj_3586;
    wire encoder1_position_28;
    wire data_out_frame_5_6;
    wire data_out_frame_29_3;
    wire \c0.data_out_frame_28_3 ;
    wire \c0.n9753 ;
    wire \c0.n26_adj_3382_cascade_ ;
    wire \c0.n21314 ;
    wire \c0.n21316 ;
    wire data_out_frame_5_4;
    wire \c0.n21465 ;
    wire \c0.data_out_frame_5_0 ;
    wire control_mode_5;
    wire \c0.n21638 ;
    wire \c0.n11_adj_3462 ;
    wire data_out_frame_5_2;
    wire \c0.rx.n9 ;
    wire n12920;
    wire \c0.n70 ;
    wire \c0.n15850 ;
    wire \c0.n21231 ;
    wire \c0.n12254 ;
    wire encoder1_position_12;
    wire data_out_frame_12_4;
    wire data_out_frame_5_7;
    wire \c0.n5_adj_3475 ;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.n21576_cascade_ ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n21302_cascade_ ;
    wire \c0.n21304_cascade_ ;
    wire \c0.n21572 ;
    wire n9;
    wire \c0.n9755 ;
    wire data_out_frame_28_5;
    wire \c0.n21308 ;
    wire byte_transmit_counter_4;
    wire byte_transmit_counter_3;
    wire \c0.n21310_cascade_ ;
    wire \c0.n21568 ;
    wire n9_adj_3590;
    wire \c0.rx.n11302 ;
    wire \c0.rx.n11302_cascade_ ;
    wire encoder1_position_0;
    wire data_out_frame_13_0;
    wire \c0.rx.n21451_cascade_ ;
    wire \c0.rx.n15906_cascade_ ;
    wire \c0.rx.n20851 ;
    wire \c0.rx.n32 ;
    wire \c0.rx.n20964 ;
    wire \c0.rx.n15906 ;
    wire r_SM_Main_2_N_2473_2_cascade_;
    wire \c0.rx.n15926 ;
    wire \c0.rx.n35_cascade_ ;
    wire r_SM_Main_0;
    wire \c0.rx.n12_cascade_ ;
    wire r_SM_Main_1;
    wire r_SM_Main_2;
    wire \c0.rx.n21406_cascade_ ;
    wire r_SM_Main_2_N_2473_2;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.r_Clock_Count_0 ;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n8 ;
    wire n12914;
    wire n12917;
    wire \c0.n11440 ;
    wire \c0.n11317_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n21267 ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire \c0.n42_adj_3256 ;
    wire \c0.n1_adj_3002 ;
    wire \c0.n21053 ;
    wire \c0.n11_adj_3093 ;
    wire \c0.n15701_cascade_ ;
    wire n11421_cascade_;
    wire \c0.n11422 ;
    wire \c0.n3632 ;
    wire \c0.n9389 ;
    wire \c0.n3 ;
    wire \c0.n11427 ;
    wire \c0.n15874 ;
    wire \c0.n121 ;
    wire \c0.n103 ;
    wire \c0.n63_adj_3084 ;
    wire \c0.n19_adj_3252 ;
    wire \c0.n21_adj_3253 ;
    wire \c0.n19_adj_3252_cascade_ ;
    wire \c0.n63_adj_3083 ;
    wire \c0.n7804 ;
    wire \c0.n21281_cascade_ ;
    wire \c0.n108 ;
    wire \c0.n108_cascade_ ;
    wire \c0.n92_adj_3254 ;
    wire data_in_1_2;
    wire \c0.n26_adj_3107 ;
    wire \c0.n38_adj_3328 ;
    wire \c0.n21279_cascade_ ;
    wire \c0.n21255_cascade_ ;
    wire \c0.n37_adj_3332 ;
    wire \c0.n63_adj_3417_cascade_ ;
    wire \c0.n5_adj_3040_cascade_ ;
    wire \c0.n30_adj_3264 ;
    wire \c0.data_in_frame_5_0 ;
    wire \c0.data_in_frame_9_7 ;
    wire \c0.n19115_cascade_ ;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.n63_adj_3146 ;
    wire \c0.n20_adj_3437_cascade_ ;
    wire n21222_cascade_;
    wire control_mode_6;
    wire control_mode_2;
    wire control_mode_4;
    wire control_mode_3;
    wire control_mode_7;
    wire \c0.n9_cascade_ ;
    wire \c0.n16_adj_3008_cascade_ ;
    wire \c0.n9 ;
    wire \c0.n19449_cascade_ ;
    wire control_mode_0;
    wire FRAME_MATCHER_state_31_N_1800_2;
    wire FRAME_MATCHER_state_2;
    wire \c0.n15499 ;
    wire \c0.n13_adj_3016 ;
    wire \c0.FRAME_MATCHER_rx_data_ready_prev ;
    wire \c0.n19111_cascade_ ;
    wire \c0.n19493 ;
    wire \c0.n16 ;
    wire \c0.n24 ;
    wire \c0.n28_cascade_ ;
    wire \c0.n12026_cascade_ ;
    wire \c0.n10_cascade_ ;
    wire \c0.n21104 ;
    wire n3846_cascade_;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.n6_adj_2995 ;
    wire \c0.rx.n11455 ;
    wire \c0.rx.r_SM_Main_2_N_2479_0 ;
    wire n3792;
    wire n12911;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n15860 ;
    wire \c0.n19449 ;
    wire n12492;
    wire n12835;
    wire r_Bit_Index_0;
    wire \c0.n22_adj_3276_cascade_ ;
    wire \c0.n36_adj_3277_cascade_ ;
    wire \c0.n20415_cascade_ ;
    wire \c0.n14_adj_3407_cascade_ ;
    wire \c0.n100_adj_3403 ;
    wire \c0.n18_adj_3412 ;
    wire \c0.n20300_cascade_ ;
    wire \c0.n20300 ;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n3235 ;
    wire \c0.data_in_frame_28_6 ;
    wire \c0.n17947_cascade_ ;
    wire \c0.n20793 ;
    wire \c0.n10_adj_3242_cascade_ ;
    wire data_in_0_2;
    wire \c0.n14_adj_3243 ;
    wire \c0.n105 ;
    wire data_in_3_3;
    wire data_in_3_1;
    wire data_in_0_7;
    wire data_in_1_6;
    wire \c0.n18_adj_3229 ;
    wire \c0.n11446 ;
    wire \c0.n21108_cascade_ ;
    wire \c0.n12_adj_3248 ;
    wire data_in_3_5;
    wire \c0.n20_adj_3250 ;
    wire data_in_2_3;
    wire data_in_1_3;
    wire data_in_0_6;
    wire data_in_0_3;
    wire \c0.n18_adj_3246 ;
    wire \c0.n20_cascade_ ;
    wire \c0.n16_adj_3247 ;
    wire \c0.n11311 ;
    wire data_in_3_2;
    wire data_in_0_5;
    wire \c0.n5_adj_2999 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.n18655 ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.n20224_cascade_ ;
    wire \c0.n19_cascade_ ;
    wire \c0.n20246_cascade_ ;
    wire \c0.n24_adj_3327 ;
    wire \c0.n23_adj_3039_cascade_ ;
    wire \c0.n23_adj_3039 ;
    wire \c0.n30_adj_3042 ;
    wire data_out_frame_29_2;
    wire \c0.n18428_cascade_ ;
    wire \c0.n29_adj_3446 ;
    wire data_out_frame_28_2;
    wire \c0.data_out_frame_28__0__N_708_cascade_ ;
    wire \c0.data_out_frame_28__0__N_708 ;
    wire \c0.data_out_frame_29_0 ;
    wire \c0.data_out_frame_29_1 ;
    wire data_out_frame_28_1;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n26_adj_3103 ;
    wire \c0.n20209 ;
    wire \c0.n20204 ;
    wire \c0.n19217_cascade_ ;
    wire \c0.n66 ;
    wire n21222;
    wire control_mode_1;
    wire \c0.n16_adj_3018 ;
    wire \c0.n32_adj_3493_cascade_ ;
    wire \c0.n36_adj_3547_cascade_ ;
    wire \c0.n63_adj_3417 ;
    wire \c0.n38_adj_3548_cascade_ ;
    wire \c0.n34_adj_3411 ;
    wire \c0.n18443_cascade_ ;
    wire \c0.n25_adj_3495 ;
    wire \c0.data_in_frame_9_4 ;
    wire \c0.n25_adj_3495_cascade_ ;
    wire \c0.n6_adj_3005 ;
    wire \c0.n13 ;
    wire \c0.n20_adj_3539 ;
    wire \c0.n12_adj_3001_cascade_ ;
    wire \c0.n20403_cascade_ ;
    wire \c0.n10_adj_3514 ;
    wire \c0.n20398_cascade_ ;
    wire \c0.n4_adj_3071 ;
    wire \c0.n5_adj_3003 ;
    wire \c0.n36_adj_3267_cascade_ ;
    wire \c0.n94 ;
    wire \c0.n12_adj_3004 ;
    wire data_in_frame_18_6;
    wire n4_adj_3595;
    wire \c0.n14_adj_3434 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n14 ;
    wire \c0.n18667 ;
    wire \c0.n61_cascade_ ;
    wire \c0.n50 ;
    wire \c0.n61 ;
    wire \c0.n86_adj_3393_cascade_ ;
    wire \c0.n95_cascade_ ;
    wire \c0.n15_adj_3441 ;
    wire data_in_3_7;
    wire data_in_frame_16_6;
    wire \c0.data_in_frame_28_4 ;
    wire \c0.n20931 ;
    wire \c0.n18537 ;
    wire \c0.n20370 ;
    wire \c0.data_in_frame_29_7 ;
    wire \c0.data_in_frame_29_6 ;
    wire \c0.n10_adj_3152_cascade_ ;
    wire \c0.n21117 ;
    wire \c0.data_in_frame_29_0 ;
    wire \c0.n21117_cascade_ ;
    wire \c0.n18 ;
    wire \c0.n5_adj_3142 ;
    wire \c0.n5_adj_3142_cascade_ ;
    wire \c0.n22_adj_3305_cascade_ ;
    wire \c0.n37_adj_3309_cascade_ ;
    wire \c0.n21099_cascade_ ;
    wire \c0.n18_adj_3314 ;
    wire \c0.n10_adj_3353_cascade_ ;
    wire \c0.n21111 ;
    wire \c0.n9_adj_3352_cascade_ ;
    wire \c0.n21051 ;
    wire \c0.data_in_frame_27_7 ;
    wire \c0.data_in_frame_27_6 ;
    wire \c0.data_in_frame_26_4 ;
    wire data_in_2_2;
    wire \c0.n10_adj_3238 ;
    wire \c0.n110 ;
    wire data_in_2_5;
    wire data_in_1_5;
    wire \c0.n160 ;
    wire data_in_2_0;
    wire data_in_1_0;
    wire \c0.n12_adj_3230 ;
    wire data_in_2_7;
    wire \c0.n11443 ;
    wire data_in_0_1;
    wire FRAME_MATCHER_state_1;
    wire n4_adj_3596;
    wire n11421;
    wire n1295;
    wire \c0.n26 ;
    wire \c0.n5_adj_3044 ;
    wire \c0.n25_adj_3045 ;
    wire \c0.n14_adj_3073_cascade_ ;
    wire \c0.n10_adj_3068 ;
    wire \c0.n22_adj_3041 ;
    wire \c0.n21079 ;
    wire \c0.n11516 ;
    wire \c0.n14_adj_3480 ;
    wire \c0.n13_adj_3490_cascade_ ;
    wire \c0.n13_adj_3546 ;
    wire \c0.n15497 ;
    wire \c0.n14_adj_3459 ;
    wire \c0.n6_adj_3453 ;
    wire \c0.n39_adj_3398_cascade_ ;
    wire \c0.n13_adj_3526 ;
    wire \c0.n14_adj_3525 ;
    wire \c0.n15_adj_3543 ;
    wire \c0.n13_adj_3526_cascade_ ;
    wire \c0.n11_adj_3394 ;
    wire \c0.n28_adj_3519 ;
    wire \c0.n16_adj_3416_cascade_ ;
    wire \c0.n16_adj_3542 ;
    wire \c0.n5_adj_3528 ;
    wire \c0.n78_cascade_ ;
    wire \c0.n30_adj_3119_cascade_ ;
    wire \c0.n20088 ;
    wire \c0.n20055_cascade_ ;
    wire \c0.n5_adj_3099 ;
    wire \c0.n37_adj_3110_cascade_ ;
    wire \c0.n22_adj_3115 ;
    wire \c0.n6_adj_3024_cascade_ ;
    wire \c0.n18435_cascade_ ;
    wire \c0.data_in_frame_10_2 ;
    wire \c0.n14_adj_3007 ;
    wire \c0.n31_adj_3121 ;
    wire \c0.n27 ;
    wire \c0.n28_adj_3120_cascade_ ;
    wire \c0.n33_adj_3122 ;
    wire \c0.n20052_cascade_ ;
    wire \c0.n10_adj_3129_cascade_ ;
    wire \c0.n18400_cascade_ ;
    wire \c0.n5_adj_3040 ;
    wire \c0.n42_adj_3560 ;
    wire \c0.n35_adj_3342_cascade_ ;
    wire \c0.n39_adj_3339 ;
    wire \c0.n12_adj_3015 ;
    wire \c0.n44_adj_3561_cascade_ ;
    wire \c0.n13_adj_3017 ;
    wire \c0.n21118 ;
    wire data_in_frame_18_2;
    wire \c0.n21118_cascade_ ;
    wire \c0.n13_adj_3139 ;
    wire \c0.n36_adj_3267 ;
    wire \c0.n96_adj_3418_cascade_ ;
    wire \c0.n99_adj_3424 ;
    wire \c0.n77_adj_3415 ;
    wire \c0.n20801_cascade_ ;
    wire \c0.n96_adj_3401_cascade_ ;
    wire \c0.n99 ;
    wire \c0.n47_adj_3408 ;
    wire \c0.n18435 ;
    wire \c0.n42_adj_3064_cascade_ ;
    wire \c0.n15489_cascade_ ;
    wire \c0.data_in_frame_15_2 ;
    wire encoder0_position_31;
    wire data_out_frame_6_7;
    wire data_in_frame_23_2;
    wire \c0.n13_adj_3405_cascade_ ;
    wire \c0.data_in_frame_27_0 ;
    wire \c0.n17880_cascade_ ;
    wire \c0.n19342_cascade_ ;
    wire \c0.n12035 ;
    wire \c0.n19496_cascade_ ;
    wire \c0.n15_adj_3395 ;
    wire \c0.n19342 ;
    wire \c0.n36_adj_3307_cascade_ ;
    wire \c0.n39_adj_3312 ;
    wire \c0.n29_adj_3148 ;
    wire \c0.n78_adj_3357 ;
    wire \c0.n75_cascade_ ;
    wire \c0.n93_adj_3373_cascade_ ;
    wire \c0.n96_adj_3419 ;
    wire \c0.n23_adj_3222_cascade_ ;
    wire \c0.n76 ;
    wire \c0.n34 ;
    wire \c0.n19403 ;
    wire \c0.data_in_frame_26_6 ;
    wire \c0.n38_adj_3051 ;
    wire \c0.n38_adj_3051_cascade_ ;
    wire \c0.n19496 ;
    wire \c0.n17947 ;
    wire \c0.n60_adj_3065 ;
    wire \c0.n64 ;
    wire \c0.n51_cascade_ ;
    wire \c0.n32_adj_3052 ;
    wire \c0.n45_adj_3284 ;
    wire \c0.n40_adj_3282 ;
    wire \c0.n20930 ;
    wire \c0.n15_adj_3297_cascade_ ;
    wire \c0.n21003 ;
    wire \c0.n21_adj_3300_cascade_ ;
    wire \c0.n23_adj_3304 ;
    wire \c0.n21247_cascade_ ;
    wire \c0.n24_adj_3298 ;
    wire \c0.n14_adj_3354 ;
    wire data_in_3_4;
    wire data_in_0_0;
    wire data_in_1_7;
    wire \c0.n10_adj_3231 ;
    wire data_in_2_1;
    wire data_in_1_1;
    wire r_Bit_Index_2;
    wire r_Bit_Index_1;
    wire n4;
    wire n4_adj_3579;
    wire \c0.n9_adj_3025 ;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.n9_adj_3351 ;
    wire \c0.data_in_frame_4_6 ;
    wire \c0.n11_adj_3507 ;
    wire \c0.n13_adj_3504 ;
    wire \c0.n12131_cascade_ ;
    wire \c0.n12131 ;
    wire \c0.n19415 ;
    wire \c0.n19415_cascade_ ;
    wire \c0.n54_adj_3502 ;
    wire \c0.n39_adj_3398 ;
    wire \c0.n14_adj_3371 ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.n10_adj_3538_cascade_ ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.n22_adj_3356_cascade_ ;
    wire \c0.n13_adj_3513 ;
    wire \c0.n23_adj_3021 ;
    wire \c0.n23_adj_3021_cascade_ ;
    wire \c0.n26_adj_3114_cascade_ ;
    wire \c0.n24_adj_3011 ;
    wire \c0.n22 ;
    wire \c0.n22_adj_3356 ;
    wire \c0.n22_adj_3022 ;
    wire \c0.data_in_frame_12_4 ;
    wire \c0.n18_adj_3372 ;
    wire \c0.n88 ;
    wire \c0.n33 ;
    wire \c0.n20029 ;
    wire \c0.n26_adj_3114 ;
    wire \c0.n30 ;
    wire \c0.n18422 ;
    wire \c0.n18422_cascade_ ;
    wire \c0.n19433_cascade_ ;
    wire \c0.data_in_frame_10_3 ;
    wire \c0.n11891_cascade_ ;
    wire \c0.n44_adj_3117 ;
    wire \c0.n43_adj_3116 ;
    wire \c0.n27_adj_3118_cascade_ ;
    wire \c0.n20052 ;
    wire \c0.data_in_frame_14_5 ;
    wire \c0.n11_adj_3340 ;
    wire \c0.n19916_cascade_ ;
    wire \c0.n18_adj_3369 ;
    wire \c0.n19477_cascade_ ;
    wire \c0.n12_adj_3348_cascade_ ;
    wire \c0.n21045_cascade_ ;
    wire \c0.n27_adj_3118 ;
    wire \c0.n19_adj_3303 ;
    wire \c0.n12 ;
    wire \c0.n12_adj_3477 ;
    wire \c0.data_in_frame_14_4 ;
    wire \c0.n21110_cascade_ ;
    wire \c0.n20246 ;
    wire \c0.data_in_frame_14_3 ;
    wire \c0.n67_adj_3063 ;
    wire \c0.n20490 ;
    wire \c0.n19433 ;
    wire \c0.n42_adj_3064 ;
    wire \c0.n12_adj_3518 ;
    wire \c0.n12_adj_3517_cascade_ ;
    wire data_in_frame_18_5;
    wire \c0.n21_adj_3337 ;
    wire \c0.n20_adj_3487 ;
    wire \c0.n20451_cascade_ ;
    wire \c0.n5_adj_3220 ;
    wire data_in_frame_18_1;
    wire \c0.n27_adj_3529_cascade_ ;
    wire \c0.n32_adj_3530_cascade_ ;
    wire \c0.n19244_cascade_ ;
    wire \c0.n85_adj_3074 ;
    wire \c0.n85_adj_3074_cascade_ ;
    wire \c0.n10_adj_3474 ;
    wire \c0.n20801 ;
    wire \c0.n49 ;
    wire \c0.n48_adj_3409 ;
    wire \c0.n22_adj_3287_cascade_ ;
    wire \c0.n39_adj_3050 ;
    wire \c0.n19384 ;
    wire \c0.n13_adj_3463 ;
    wire \c0.n10 ;
    wire \c0.n19384_cascade_ ;
    wire data_in_frame_16_5;
    wire data_in_frame_19_0;
    wire \c0.n9_adj_3430_cascade_ ;
    wire \c0.n10_adj_3445 ;
    wire \c0.n9_adj_3430 ;
    wire \c0.n14_adj_3421 ;
    wire \c0.n18433_cascade_ ;
    wire \c0.n19511 ;
    wire \c0.n19511_cascade_ ;
    wire \c0.n21110 ;
    wire \c0.n20_adj_3448 ;
    wire \c0.n20431 ;
    wire \c0.n64_adj_3512 ;
    wire data_in_frame_16_4;
    wire \c0.n7_adj_3440 ;
    wire \c0.data_in_frame_13_0 ;
    wire \c0.n11_adj_3219 ;
    wire \c0.n13_adj_3221 ;
    wire data_in_frame_23_3;
    wire \c0.n25_adj_3524 ;
    wire \c0.n21044_cascade_ ;
    wire \c0.data_in_frame_26_7 ;
    wire \c0.n16_adj_3109_cascade_ ;
    wire \c0.n21071 ;
    wire \c0.n20479 ;
    wire \c0.n77 ;
    wire \c0.n34_adj_3096 ;
    wire \c0.n32_adj_3095 ;
    wire \c0.n18457_cascade_ ;
    wire \c0.n23_adj_3222 ;
    wire \c0.n43_adj_3280_cascade_ ;
    wire \c0.n41_adj_3281 ;
    wire \c0.n50_adj_3283 ;
    wire \c0.n18457 ;
    wire \c0.n21076 ;
    wire \c0.n33_adj_3308 ;
    wire \c0.n18417 ;
    wire \c0.n18417_cascade_ ;
    wire \c0.n19_adj_3292 ;
    wire \c0.data_in_frame_29_4 ;
    wire \c0.data_in_frame_29_2 ;
    wire \c0.data_in_frame_29_1 ;
    wire \c0.data_in_frame_28_1 ;
    wire \c0.data_in_frame_28_0 ;
    wire \c0.n20324 ;
    wire \c0.n14_adj_3349 ;
    wire \c0.n7_adj_3078 ;
    wire \c0.n17880 ;
    wire \c0.n26_adj_3523 ;
    wire data_in_0_4;
    wire n20896;
    wire \c0.n12085 ;
    wire \c0.n11865 ;
    wire \c0.n12085_cascade_ ;
    wire \c0.n6495 ;
    wire data_in_2_4;
    wire data_in_1_4;
    wire \c0.n6_adj_3343 ;
    wire \c0.data_out_frame_28_7 ;
    wire n8112;
    wire \c0.data_in_frame_4_3 ;
    wire \c0.data_in_frame_4_2 ;
    wire \c0.data_in_frame_6_4 ;
    wire \c0.n13_adj_3496_cascade_ ;
    wire \c0.data_in_frame_2_2 ;
    wire data_in_frame_0_0;
    wire \c0.n19277 ;
    wire \c0.data_in_frame_2_0 ;
    wire \c0.n8_adj_3397 ;
    wire \c0.n11833_cascade_ ;
    wire \c0.n92_cascade_ ;
    wire \c0.n80 ;
    wire \c0.n19196 ;
    wire \c0.data_in_frame_4_5 ;
    wire \c0.n54 ;
    wire \c0.n90 ;
    wire \c0.n98 ;
    wire \c0.n21277 ;
    wire \c0.n4_adj_3406 ;
    wire \c0.n14_adj_3476_cascade_ ;
    wire \c0.data_in_frame_7_3 ;
    wire \c0.n19508 ;
    wire \c0.n10_adj_3538 ;
    wire \c0.n85 ;
    wire \c0.n37 ;
    wire \c0.n67_cascade_ ;
    wire \c0.n96 ;
    wire \c0.n83 ;
    wire \c0.n40_adj_3032 ;
    wire \c0.n100_cascade_ ;
    wire \c0.n102 ;
    wire \c0.n4_adj_3009 ;
    wire \c0.n21_adj_3010 ;
    wire \c0.n28_adj_3023 ;
    wire \c0.n17_adj_3508 ;
    wire \c0.n19966 ;
    wire \c0.n30_adj_3075 ;
    wire \c0.n32_adj_3077_cascade_ ;
    wire \c0.n19372 ;
    wire \c0.n21047_cascade_ ;
    wire \c0.n42_adj_3111 ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.n10_adj_3014_cascade_ ;
    wire \c0.n40 ;
    wire \c0.n16_adj_3218_cascade_ ;
    wire \c0.data_in_frame_12_2 ;
    wire \c0.n7_adj_3491 ;
    wire \c0.n30_adj_3531 ;
    wire \c0.n12_adj_3034 ;
    wire \c0.n31_adj_3532 ;
    wire \c0.n11537 ;
    wire \c0.data_in_frame_15_6 ;
    wire \c0.n16_adj_3481_cascade_ ;
    wire \c0.n11815_cascade_ ;
    wire \c0.n19291 ;
    wire data_in_frame_16_1;
    wire \c0.n12056_cascade_ ;
    wire \c0.n12_adj_3249 ;
    wire \c0.n12_adj_3249_cascade_ ;
    wire \c0.n12056 ;
    wire \c0.n19301 ;
    wire \c0.n19301_cascade_ ;
    wire \c0.n31_adj_3126_cascade_ ;
    wire \c0.n19427 ;
    wire \c0.n19551 ;
    wire \c0.n27_adj_3455 ;
    wire \c0.n46_cascade_ ;
    wire \c0.n46 ;
    wire \c0.n8 ;
    wire \c0.n84 ;
    wire \c0.n19824_cascade_ ;
    wire \c0.n29 ;
    wire \c0.n18_adj_3360_cascade_ ;
    wire \c0.n32_adj_3362_cascade_ ;
    wire \c0.n20112_cascade_ ;
    wire \c0.data_in_frame_13_1 ;
    wire \c0.n18398_cascade_ ;
    wire \c0.n37_adj_3390_cascade_ ;
    wire \c0.n37_adj_3390 ;
    wire \c0.n60_adj_3368_cascade_ ;
    wire \c0.n51_adj_3376 ;
    wire \c0.n19916 ;
    wire \c0.n18443 ;
    wire \c0.n39_adj_3334 ;
    wire \c0.n19_adj_3336 ;
    wire \c0.n39_adj_3334_cascade_ ;
    wire \c0.n25_adj_3431 ;
    wire \c0.n42_adj_3367 ;
    wire \c0.n43_adj_3386 ;
    wire \c0.n40_adj_3366 ;
    wire \c0.n30_adj_3429 ;
    wire \c0.n35_adj_3274_cascade_ ;
    wire \c0.n59 ;
    wire \c0.n30_adj_3392 ;
    wire \c0.n21047 ;
    wire \c0.n12_adj_3049 ;
    wire \c0.n91 ;
    wire \c0.n35_adj_3274 ;
    wire \c0.n17_adj_3451 ;
    wire \c0.n20403 ;
    wire \c0.n22_adj_3450 ;
    wire \c0.n24_adj_3427_cascade_ ;
    wire \c0.data_in_frame_17_0 ;
    wire \c0.n32_adj_3057_cascade_ ;
    wire \c0.n33_adj_3289 ;
    wire \c0.n10_adj_3555 ;
    wire \c0.n4_adj_3522 ;
    wire \c0.n55_adj_3273 ;
    wire \c0.n19514 ;
    wire \c0.n20965_cascade_ ;
    wire \c0.n40_adj_3323 ;
    wire \c0.data_in_frame_27_3 ;
    wire \c0.n20336_cascade_ ;
    wire \c0.n61_adj_3387 ;
    wire \c0.n63_adj_3391 ;
    wire \c0.n21034_cascade_ ;
    wire \c0.n12134 ;
    wire \c0.n58_adj_3381 ;
    wire \c0.n43_adj_3330 ;
    wire \c0.n50_adj_3331 ;
    wire \c0.n35_adj_3266 ;
    wire \c0.n33_adj_3097 ;
    wire \c0.n9_adj_3240 ;
    wire \c0.n20112 ;
    wire \c0.n32_adj_3236 ;
    wire \c0.n28_adj_3245 ;
    wire \c0.n27_adj_3241_cascade_ ;
    wire \c0.n13_adj_3244 ;
    wire \c0.n19_adj_3135 ;
    wire \c0.n19_adj_3135_cascade_ ;
    wire \c0.n24_adj_3134 ;
    wire \c0.n86 ;
    wire \c0.n22_adj_3136_cascade_ ;
    wire \c0.n11936_cascade_ ;
    wire \c0.data_in_frame_27_4 ;
    wire \c0.data_in_frame_27_5 ;
    wire \c0.n17_adj_3318 ;
    wire \c0.n11936 ;
    wire \c0.n12_adj_3141 ;
    wire data_in_frame_24_6;
    wire data_in_frame_24_4;
    wire \c0.n19465_cascade_ ;
    wire \c0.n17 ;
    wire \c0.n21044 ;
    wire \c0.n19703 ;
    wire \c0.n19703_cascade_ ;
    wire \c0.n44_adj_3278 ;
    wire \c0.data_in_frame_25_1 ;
    wire \c0.n18377 ;
    wire \c0.data_in_frame_25_2 ;
    wire \c0.data_in_frame_25_3 ;
    wire \c0.n19400 ;
    wire \c0.data_in_frame_26_5 ;
    wire \c0.n17840 ;
    wire data_in_3_0;
    wire \c0.n12_adj_3498 ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire \c0.n6_adj_3149 ;
    wire \c0.data_in_frame_8_6 ;
    wire \c0.data_in_frame_4_0 ;
    wire \c0.n17_adj_3113 ;
    wire \c0.n5_adj_3030 ;
    wire \c0.n60_cascade_ ;
    wire \c0.n93 ;
    wire \c0.data_in_frame_6_1 ;
    wire \c0.n5_adj_3028 ;
    wire \c0.n19443 ;
    wire \c0.n11687 ;
    wire \c0.n20313 ;
    wire \c0.n8_adj_3066_cascade_ ;
    wire \c0.n19170 ;
    wire \c0.n19170_cascade_ ;
    wire \c0.data_in_frame_8_2 ;
    wire \c0.n21_adj_3053 ;
    wire \c0.n21 ;
    wire \c0.data_in_frame_5_4 ;
    wire \c0.n25 ;
    wire \c0.n89 ;
    wire \c0.data_in_frame_3_1 ;
    wire data_in_frame_0_5;
    wire \c0.n33_adj_3088 ;
    wire \c0.n15_adj_3545 ;
    wire \c0.n24_adj_3013 ;
    wire \c0.data_in_frame_3_3 ;
    wire \c0.data_in_frame_3_2 ;
    wire data_out_frame_29__3__N_647;
    wire \c0.n29_adj_3216 ;
    wire \c0.n78 ;
    wire \c0.n37_adj_3215 ;
    wire \c0.n29_adj_3216_cascade_ ;
    wire \c0.n44_adj_3217 ;
    wire \c0.n36_adj_3212_cascade_ ;
    wire \c0.n41_adj_3213 ;
    wire \c0.n20340 ;
    wire \c0.n11651_cascade_ ;
    wire \c0.n27_adj_3082 ;
    wire \c0.n11800 ;
    wire \c0.n31 ;
    wire \c0.n37_adj_3153 ;
    wire \c0.n35_adj_3233 ;
    wire \c0.n60 ;
    wire \c0.n52_adj_3223_cascade_ ;
    wire \c0.n60_adj_3503 ;
    wire \c0.n52_adj_3402 ;
    wire \c0.data_in_frame_7_4 ;
    wire \c0.n20391 ;
    wire \c0.n4 ;
    wire \c0.n12026 ;
    wire \c0.n5 ;
    wire \c0.n4_cascade_ ;
    wire \c0.data_in_frame_11_4 ;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.data_in_frame_21_0 ;
    wire \c0.n16_adj_3218 ;
    wire \c0.n48 ;
    wire \c0.data_in_frame_5_1 ;
    wire \c0.n20224 ;
    wire \c0.n5_adj_3549 ;
    wire \c0.data_in_frame_4_7 ;
    wire \c0.n11613 ;
    wire \c0.data_in_frame_17_6 ;
    wire data_in_frame_18_0;
    wire \c0.n11613_cascade_ ;
    wire \c0.n19477 ;
    wire \c0.n17_adj_3482 ;
    wire \c0.data_in_frame_13_6 ;
    wire \c0.data_in_frame_13_5 ;
    wire \c0.n20826 ;
    wire \c0.n54_adj_3234 ;
    wire \c0.n43_adj_3232_cascade_ ;
    wire \c0.n17849 ;
    wire \c0.n49_adj_3237 ;
    wire \c0.n7_adj_3225_cascade_ ;
    wire \c0.data_in_frame_15_4 ;
    wire \c0.n7_adj_3225 ;
    wire \c0.n44_adj_3226 ;
    wire \c0.data_in_frame_10_4 ;
    wire \c0.data_in_frame_8_1 ;
    wire \c0.n41_adj_3365 ;
    wire \c0.n22_adj_3287 ;
    wire \c0.n47_adj_3286_cascade_ ;
    wire \c0.n51_adj_3290 ;
    wire \c0.n52_adj_3288_cascade_ ;
    wire \c0.n6_adj_3291 ;
    wire \c0.data_in_frame_11_6 ;
    wire \c0.n19909_cascade_ ;
    wire \c0.n87 ;
    wire \c0.n6_adj_3137 ;
    wire \c0.n35_adj_3098 ;
    wire \c0.n19909 ;
    wire \c0.n19223 ;
    wire \c0.n12218 ;
    wire \c0.n7_adj_3047_cascade_ ;
    wire \c0.n28_adj_3059_cascade_ ;
    wire \c0.n36_adj_3452 ;
    wire \c0.n47 ;
    wire \c0.n17819 ;
    wire \c0.n20321 ;
    wire \c0.n19824 ;
    wire \c0.n12_adj_3469 ;
    wire \c0.n29_adj_3461_cascade_ ;
    wire \c0.n25_adj_3035 ;
    wire \c0.n23_adj_3364 ;
    wire \c0.n24_adj_3335 ;
    wire \c0.n36_adj_3470_cascade_ ;
    wire \c0.n22_adj_3341 ;
    wire \c0.n11_adj_3124_cascade_ ;
    wire \c0.n32_adj_3465 ;
    wire \c0.n33_adj_3315 ;
    wire \c0.n49_adj_3316 ;
    wire \c0.n35_adj_3317 ;
    wire \c0.data_in_frame_17_1 ;
    wire \c0.n17871 ;
    wire \c0.n22_adj_3363 ;
    wire \c0.n22_adj_3363_cascade_ ;
    wire \c0.n30_adj_3468 ;
    wire \c0.n65 ;
    wire \c0.n70_adj_3087_cascade_ ;
    wire \c0.n20339 ;
    wire \c0.n27_adj_3311 ;
    wire \c0.n7_adj_3094 ;
    wire \c0.n20_adj_3293 ;
    wire \c0.n33_adj_3279 ;
    wire \c0.n30_adj_3295 ;
    wire \c0.n32_adj_3294_cascade_ ;
    wire \c0.n21075 ;
    wire \c0.n7_adj_3079 ;
    wire \c0.n29_adj_3299 ;
    wire \c0.n19_adj_3320 ;
    wire \c0.n20336 ;
    wire \c0.n18379 ;
    wire \c0.n21034 ;
    wire \c0.n57 ;
    wire \c0.n24_adj_3427 ;
    wire \c0.n11714 ;
    wire \c0.n22_adj_3296 ;
    wire \c0.n19159_cascade_ ;
    wire \c0.n11632 ;
    wire \c0.n19159 ;
    wire \c0.data_in_frame_28_7 ;
    wire \c0.n79 ;
    wire \c0.n10_adj_3207 ;
    wire \c0.n11_adj_3206 ;
    wire \c0.n11776_cascade_ ;
    wire \c0.n6_adj_3319 ;
    wire data_in_frame_24_7;
    wire \c0.n12206 ;
    wire \c0.n19268 ;
    wire \c0.n19268_cascade_ ;
    wire \c0.n20_adj_3301 ;
    wire \c0.n7_adj_3054 ;
    wire \c0.n11601 ;
    wire \c0.n19764 ;
    wire \c0.n42_adj_3055 ;
    wire \c0.n11815 ;
    wire \c0.n4_adj_3100 ;
    wire \c0.data_in_frame_25_0 ;
    wire \c0.n19436 ;
    wire data_in_frame_22_4;
    wire \c0.n19436_cascade_ ;
    wire \c0.n11776 ;
    wire \c0.n6_adj_3112 ;
    wire \c0.n19151 ;
    wire \c0.n20933 ;
    wire rx_data_ready;
    wire data_in_3_6;
    wire data_in_2_6;
    wire \c0.n25_adj_3048 ;
    wire \c0.n19312 ;
    wire \c0.n20512 ;
    wire \c0.n19202 ;
    wire \c0.n12_adj_3210_cascade_ ;
    wire \c0.n18433 ;
    wire \c0.n17834 ;
    wire \c0.n21767 ;
    wire data_in_frame_22_6;
    wire data_in_frame_23_0;
    wire data_in_frame_23_4;
    wire n19126;
    wire \c0.data_in_frame_11_0 ;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.n34_adj_3326 ;
    wire \c0.n13_adj_3344 ;
    wire \c0.n23_adj_3076 ;
    wire \c0.n19424 ;
    wire \c0.n7_adj_3029 ;
    wire data_in_frame_0_4;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.data_in_frame_4_4 ;
    wire \c0.n8_adj_3345 ;
    wire \c0.n7_adj_3520 ;
    wire \c0.n9_adj_3346 ;
    wire \c0.n8_adj_3345_cascade_ ;
    wire \c0.n11626_cascade_ ;
    wire \c0.data_in_frame_8_7 ;
    wire data_in_frame_1_1;
    wire \c0.n19970 ;
    wire \c0.n6_adj_3501 ;
    wire \c0.data_in_frame_6_3 ;
    wire \c0.n11478_cascade_ ;
    wire \c0.n81 ;
    wire data_in_frame_1_6;
    wire \c0.n11526 ;
    wire \c0.data_in_frame_6_5 ;
    wire \c0.n11549 ;
    wire \c0.n11651 ;
    wire \c0.n27_adj_3457 ;
    wire data_in_frame_1_7;
    wire \c0.n12_adj_3378 ;
    wire \c0.n11626 ;
    wire \c0.n21_adj_3205 ;
    wire \c0.n28_adj_3428 ;
    wire data_in_frame_1_5;
    wire \c0.n7_adj_3509 ;
    wire \c0.n7_adj_3509_cascade_ ;
    wire \c0.n10_adj_3012 ;
    wire \c0.n45 ;
    wire \c0.data_in_frame_4_1 ;
    wire data_in_frame_0_6;
    wire data_in_frame_1_0;
    wire \c0.n20341 ;
    wire \c0.n58_adj_3497 ;
    wire \c0.n56_adj_3505 ;
    wire \c0.n64_adj_3506 ;
    wire \c0.n19217 ;
    wire \c0.n4_adj_3036_cascade_ ;
    wire \c0.n57_adj_3499 ;
    wire \c0.n6_adj_3019 ;
    wire \c0.data_in_frame_7_5 ;
    wire \c0.n6_adj_3019_cascade_ ;
    wire \c0.n20386 ;
    wire \c0.data_in_frame_9_6 ;
    wire \c0.data_in_frame_3_7 ;
    wire \c0.data_in_frame_5_5 ;
    wire \c0.data_in_frame_5_3 ;
    wire n11461;
    wire \c0.n23 ;
    wire \c0.n51_adj_3426 ;
    wire n15645;
    wire r_Rx_Data;
    wire n11466;
    wire \c0.data_in_frame_13_7 ;
    wire \c0.n13_adj_3541 ;
    wire \c0.data_in_frame_13_2 ;
    wire \c0.data_in_frame_9_5 ;
    wire \c0.n9_adj_3211 ;
    wire data_in_frame_0_1;
    wire \c0.n17_adj_3544 ;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.n11858_cascade_ ;
    wire \c0.n19446 ;
    wire \c0.n19446_cascade_ ;
    wire \c0.data_out_frame_0__7__N_1537 ;
    wire \c0.n11982 ;
    wire \c0.n33_adj_3209_cascade_ ;
    wire \c0.n5598 ;
    wire \c0.data_in_frame_17_7 ;
    wire \c0.n9_adj_3350 ;
    wire \c0.n29_adj_3533 ;
    wire \c0.n33_adj_3209 ;
    wire \c0.n12209 ;
    wire \c0.n9_adj_3027 ;
    wire \c0.n45_adj_3224 ;
    wire \c0.data_in_frame_7_6 ;
    wire \c0.n15 ;
    wire \c0.n5753 ;
    wire \c0.data_in_frame_14_0 ;
    wire \c0.data_in_frame_12_0 ;
    wire \c0.n20055 ;
    wire \c0.n20_adj_3536_cascade_ ;
    wire \c0.n12_adj_3558_cascade_ ;
    wire \c0.data_in_frame_8_5 ;
    wire \c0.data_in_frame_12_7 ;
    wire \c0.n5_adj_3031 ;
    wire \c0.n19359_cascade_ ;
    wire \c0.data_in_frame_8_4 ;
    wire \c0.n11478 ;
    wire \c0.n19199 ;
    wire \c0.data_in_frame_10_5 ;
    wire \c0.n19199_cascade_ ;
    wire \c0.n19_adj_3540 ;
    wire \c0.data_in_frame_14_1 ;
    wire \c0.data_in_frame_15_7 ;
    wire \c0.data_in_frame_14_2 ;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.n20981 ;
    wire \c0.n25_adj_3157 ;
    wire \c0.n69 ;
    wire \c0.n28_adj_3059 ;
    wire \c0.n38_adj_3058_cascade_ ;
    wire \c0.n32_adj_3060 ;
    wire \c0.n8_adj_3061_cascade_ ;
    wire \c0.n52 ;
    wire \c0.n8_adj_3061 ;
    wire \c0.n43_adj_3285_cascade_ ;
    wire \c0.n53 ;
    wire \c0.n4_adj_3123 ;
    wire data_in_frame_16_7;
    wire \c0.data_in_frame_12_5 ;
    wire \c0.n12_adj_3554_cascade_ ;
    wire \c0.n20151 ;
    wire \c0.n20542 ;
    wire \c0.n20542_cascade_ ;
    wire \c0.n45_adj_3423 ;
    wire \c0.n25_adj_3510_cascade_ ;
    wire \c0.n58_adj_3511 ;
    wire \c0.n20085 ;
    wire \c0.n19244 ;
    wire \c0.n88_adj_3422 ;
    wire \c0.n25_adj_3510 ;
    wire \c0.n56 ;
    wire \c0.n44_adj_3125 ;
    wire \c0.n11_adj_3124 ;
    wire \c0.n48_adj_3313 ;
    wire \c0.n35_cascade_ ;
    wire \c0.n67_adj_3092 ;
    wire \c0.n43_adj_3089 ;
    wire \c0.n41_adj_3085 ;
    wire \c0.n42_adj_3086 ;
    wire \c0.n60_adj_3127 ;
    wire \c0.n55_adj_3128_cascade_ ;
    wire \c0.n19749 ;
    wire \c0.n58 ;
    wire \c0.n16_adj_3489 ;
    wire \c0.n31_adj_3126 ;
    wire \c0.n10_adj_3425_cascade_ ;
    wire \c0.n42_adj_3130 ;
    wire \c0.n92_adj_3272 ;
    wire \c0.n39_adj_3269 ;
    wire \c0.n36_adj_3275 ;
    wire \c0.n38_adj_3270 ;
    wire \c0.n39_adj_3269_cascade_ ;
    wire \c0.n37_adj_3268 ;
    wire \c0.n94_adj_3375 ;
    wire \c0.n92_adj_3377_cascade_ ;
    wire \c0.n91_adj_3389 ;
    wire \c0.n100_adj_3420 ;
    wire \c0.n11942 ;
    wire \c0.n12_adj_3208 ;
    wire \c0.n10_adj_3425 ;
    wire \c0.n82 ;
    wire \c0.n93_adj_3385 ;
    wire \c0.n32_adj_3057 ;
    wire \c0.n62 ;
    wire \c0.n68 ;
    wire \c0.n19502 ;
    wire \c0.n20_adj_3536 ;
    wire \c0.n23_adj_3534 ;
    wire \c0.n40_adj_3374 ;
    wire \c0.n38_adj_3062_cascade_ ;
    wire \c0.n39_adj_3384 ;
    wire \c0.n93_adj_3329 ;
    wire \c0.data_in_frame_8_3 ;
    wire \c0.n19505 ;
    wire \c0.n26_adj_3537 ;
    wire \c0.n20917_cascade_ ;
    wire \c0.n19524 ;
    wire \c0.n6_adj_3433_cascade_ ;
    wire \c0.n18375_cascade_ ;
    wire \c0.n38_adj_3062 ;
    wire \c0.n83_adj_3442 ;
    wire data_in_frame_18_7;
    wire \c0.n12052 ;
    wire \c0.n19_adj_3056 ;
    wire \c0.n19_adj_3056_cascade_ ;
    wire \c0.n21045 ;
    wire \c0.n29_adj_3454 ;
    wire \c0.n18398 ;
    wire \c0.n6_adj_3239 ;
    wire data_in_frame_22_2;
    wire \c0.n19354 ;
    wire data_in_frame_22_7;
    wire data_in_frame_22_3;
    wire data_in_frame_24_0;
    wire \c0.data_in_frame_26_2 ;
    wire \c0.n18431 ;
    wire \c0.n15701 ;
    wire \c0.n7_adj_3047 ;
    wire \c0.n20965 ;
    wire \c0.data_in_frame_26_0 ;
    wire \c0.data_in_frame_27_1 ;
    wire \c0.data_in_frame_27_2 ;
    wire \c0.data_in_frame_28_2 ;
    wire \c0.n20709 ;
    wire \c0.n17942 ;
    wire \c0.n77_adj_3396_cascade_ ;
    wire \c0.n90_adj_3400 ;
    wire \c0.data_in_frame_25_7 ;
    wire \c0.data_in_frame_25_5 ;
    wire \c0.data_in_frame_25_4 ;
    wire \c0.n19214_cascade_ ;
    wire data_in_frame_24_5;
    wire \c0.n12_adj_3214 ;
    wire \c0.data_in_frame_25_6 ;
    wire \c0.n5784 ;
    wire \c0.n11833 ;
    wire \c0.n19456 ;
    wire \c0.n5595 ;
    wire n2108;
    wire \c0.n6_adj_3140 ;
    wire \c0.data_in_frame_6_0 ;
    wire \c0.data_in_frame_6_2 ;
    wire data_in_frame_1_2;
    wire \c0.n9_adj_3101 ;
    wire FRAME_MATCHER_i_0;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire n19100;
    wire \c0.n20095 ;
    wire data_in_frame_0_3;
    wire \c0.n5240 ;
    wire \c0.n7_cascade_ ;
    wire \c0.n9_adj_3038 ;
    wire \c0.data_in_frame_6_7 ;
    wire \c0.n19098 ;
    wire \c0.n9_adj_3251 ;
    wire \c0.data_in_frame_3_4 ;
    wire \c0.n12_adj_2998 ;
    wire \c0.n19176 ;
    wire \c0.n11953 ;
    wire \c0.data_in_frame_5_2 ;
    wire data_in_frame_1_3;
    wire \c0.n55_adj_3500 ;
    wire data_in_frame_0_2;
    wire \c0.n7 ;
    wire \c0.n19241 ;
    wire \c0.data_in_frame_2_4 ;
    wire data_in_frame_1_4;
    wire \c0.n6_adj_3037 ;
    wire \c0.data_in_frame_5_7 ;
    wire \c0.n4_adj_3036 ;
    wire \c0.n6_adj_3037_cascade_ ;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.n19560 ;
    wire \c0.data_out_frame_0__7__N_1540 ;
    wire \c0.data_in_frame_6_6 ;
    wire \c0.n19258 ;
    wire \c0.data_in_frame_8_0 ;
    wire \c0.data_in_frame_7_7 ;
    wire \c0.data_in_frame_5_6 ;
    wire \c0.n8_adj_3020 ;
    wire \c0.data_in_frame_13_3 ;
    wire \c0.data_in_frame_9_2 ;
    wire \c0.n19115 ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.data_in_frame_11_5 ;
    wire \c0.n5_adj_3043 ;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.data_in_frame_9_0 ;
    wire \c0.data_in_frame_11_3 ;
    wire \c0.data_in_frame_13_4 ;
    wire \c0.n11_adj_3492 ;
    wire \c0.n11_adj_3492_cascade_ ;
    wire data_in_frame_16_0;
    wire \c0.n20_adj_3527 ;
    wire \c0.data_in_frame_11_1 ;
    wire \c0.n19229 ;
    wire \c0.data_in_frame_11_2 ;
    wire \c0.n19134 ;
    wire \c0.data_in_frame_10_7 ;
    wire \c0.n19131 ;
    wire \c0.data_in_frame_11_7 ;
    wire \c0.n15489 ;
    wire \c0.n19140 ;
    wire \c0.data_in_frame_15_5 ;
    wire \c0.n9_adj_3552_cascade_ ;
    wire data_in_frame_18_3;
    wire n19129;
    wire data_in_frame_18_4;
    wire \c0.data_in_frame_12_1 ;
    wire \c0.n7_adj_3000 ;
    wire \c0.n19430 ;
    wire \c0.n7_adj_3000_cascade_ ;
    wire data_in_frame_16_3;
    wire \c0.n6 ;
    wire \c0.n19187 ;
    wire \c0.n46_adj_3443 ;
    wire \c0.data_in_frame_15_0 ;
    wire \c0.n40_adj_3413 ;
    wire \c0.n45_adj_3138 ;
    wire \c0.n19381 ;
    wire \c0.data_in_frame_7_0 ;
    wire \c0.n7_adj_3355 ;
    wire \c0.data_in_frame_17_5 ;
    wire \c0.n11590 ;
    wire \c0.n14_adj_3449 ;
    wire rx_data_0;
    wire \c0.data_in_frame_15_1 ;
    wire \c0.data_in_frame_14_7 ;
    wire \c0.data_in_frame_14_6 ;
    wire \c0.n19554 ;
    wire \c0.data_in_frame_17_4 ;
    wire \c0.n18_adj_3235 ;
    wire \c0.data_in_frame_15_3 ;
    wire \c0.n10_adj_3483 ;
    wire \c0.n18420 ;
    wire \c0.n19251 ;
    wire \c0.n7_adj_3347 ;
    wire \c0.data_in_frame_10_6 ;
    wire \c0.n19359 ;
    wire \c0.data_in_frame_12_6 ;
    wire \c0.n22_adj_3535 ;
    wire \c0.data_in_frame_20_1 ;
    wire \c0.n12_adj_3265 ;
    wire \c0.data_in_frame_12_3 ;
    wire data_in_frame_19_2;
    wire data_in_frame_19_5;
    wire data_in_frame_19_1;
    wire \c0.n6166 ;
    wire n19130;
    wire data_in_frame_16_2;
    wire \c0.data_in_frame_28_5 ;
    wire \c0.n19111 ;
    wire \c0.data_in_frame_29_3 ;
    wire \c0.n12_adj_3006 ;
    wire \c0.data_in_frame_29_5 ;
    wire \c0.n15_adj_3432 ;
    wire \c0.n20503 ;
    wire data_in_frame_23_1;
    wire \c0.n20503_cascade_ ;
    wire \c0.n12_adj_3494 ;
    wire \c0.n27_adj_3399 ;
    wire \c0.data_in_frame_28_3 ;
    wire \c0.n27_adj_3399_cascade_ ;
    wire \c0.data_in_frame_26_1 ;
    wire \c0.n78_adj_3414 ;
    wire data_in_frame_23_6;
    wire data_in_frame_23_5;
    wire \c0.n19487 ;
    wire data_in_frame_23_7;
    wire \c0.n11971 ;
    wire \c0.n19484 ;
    wire \c0.n7_adj_3072_cascade_ ;
    wire \c0.n18413_cascade_ ;
    wire \c0.data_in_frame_26_3 ;
    wire n19127;
    wire data_in_frame_22_5;
    wire \c0.n9_adj_3069 ;
    wire \c0.n20451 ;
    wire \c0.n8_adj_3070 ;
    wire \c0.n19315 ;
    wire \c0.n26_adj_3550 ;
    wire \c0.n27_adj_3551 ;
    wire \c0.n25_adj_3553 ;
    wire \c0.n49_adj_3358 ;
    wire \c0.n17832 ;
    wire \c0.n40_adj_3271 ;
    wire rx_data_6;
    wire rx_data_2;
    wire \c0.n19474 ;
    wire \c0.data_in_frame_17_2 ;
    wire \c0.data_in_frame_17_3 ;
    wire \c0.n14_adj_3436 ;
    wire \c0.data_in_frame_20_4 ;
    wire \c0.n19274 ;
    wire \c0.data_in_frame_20_3 ;
    wire \c0.n54_adj_3388 ;
    wire \c0.n32_adj_3310 ;
    wire \c0.n43_adj_3131 ;
    wire rx_data_5;
    wire \c0.data_in_frame_20_2 ;
    wire \c0.n20840 ;
    wire \c0.n22_adj_3322 ;
    wire \c0.n22_adj_3322_cascade_ ;
    wire \c0.n36_adj_3090 ;
    wire \c0.data_in_frame_21_2 ;
    wire \c0.n29_adj_3383 ;
    wire \c0.n20917 ;
    wire \c0.data_in_frame_20_0 ;
    wire \c0.n4_adj_3435 ;
    wire \c0.n6_adj_3091 ;
    wire \c0.n18375 ;
    wire \c0.n6_adj_3091_cascade_ ;
    wire \c0.n17900 ;
    wire \c0.data_in_frame_21_3 ;
    wire \c0.data_in_frame_21_5 ;
    wire \c0.n19321 ;
    wire \c0.n12037 ;
    wire data_in_frame_19_7;
    wire rx_data_3;
    wire n19128;
    wire data_in_frame_19_3;
    wire \c0.n19162 ;
    wire data_in_frame_22_1;
    wire \c0.n20332 ;
    wire data_in_frame_24_1;
    wire data_in_frame_24_3;
    wire \c0.n20332_cascade_ ;
    wire \c0.n18413 ;
    wire \c0.n36 ;
    wire \c0.n20642 ;
    wire \c0.n18525 ;
    wire data_in_frame_24_2;
    wire \c0.n18498 ;
    wire \c0.n10_adj_3410 ;
    wire \c0.data_in_frame_20_7 ;
    wire \c0.data_in_frame_20_6 ;
    wire \c0.n20576 ;
    wire \c0.n12_adj_3439 ;
    wire data_in_frame_22_0;
    wire \c0.n18415 ;
    wire \c0.n4_adj_3067_cascade_ ;
    wire \c0.n6009 ;
    wire \c0.n19369 ;
    wire data_in_frame_19_4;
    wire \c0.n11669 ;
    wire rx_data_4;
    wire \c0.data_in_frame_21_6 ;
    wire \c0.data_in_frame_20_5 ;
    wire \c0.data_in_frame_21_4 ;
    wire \c0.n11939_cascade_ ;
    wire data_in_frame_19_6;
    wire \c0.n13_adj_3485 ;
    wire rx_data_7;
    wire \c0.data_in_frame_21_7 ;
    wire \c0.n19107 ;
    wire \c0.n12_adj_3361 ;
    wire rx_data_1;
    wire \c0.data_in_frame_21_1 ;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__73031),
            .DIN(N__73030),
            .DOUT(N__73029),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__73031),
            .PADOUT(N__73030),
            .PADIN(N__73029),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24736),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_12_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_12_pad_iopad (
            .OE(N__73022),
            .DIN(N__73021),
            .DOUT(N__73020),
            .PACKAGEPIN(PIN_12));
    defparam PIN_12_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_12_pad_preio (
            .PADOEN(N__73022),
            .PADOUT(N__73021),
            .PADIN(N__73020),
            .CLOCKENABLE(),
            .DIN0(PIN_12_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_13_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_13_pad_iopad (
            .OE(N__73013),
            .DIN(N__73012),
            .DOUT(N__73011),
            .PACKAGEPIN(PIN_13));
    defparam PIN_13_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_13_pad_preio (
            .PADOEN(N__73013),
            .PADOUT(N__73012),
            .PADIN(N__73011),
            .CLOCKENABLE(),
            .DIN0(PIN_13_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_1_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_1_pad_iopad (
            .OE(N__73004),
            .DIN(N__73003),
            .DOUT(N__73002),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_1_pad_preio (
            .PADOEN(N__73004),
            .PADOUT(N__73003),
            .PADIN(N__73002),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_22_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_22_pad_iopad (
            .OE(N__72995),
            .DIN(N__72994),
            .DOUT(N__72993),
            .PACKAGEPIN(PIN_22));
    defparam PIN_22_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_22_pad_preio (
            .PADOEN(N__72995),
            .PADOUT(N__72994),
            .PADIN(N__72993),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_23_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_23_pad_iopad (
            .OE(N__72986),
            .DIN(N__72985),
            .DOUT(N__72984),
            .PACKAGEPIN(PIN_23));
    defparam PIN_23_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_23_pad_preio (
            .PADOEN(N__72986),
            .PADOUT(N__72985),
            .PADIN(N__72984),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_24_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_24_pad_iopad (
            .OE(N__72977),
            .DIN(N__72976),
            .DOUT(N__72975),
            .PACKAGEPIN(PIN_24));
    defparam PIN_24_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_24_pad_preio (
            .PADOEN(N__72977),
            .PADOUT(N__72976),
            .PADIN(N__72975),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__72968),
            .DIN(N__72967),
            .DOUT(N__72966),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__72968),
            .PADOUT(N__72967),
            .PADIN(N__72966),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_3_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_3_pad_iopad (
            .OE(N__72959),
            .DIN(N__72958),
            .DOUT(N__72957),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_3_pad_preio (
            .PADOEN(N__72959),
            .PADOUT(N__72958),
            .PADIN(N__72957),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_7_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_7_pad_iopad (
            .OE(N__72950),
            .DIN(N__72949),
            .DOUT(N__72948),
            .PACKAGEPIN(PIN_7));
    defparam PIN_7_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_7_pad_preio (
            .PADOEN(N__72950),
            .PADOUT(N__72949),
            .PADIN(N__72948),
            .CLOCKENABLE(),
            .DIN0(PIN_7_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_8_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_8_pad_iopad (
            .OE(N__72941),
            .DIN(N__72940),
            .DOUT(N__72939),
            .PACKAGEPIN(PIN_8));
    defparam PIN_8_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_8_pad_preio (
            .PADOEN(N__72941),
            .PADOUT(N__72940),
            .PADIN(N__72939),
            .CLOCKENABLE(),
            .DIN0(PIN_8_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__72932),
            .DIN(N__72931),
            .DOUT(N__72930),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__72932),
            .PADOUT(N__72931),
            .PADIN(N__72930),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__72923),
            .DIN(N__72922),
            .DOUT(N__72921),
            .PACKAGEPIN(PIN_4));
    defparam hall1_input_preio.PIN_TYPE=6'b000001;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__72923),
            .PADOUT(N__72922),
            .PADIN(N__72921),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__72914),
            .DIN(N__72913),
            .DOUT(N__72912),
            .PACKAGEPIN(PIN_5));
    defparam hall2_input_preio.PIN_TYPE=6'b000001;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__72914),
            .PADOUT(N__72913),
            .PADIN(N__72912),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__72905),
            .DIN(N__72904),
            .DOUT(N__72903),
            .PACKAGEPIN(PIN_6));
    defparam hall3_input_preio.PIN_TYPE=6'b000001;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__72905),
            .PADOUT(N__72904),
            .PADIN(N__72903),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__72896),
            .DIN(N__72895),
            .DOUT(N__72894),
            .PACKAGEPIN(PIN_11));
    defparam rx_input_preio.PIN_TYPE=6'b000001;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__72896),
            .PADOUT(N__72895),
            .PADIN(N__72894),
            .CLOCKENABLE(),
            .DIN0(LED_c),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__72887),
            .DIN(N__72886),
            .DOUT(N__72885),
            .PACKAGEPIN(PIN_10));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__72887),
            .PADOUT(N__72886),
            .PADIN(N__72885),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34183),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__24745));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__72878),
            .DIN(N__72877),
            .DOUT(N__72876),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__72878),
            .PADOUT(N__72877),
            .PADIN(N__72876),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__18132 (
            .O(N__72859),
            .I(N__72855));
    InMux I__18131 (
            .O(N__72858),
            .I(N__72852));
    LocalMux I__18130 (
            .O(N__72855),
            .I(N__72848));
    LocalMux I__18129 (
            .O(N__72852),
            .I(N__72845));
    CascadeMux I__18128 (
            .O(N__72851),
            .I(N__72841));
    Span4Mux_h I__18127 (
            .O(N__72848),
            .I(N__72838));
    Span4Mux_v I__18126 (
            .O(N__72845),
            .I(N__72835));
    CascadeMux I__18125 (
            .O(N__72844),
            .I(N__72828));
    InMux I__18124 (
            .O(N__72841),
            .I(N__72824));
    Span4Mux_v I__18123 (
            .O(N__72838),
            .I(N__72819));
    Span4Mux_h I__18122 (
            .O(N__72835),
            .I(N__72819));
    InMux I__18121 (
            .O(N__72834),
            .I(N__72812));
    InMux I__18120 (
            .O(N__72833),
            .I(N__72812));
    InMux I__18119 (
            .O(N__72832),
            .I(N__72812));
    InMux I__18118 (
            .O(N__72831),
            .I(N__72809));
    InMux I__18117 (
            .O(N__72828),
            .I(N__72806));
    InMux I__18116 (
            .O(N__72827),
            .I(N__72803));
    LocalMux I__18115 (
            .O(N__72824),
            .I(N__72800));
    Sp12to4 I__18114 (
            .O(N__72819),
            .I(N__72795));
    LocalMux I__18113 (
            .O(N__72812),
            .I(N__72795));
    LocalMux I__18112 (
            .O(N__72809),
            .I(N__72790));
    LocalMux I__18111 (
            .O(N__72806),
            .I(N__72790));
    LocalMux I__18110 (
            .O(N__72803),
            .I(data_in_frame_19_4));
    Odrv4 I__18109 (
            .O(N__72800),
            .I(data_in_frame_19_4));
    Odrv12 I__18108 (
            .O(N__72795),
            .I(data_in_frame_19_4));
    Odrv4 I__18107 (
            .O(N__72790),
            .I(data_in_frame_19_4));
    InMux I__18106 (
            .O(N__72781),
            .I(N__72778));
    LocalMux I__18105 (
            .O(N__72778),
            .I(\c0.n11669 ));
    InMux I__18104 (
            .O(N__72775),
            .I(N__72771));
    InMux I__18103 (
            .O(N__72774),
            .I(N__72768));
    LocalMux I__18102 (
            .O(N__72771),
            .I(N__72761));
    LocalMux I__18101 (
            .O(N__72768),
            .I(N__72761));
    InMux I__18100 (
            .O(N__72767),
            .I(N__72756));
    InMux I__18099 (
            .O(N__72766),
            .I(N__72756));
    Span4Mux_h I__18098 (
            .O(N__72761),
            .I(N__72749));
    LocalMux I__18097 (
            .O(N__72756),
            .I(N__72749));
    CascadeMux I__18096 (
            .O(N__72755),
            .I(N__72745));
    InMux I__18095 (
            .O(N__72754),
            .I(N__72741));
    Span4Mux_v I__18094 (
            .O(N__72749),
            .I(N__72734));
    InMux I__18093 (
            .O(N__72748),
            .I(N__72730));
    InMux I__18092 (
            .O(N__72745),
            .I(N__72726));
    InMux I__18091 (
            .O(N__72744),
            .I(N__72723));
    LocalMux I__18090 (
            .O(N__72741),
            .I(N__72720));
    InMux I__18089 (
            .O(N__72740),
            .I(N__72717));
    InMux I__18088 (
            .O(N__72739),
            .I(N__72712));
    InMux I__18087 (
            .O(N__72738),
            .I(N__72712));
    InMux I__18086 (
            .O(N__72737),
            .I(N__72707));
    Span4Mux_h I__18085 (
            .O(N__72734),
            .I(N__72704));
    InMux I__18084 (
            .O(N__72733),
            .I(N__72701));
    LocalMux I__18083 (
            .O(N__72730),
            .I(N__72694));
    InMux I__18082 (
            .O(N__72729),
            .I(N__72691));
    LocalMux I__18081 (
            .O(N__72726),
            .I(N__72686));
    LocalMux I__18080 (
            .O(N__72723),
            .I(N__72686));
    Span4Mux_v I__18079 (
            .O(N__72720),
            .I(N__72681));
    LocalMux I__18078 (
            .O(N__72717),
            .I(N__72681));
    LocalMux I__18077 (
            .O(N__72712),
            .I(N__72678));
    InMux I__18076 (
            .O(N__72711),
            .I(N__72674));
    InMux I__18075 (
            .O(N__72710),
            .I(N__72669));
    LocalMux I__18074 (
            .O(N__72707),
            .I(N__72666));
    Span4Mux_h I__18073 (
            .O(N__72704),
            .I(N__72661));
    LocalMux I__18072 (
            .O(N__72701),
            .I(N__72661));
    InMux I__18071 (
            .O(N__72700),
            .I(N__72656));
    InMux I__18070 (
            .O(N__72699),
            .I(N__72653));
    InMux I__18069 (
            .O(N__72698),
            .I(N__72650));
    InMux I__18068 (
            .O(N__72697),
            .I(N__72646));
    Span4Mux_v I__18067 (
            .O(N__72694),
            .I(N__72641));
    LocalMux I__18066 (
            .O(N__72691),
            .I(N__72641));
    Span4Mux_v I__18065 (
            .O(N__72686),
            .I(N__72636));
    Span4Mux_h I__18064 (
            .O(N__72681),
            .I(N__72636));
    Span4Mux_h I__18063 (
            .O(N__72678),
            .I(N__72633));
    InMux I__18062 (
            .O(N__72677),
            .I(N__72630));
    LocalMux I__18061 (
            .O(N__72674),
            .I(N__72627));
    InMux I__18060 (
            .O(N__72673),
            .I(N__72622));
    InMux I__18059 (
            .O(N__72672),
            .I(N__72622));
    LocalMux I__18058 (
            .O(N__72669),
            .I(N__72615));
    Span4Mux_v I__18057 (
            .O(N__72666),
            .I(N__72615));
    Span4Mux_v I__18056 (
            .O(N__72661),
            .I(N__72615));
    InMux I__18055 (
            .O(N__72660),
            .I(N__72607));
    InMux I__18054 (
            .O(N__72659),
            .I(N__72604));
    LocalMux I__18053 (
            .O(N__72656),
            .I(N__72601));
    LocalMux I__18052 (
            .O(N__72653),
            .I(N__72598));
    LocalMux I__18051 (
            .O(N__72650),
            .I(N__72595));
    InMux I__18050 (
            .O(N__72649),
            .I(N__72592));
    LocalMux I__18049 (
            .O(N__72646),
            .I(N__72589));
    Span4Mux_v I__18048 (
            .O(N__72641),
            .I(N__72584));
    Span4Mux_h I__18047 (
            .O(N__72636),
            .I(N__72584));
    Span4Mux_h I__18046 (
            .O(N__72633),
            .I(N__72575));
    LocalMux I__18045 (
            .O(N__72630),
            .I(N__72575));
    Span4Mux_h I__18044 (
            .O(N__72627),
            .I(N__72575));
    LocalMux I__18043 (
            .O(N__72622),
            .I(N__72575));
    Sp12to4 I__18042 (
            .O(N__72615),
            .I(N__72572));
    InMux I__18041 (
            .O(N__72614),
            .I(N__72569));
    InMux I__18040 (
            .O(N__72613),
            .I(N__72566));
    InMux I__18039 (
            .O(N__72612),
            .I(N__72563));
    InMux I__18038 (
            .O(N__72611),
            .I(N__72558));
    InMux I__18037 (
            .O(N__72610),
            .I(N__72558));
    LocalMux I__18036 (
            .O(N__72607),
            .I(N__72549));
    LocalMux I__18035 (
            .O(N__72604),
            .I(N__72549));
    Span4Mux_v I__18034 (
            .O(N__72601),
            .I(N__72549));
    Span4Mux_v I__18033 (
            .O(N__72598),
            .I(N__72549));
    Span4Mux_h I__18032 (
            .O(N__72595),
            .I(N__72546));
    LocalMux I__18031 (
            .O(N__72592),
            .I(N__72541));
    Span4Mux_v I__18030 (
            .O(N__72589),
            .I(N__72541));
    Span4Mux_v I__18029 (
            .O(N__72584),
            .I(N__72538));
    Span4Mux_v I__18028 (
            .O(N__72575),
            .I(N__72535));
    Span12Mux_h I__18027 (
            .O(N__72572),
            .I(N__72532));
    LocalMux I__18026 (
            .O(N__72569),
            .I(N__72528));
    LocalMux I__18025 (
            .O(N__72566),
            .I(N__72525));
    LocalMux I__18024 (
            .O(N__72563),
            .I(N__72522));
    LocalMux I__18023 (
            .O(N__72558),
            .I(N__72517));
    Span4Mux_h I__18022 (
            .O(N__72549),
            .I(N__72517));
    Span4Mux_h I__18021 (
            .O(N__72546),
            .I(N__72510));
    Span4Mux_h I__18020 (
            .O(N__72541),
            .I(N__72510));
    Span4Mux_v I__18019 (
            .O(N__72538),
            .I(N__72510));
    Sp12to4 I__18018 (
            .O(N__72535),
            .I(N__72505));
    Span12Mux_v I__18017 (
            .O(N__72532),
            .I(N__72505));
    InMux I__18016 (
            .O(N__72531),
            .I(N__72502));
    Span4Mux_h I__18015 (
            .O(N__72528),
            .I(N__72499));
    Span4Mux_v I__18014 (
            .O(N__72525),
            .I(N__72496));
    Span4Mux_h I__18013 (
            .O(N__72522),
            .I(N__72491));
    Span4Mux_v I__18012 (
            .O(N__72517),
            .I(N__72491));
    Sp12to4 I__18011 (
            .O(N__72510),
            .I(N__72486));
    Span12Mux_h I__18010 (
            .O(N__72505),
            .I(N__72486));
    LocalMux I__18009 (
            .O(N__72502),
            .I(rx_data_4));
    Odrv4 I__18008 (
            .O(N__72499),
            .I(rx_data_4));
    Odrv4 I__18007 (
            .O(N__72496),
            .I(rx_data_4));
    Odrv4 I__18006 (
            .O(N__72491),
            .I(rx_data_4));
    Odrv12 I__18005 (
            .O(N__72486),
            .I(rx_data_4));
    InMux I__18004 (
            .O(N__72475),
            .I(N__72468));
    InMux I__18003 (
            .O(N__72474),
            .I(N__72468));
    CascadeMux I__18002 (
            .O(N__72473),
            .I(N__72463));
    LocalMux I__18001 (
            .O(N__72468),
            .I(N__72460));
    InMux I__18000 (
            .O(N__72467),
            .I(N__72455));
    InMux I__17999 (
            .O(N__72466),
            .I(N__72455));
    InMux I__17998 (
            .O(N__72463),
            .I(N__72452));
    Span4Mux_v I__17997 (
            .O(N__72460),
            .I(N__72449));
    LocalMux I__17996 (
            .O(N__72455),
            .I(N__72446));
    LocalMux I__17995 (
            .O(N__72452),
            .I(\c0.data_in_frame_21_6 ));
    Odrv4 I__17994 (
            .O(N__72449),
            .I(\c0.data_in_frame_21_6 ));
    Odrv4 I__17993 (
            .O(N__72446),
            .I(\c0.data_in_frame_21_6 ));
    InMux I__17992 (
            .O(N__72439),
            .I(N__72434));
    InMux I__17991 (
            .O(N__72438),
            .I(N__72429));
    InMux I__17990 (
            .O(N__72437),
            .I(N__72429));
    LocalMux I__17989 (
            .O(N__72434),
            .I(N__72426));
    LocalMux I__17988 (
            .O(N__72429),
            .I(N__72421));
    Span4Mux_v I__17987 (
            .O(N__72426),
            .I(N__72418));
    InMux I__17986 (
            .O(N__72425),
            .I(N__72415));
    InMux I__17985 (
            .O(N__72424),
            .I(N__72412));
    Span12Mux_s11_v I__17984 (
            .O(N__72421),
            .I(N__72409));
    Span4Mux_v I__17983 (
            .O(N__72418),
            .I(N__72404));
    LocalMux I__17982 (
            .O(N__72415),
            .I(N__72404));
    LocalMux I__17981 (
            .O(N__72412),
            .I(\c0.data_in_frame_20_5 ));
    Odrv12 I__17980 (
            .O(N__72409),
            .I(\c0.data_in_frame_20_5 ));
    Odrv4 I__17979 (
            .O(N__72404),
            .I(\c0.data_in_frame_20_5 ));
    CascadeMux I__17978 (
            .O(N__72397),
            .I(N__72394));
    InMux I__17977 (
            .O(N__72394),
            .I(N__72389));
    CascadeMux I__17976 (
            .O(N__72393),
            .I(N__72386));
    InMux I__17975 (
            .O(N__72392),
            .I(N__72382));
    LocalMux I__17974 (
            .O(N__72389),
            .I(N__72379));
    InMux I__17973 (
            .O(N__72386),
            .I(N__72376));
    InMux I__17972 (
            .O(N__72385),
            .I(N__72373));
    LocalMux I__17971 (
            .O(N__72382),
            .I(N__72370));
    Span4Mux_v I__17970 (
            .O(N__72379),
            .I(N__72366));
    LocalMux I__17969 (
            .O(N__72376),
            .I(N__72359));
    LocalMux I__17968 (
            .O(N__72373),
            .I(N__72359));
    Span4Mux_v I__17967 (
            .O(N__72370),
            .I(N__72359));
    InMux I__17966 (
            .O(N__72369),
            .I(N__72356));
    Odrv4 I__17965 (
            .O(N__72366),
            .I(\c0.data_in_frame_21_4 ));
    Odrv4 I__17964 (
            .O(N__72359),
            .I(\c0.data_in_frame_21_4 ));
    LocalMux I__17963 (
            .O(N__72356),
            .I(\c0.data_in_frame_21_4 ));
    CascadeMux I__17962 (
            .O(N__72349),
            .I(\c0.n11939_cascade_ ));
    InMux I__17961 (
            .O(N__72346),
            .I(N__72343));
    LocalMux I__17960 (
            .O(N__72343),
            .I(N__72339));
    CascadeMux I__17959 (
            .O(N__72342),
            .I(N__72332));
    Span4Mux_v I__17958 (
            .O(N__72339),
            .I(N__72329));
    InMux I__17957 (
            .O(N__72338),
            .I(N__72324));
    InMux I__17956 (
            .O(N__72337),
            .I(N__72324));
    InMux I__17955 (
            .O(N__72336),
            .I(N__72319));
    InMux I__17954 (
            .O(N__72335),
            .I(N__72319));
    InMux I__17953 (
            .O(N__72332),
            .I(N__72316));
    Sp12to4 I__17952 (
            .O(N__72329),
            .I(N__72309));
    LocalMux I__17951 (
            .O(N__72324),
            .I(N__72309));
    LocalMux I__17950 (
            .O(N__72319),
            .I(N__72309));
    LocalMux I__17949 (
            .O(N__72316),
            .I(data_in_frame_19_6));
    Odrv12 I__17948 (
            .O(N__72309),
            .I(data_in_frame_19_6));
    InMux I__17947 (
            .O(N__72304),
            .I(N__72301));
    LocalMux I__17946 (
            .O(N__72301),
            .I(N__72298));
    Odrv4 I__17945 (
            .O(N__72298),
            .I(\c0.n13_adj_3485 ));
    InMux I__17944 (
            .O(N__72295),
            .I(N__72288));
    InMux I__17943 (
            .O(N__72294),
            .I(N__72280));
    InMux I__17942 (
            .O(N__72293),
            .I(N__72277));
    InMux I__17941 (
            .O(N__72292),
            .I(N__72274));
    InMux I__17940 (
            .O(N__72291),
            .I(N__72271));
    LocalMux I__17939 (
            .O(N__72288),
            .I(N__72267));
    InMux I__17938 (
            .O(N__72287),
            .I(N__72262));
    InMux I__17937 (
            .O(N__72286),
            .I(N__72262));
    InMux I__17936 (
            .O(N__72285),
            .I(N__72257));
    InMux I__17935 (
            .O(N__72284),
            .I(N__72251));
    InMux I__17934 (
            .O(N__72283),
            .I(N__72248));
    LocalMux I__17933 (
            .O(N__72280),
            .I(N__72243));
    LocalMux I__17932 (
            .O(N__72277),
            .I(N__72243));
    LocalMux I__17931 (
            .O(N__72274),
            .I(N__72238));
    LocalMux I__17930 (
            .O(N__72271),
            .I(N__72235));
    CascadeMux I__17929 (
            .O(N__72270),
            .I(N__72232));
    Span4Mux_h I__17928 (
            .O(N__72267),
            .I(N__72228));
    LocalMux I__17927 (
            .O(N__72262),
            .I(N__72225));
    InMux I__17926 (
            .O(N__72261),
            .I(N__72222));
    InMux I__17925 (
            .O(N__72260),
            .I(N__72218));
    LocalMux I__17924 (
            .O(N__72257),
            .I(N__72214));
    InMux I__17923 (
            .O(N__72256),
            .I(N__72211));
    InMux I__17922 (
            .O(N__72255),
            .I(N__72208));
    InMux I__17921 (
            .O(N__72254),
            .I(N__72202));
    LocalMux I__17920 (
            .O(N__72251),
            .I(N__72196));
    LocalMux I__17919 (
            .O(N__72248),
            .I(N__72193));
    Span4Mux_h I__17918 (
            .O(N__72243),
            .I(N__72190));
    InMux I__17917 (
            .O(N__72242),
            .I(N__72187));
    InMux I__17916 (
            .O(N__72241),
            .I(N__72184));
    Span4Mux_v I__17915 (
            .O(N__72238),
            .I(N__72181));
    Span4Mux_v I__17914 (
            .O(N__72235),
            .I(N__72178));
    InMux I__17913 (
            .O(N__72232),
            .I(N__72175));
    InMux I__17912 (
            .O(N__72231),
            .I(N__72172));
    Span4Mux_v I__17911 (
            .O(N__72228),
            .I(N__72165));
    Span4Mux_v I__17910 (
            .O(N__72225),
            .I(N__72165));
    LocalMux I__17909 (
            .O(N__72222),
            .I(N__72165));
    InMux I__17908 (
            .O(N__72221),
            .I(N__72162));
    LocalMux I__17907 (
            .O(N__72218),
            .I(N__72159));
    InMux I__17906 (
            .O(N__72217),
            .I(N__72156));
    Span4Mux_v I__17905 (
            .O(N__72214),
            .I(N__72153));
    LocalMux I__17904 (
            .O(N__72211),
            .I(N__72150));
    LocalMux I__17903 (
            .O(N__72208),
            .I(N__72146));
    InMux I__17902 (
            .O(N__72207),
            .I(N__72141));
    InMux I__17901 (
            .O(N__72206),
            .I(N__72136));
    InMux I__17900 (
            .O(N__72205),
            .I(N__72136));
    LocalMux I__17899 (
            .O(N__72202),
            .I(N__72133));
    CascadeMux I__17898 (
            .O(N__72201),
            .I(N__72129));
    InMux I__17897 (
            .O(N__72200),
            .I(N__72125));
    InMux I__17896 (
            .O(N__72199),
            .I(N__72122));
    Span4Mux_v I__17895 (
            .O(N__72196),
            .I(N__72117));
    Span4Mux_v I__17894 (
            .O(N__72193),
            .I(N__72117));
    Span4Mux_h I__17893 (
            .O(N__72190),
            .I(N__72114));
    LocalMux I__17892 (
            .O(N__72187),
            .I(N__72105));
    LocalMux I__17891 (
            .O(N__72184),
            .I(N__72105));
    Sp12to4 I__17890 (
            .O(N__72181),
            .I(N__72105));
    Sp12to4 I__17889 (
            .O(N__72178),
            .I(N__72105));
    LocalMux I__17888 (
            .O(N__72175),
            .I(N__72100));
    LocalMux I__17887 (
            .O(N__72172),
            .I(N__72100));
    Span4Mux_h I__17886 (
            .O(N__72165),
            .I(N__72097));
    LocalMux I__17885 (
            .O(N__72162),
            .I(N__72092));
    Span4Mux_h I__17884 (
            .O(N__72159),
            .I(N__72092));
    LocalMux I__17883 (
            .O(N__72156),
            .I(N__72085));
    Span4Mux_h I__17882 (
            .O(N__72153),
            .I(N__72085));
    Span4Mux_h I__17881 (
            .O(N__72150),
            .I(N__72085));
    InMux I__17880 (
            .O(N__72149),
            .I(N__72082));
    Span4Mux_h I__17879 (
            .O(N__72146),
            .I(N__72079));
    InMux I__17878 (
            .O(N__72145),
            .I(N__72074));
    InMux I__17877 (
            .O(N__72144),
            .I(N__72074));
    LocalMux I__17876 (
            .O(N__72141),
            .I(N__72071));
    LocalMux I__17875 (
            .O(N__72136),
            .I(N__72066));
    Span4Mux_v I__17874 (
            .O(N__72133),
            .I(N__72066));
    InMux I__17873 (
            .O(N__72132),
            .I(N__72059));
    InMux I__17872 (
            .O(N__72129),
            .I(N__72059));
    InMux I__17871 (
            .O(N__72128),
            .I(N__72059));
    LocalMux I__17870 (
            .O(N__72125),
            .I(N__72054));
    LocalMux I__17869 (
            .O(N__72122),
            .I(N__72054));
    Span4Mux_v I__17868 (
            .O(N__72117),
            .I(N__72051));
    Sp12to4 I__17867 (
            .O(N__72114),
            .I(N__72046));
    Span12Mux_h I__17866 (
            .O(N__72105),
            .I(N__72046));
    Span4Mux_v I__17865 (
            .O(N__72100),
            .I(N__72043));
    Span4Mux_h I__17864 (
            .O(N__72097),
            .I(N__72036));
    Span4Mux_h I__17863 (
            .O(N__72092),
            .I(N__72036));
    Span4Mux_v I__17862 (
            .O(N__72085),
            .I(N__72036));
    LocalMux I__17861 (
            .O(N__72082),
            .I(N__72031));
    Sp12to4 I__17860 (
            .O(N__72079),
            .I(N__72031));
    LocalMux I__17859 (
            .O(N__72074),
            .I(N__72024));
    Span4Mux_h I__17858 (
            .O(N__72071),
            .I(N__72024));
    Span4Mux_v I__17857 (
            .O(N__72066),
            .I(N__72024));
    LocalMux I__17856 (
            .O(N__72059),
            .I(N__72019));
    Span12Mux_s11_v I__17855 (
            .O(N__72054),
            .I(N__72019));
    Sp12to4 I__17854 (
            .O(N__72051),
            .I(N__72014));
    Span12Mux_v I__17853 (
            .O(N__72046),
            .I(N__72014));
    Span4Mux_h I__17852 (
            .O(N__72043),
            .I(N__72009));
    Span4Mux_v I__17851 (
            .O(N__72036),
            .I(N__72009));
    Odrv12 I__17850 (
            .O(N__72031),
            .I(rx_data_7));
    Odrv4 I__17849 (
            .O(N__72024),
            .I(rx_data_7));
    Odrv12 I__17848 (
            .O(N__72019),
            .I(rx_data_7));
    Odrv12 I__17847 (
            .O(N__72014),
            .I(rx_data_7));
    Odrv4 I__17846 (
            .O(N__72009),
            .I(rx_data_7));
    InMux I__17845 (
            .O(N__71998),
            .I(N__71995));
    LocalMux I__17844 (
            .O(N__71995),
            .I(N__71989));
    InMux I__17843 (
            .O(N__71994),
            .I(N__71982));
    InMux I__17842 (
            .O(N__71993),
            .I(N__71982));
    InMux I__17841 (
            .O(N__71992),
            .I(N__71982));
    Odrv4 I__17840 (
            .O(N__71989),
            .I(\c0.data_in_frame_21_7 ));
    LocalMux I__17839 (
            .O(N__71982),
            .I(\c0.data_in_frame_21_7 ));
    InMux I__17838 (
            .O(N__71977),
            .I(N__71974));
    LocalMux I__17837 (
            .O(N__71974),
            .I(N__71966));
    CascadeMux I__17836 (
            .O(N__71973),
            .I(N__71955));
    InMux I__17835 (
            .O(N__71972),
            .I(N__71952));
    InMux I__17834 (
            .O(N__71971),
            .I(N__71949));
    InMux I__17833 (
            .O(N__71970),
            .I(N__71942));
    InMux I__17832 (
            .O(N__71969),
            .I(N__71942));
    Span4Mux_h I__17831 (
            .O(N__71966),
            .I(N__71938));
    InMux I__17830 (
            .O(N__71965),
            .I(N__71935));
    InMux I__17829 (
            .O(N__71964),
            .I(N__71929));
    InMux I__17828 (
            .O(N__71963),
            .I(N__71922));
    InMux I__17827 (
            .O(N__71962),
            .I(N__71922));
    InMux I__17826 (
            .O(N__71961),
            .I(N__71922));
    InMux I__17825 (
            .O(N__71960),
            .I(N__71917));
    InMux I__17824 (
            .O(N__71959),
            .I(N__71917));
    InMux I__17823 (
            .O(N__71958),
            .I(N__71912));
    InMux I__17822 (
            .O(N__71955),
            .I(N__71912));
    LocalMux I__17821 (
            .O(N__71952),
            .I(N__71907));
    LocalMux I__17820 (
            .O(N__71949),
            .I(N__71907));
    InMux I__17819 (
            .O(N__71948),
            .I(N__71902));
    InMux I__17818 (
            .O(N__71947),
            .I(N__71902));
    LocalMux I__17817 (
            .O(N__71942),
            .I(N__71899));
    InMux I__17816 (
            .O(N__71941),
            .I(N__71895));
    Span4Mux_v I__17815 (
            .O(N__71938),
            .I(N__71890));
    LocalMux I__17814 (
            .O(N__71935),
            .I(N__71890));
    InMux I__17813 (
            .O(N__71934),
            .I(N__71883));
    InMux I__17812 (
            .O(N__71933),
            .I(N__71883));
    InMux I__17811 (
            .O(N__71932),
            .I(N__71883));
    LocalMux I__17810 (
            .O(N__71929),
            .I(N__71876));
    LocalMux I__17809 (
            .O(N__71922),
            .I(N__71876));
    LocalMux I__17808 (
            .O(N__71917),
            .I(N__71876));
    LocalMux I__17807 (
            .O(N__71912),
            .I(N__71871));
    Span4Mux_v I__17806 (
            .O(N__71907),
            .I(N__71871));
    LocalMux I__17805 (
            .O(N__71902),
            .I(N__71863));
    Span4Mux_v I__17804 (
            .O(N__71899),
            .I(N__71863));
    CascadeMux I__17803 (
            .O(N__71898),
            .I(N__71860));
    LocalMux I__17802 (
            .O(N__71895),
            .I(N__71857));
    Span4Mux_h I__17801 (
            .O(N__71890),
            .I(N__71854));
    LocalMux I__17800 (
            .O(N__71883),
            .I(N__71851));
    Span4Mux_v I__17799 (
            .O(N__71876),
            .I(N__71846));
    Span4Mux_v I__17798 (
            .O(N__71871),
            .I(N__71846));
    InMux I__17797 (
            .O(N__71870),
            .I(N__71839));
    InMux I__17796 (
            .O(N__71869),
            .I(N__71839));
    InMux I__17795 (
            .O(N__71868),
            .I(N__71839));
    Span4Mux_v I__17794 (
            .O(N__71863),
            .I(N__71836));
    InMux I__17793 (
            .O(N__71860),
            .I(N__71833));
    Span4Mux_h I__17792 (
            .O(N__71857),
            .I(N__71830));
    Sp12to4 I__17791 (
            .O(N__71854),
            .I(N__71825));
    Span12Mux_h I__17790 (
            .O(N__71851),
            .I(N__71825));
    Span4Mux_h I__17789 (
            .O(N__71846),
            .I(N__71822));
    LocalMux I__17788 (
            .O(N__71839),
            .I(N__71817));
    Span4Mux_h I__17787 (
            .O(N__71836),
            .I(N__71817));
    LocalMux I__17786 (
            .O(N__71833),
            .I(\c0.n19107 ));
    Odrv4 I__17785 (
            .O(N__71830),
            .I(\c0.n19107 ));
    Odrv12 I__17784 (
            .O(N__71825),
            .I(\c0.n19107 ));
    Odrv4 I__17783 (
            .O(N__71822),
            .I(\c0.n19107 ));
    Odrv4 I__17782 (
            .O(N__71817),
            .I(\c0.n19107 ));
    CascadeMux I__17781 (
            .O(N__71806),
            .I(N__71803));
    InMux I__17780 (
            .O(N__71803),
            .I(N__71797));
    InMux I__17779 (
            .O(N__71802),
            .I(N__71794));
    InMux I__17778 (
            .O(N__71801),
            .I(N__71788));
    InMux I__17777 (
            .O(N__71800),
            .I(N__71783));
    LocalMux I__17776 (
            .O(N__71797),
            .I(N__71770));
    LocalMux I__17775 (
            .O(N__71794),
            .I(N__71770));
    InMux I__17774 (
            .O(N__71793),
            .I(N__71767));
    CascadeMux I__17773 (
            .O(N__71792),
            .I(N__71763));
    InMux I__17772 (
            .O(N__71791),
            .I(N__71759));
    LocalMux I__17771 (
            .O(N__71788),
            .I(N__71756));
    InMux I__17770 (
            .O(N__71787),
            .I(N__71749));
    InMux I__17769 (
            .O(N__71786),
            .I(N__71749));
    LocalMux I__17768 (
            .O(N__71783),
            .I(N__71746));
    CascadeMux I__17767 (
            .O(N__71782),
            .I(N__71741));
    CascadeMux I__17766 (
            .O(N__71781),
            .I(N__71735));
    InMux I__17765 (
            .O(N__71780),
            .I(N__71729));
    InMux I__17764 (
            .O(N__71779),
            .I(N__71729));
    InMux I__17763 (
            .O(N__71778),
            .I(N__71726));
    InMux I__17762 (
            .O(N__71777),
            .I(N__71723));
    InMux I__17761 (
            .O(N__71776),
            .I(N__71718));
    InMux I__17760 (
            .O(N__71775),
            .I(N__71718));
    Span4Mux_v I__17759 (
            .O(N__71770),
            .I(N__71713));
    LocalMux I__17758 (
            .O(N__71767),
            .I(N__71713));
    InMux I__17757 (
            .O(N__71766),
            .I(N__71710));
    InMux I__17756 (
            .O(N__71763),
            .I(N__71707));
    InMux I__17755 (
            .O(N__71762),
            .I(N__71704));
    LocalMux I__17754 (
            .O(N__71759),
            .I(N__71701));
    Span4Mux_v I__17753 (
            .O(N__71756),
            .I(N__71698));
    InMux I__17752 (
            .O(N__71755),
            .I(N__71693));
    InMux I__17751 (
            .O(N__71754),
            .I(N__71693));
    LocalMux I__17750 (
            .O(N__71749),
            .I(N__71688));
    Span4Mux_h I__17749 (
            .O(N__71746),
            .I(N__71688));
    InMux I__17748 (
            .O(N__71745),
            .I(N__71681));
    InMux I__17747 (
            .O(N__71744),
            .I(N__71681));
    InMux I__17746 (
            .O(N__71741),
            .I(N__71681));
    InMux I__17745 (
            .O(N__71740),
            .I(N__71678));
    InMux I__17744 (
            .O(N__71739),
            .I(N__71671));
    InMux I__17743 (
            .O(N__71738),
            .I(N__71671));
    InMux I__17742 (
            .O(N__71735),
            .I(N__71671));
    InMux I__17741 (
            .O(N__71734),
            .I(N__71668));
    LocalMux I__17740 (
            .O(N__71729),
            .I(N__71665));
    LocalMux I__17739 (
            .O(N__71726),
            .I(N__71662));
    LocalMux I__17738 (
            .O(N__71723),
            .I(N__71659));
    LocalMux I__17737 (
            .O(N__71718),
            .I(N__71656));
    Span4Mux_h I__17736 (
            .O(N__71713),
            .I(N__71653));
    LocalMux I__17735 (
            .O(N__71710),
            .I(N__71650));
    LocalMux I__17734 (
            .O(N__71707),
            .I(N__71647));
    LocalMux I__17733 (
            .O(N__71704),
            .I(N__71644));
    Span4Mux_v I__17732 (
            .O(N__71701),
            .I(N__71641));
    Span4Mux_h I__17731 (
            .O(N__71698),
            .I(N__71636));
    LocalMux I__17730 (
            .O(N__71693),
            .I(N__71636));
    Span4Mux_h I__17729 (
            .O(N__71688),
            .I(N__71633));
    LocalMux I__17728 (
            .O(N__71681),
            .I(N__71630));
    LocalMux I__17727 (
            .O(N__71678),
            .I(N__71625));
    LocalMux I__17726 (
            .O(N__71671),
            .I(N__71625));
    LocalMux I__17725 (
            .O(N__71668),
            .I(N__71620));
    Span4Mux_h I__17724 (
            .O(N__71665),
            .I(N__71615));
    Span4Mux_v I__17723 (
            .O(N__71662),
            .I(N__71615));
    Span4Mux_h I__17722 (
            .O(N__71659),
            .I(N__71612));
    Span4Mux_h I__17721 (
            .O(N__71656),
            .I(N__71607));
    Span4Mux_h I__17720 (
            .O(N__71653),
            .I(N__71607));
    Span4Mux_h I__17719 (
            .O(N__71650),
            .I(N__71604));
    Span4Mux_h I__17718 (
            .O(N__71647),
            .I(N__71601));
    Span4Mux_v I__17717 (
            .O(N__71644),
            .I(N__71594));
    Span4Mux_v I__17716 (
            .O(N__71641),
            .I(N__71594));
    Span4Mux_h I__17715 (
            .O(N__71636),
            .I(N__71594));
    Span4Mux_v I__17714 (
            .O(N__71633),
            .I(N__71591));
    Span12Mux_v I__17713 (
            .O(N__71630),
            .I(N__71586));
    Span12Mux_v I__17712 (
            .O(N__71625),
            .I(N__71586));
    InMux I__17711 (
            .O(N__71624),
            .I(N__71583));
    InMux I__17710 (
            .O(N__71623),
            .I(N__71580));
    Span4Mux_v I__17709 (
            .O(N__71620),
            .I(N__71573));
    Span4Mux_h I__17708 (
            .O(N__71615),
            .I(N__71573));
    Span4Mux_v I__17707 (
            .O(N__71612),
            .I(N__71573));
    Span4Mux_h I__17706 (
            .O(N__71607),
            .I(N__71570));
    Span4Mux_h I__17705 (
            .O(N__71604),
            .I(N__71563));
    Span4Mux_v I__17704 (
            .O(N__71601),
            .I(N__71563));
    Span4Mux_h I__17703 (
            .O(N__71594),
            .I(N__71563));
    Odrv4 I__17702 (
            .O(N__71591),
            .I(\c0.n12_adj_3361 ));
    Odrv12 I__17701 (
            .O(N__71586),
            .I(\c0.n12_adj_3361 ));
    LocalMux I__17700 (
            .O(N__71583),
            .I(\c0.n12_adj_3361 ));
    LocalMux I__17699 (
            .O(N__71580),
            .I(\c0.n12_adj_3361 ));
    Odrv4 I__17698 (
            .O(N__71573),
            .I(\c0.n12_adj_3361 ));
    Odrv4 I__17697 (
            .O(N__71570),
            .I(\c0.n12_adj_3361 ));
    Odrv4 I__17696 (
            .O(N__71563),
            .I(\c0.n12_adj_3361 ));
    InMux I__17695 (
            .O(N__71548),
            .I(N__71544));
    InMux I__17694 (
            .O(N__71547),
            .I(N__71540));
    LocalMux I__17693 (
            .O(N__71544),
            .I(N__71537));
    InMux I__17692 (
            .O(N__71543),
            .I(N__71531));
    LocalMux I__17691 (
            .O(N__71540),
            .I(N__71528));
    Span4Mux_v I__17690 (
            .O(N__71537),
            .I(N__71521));
    InMux I__17689 (
            .O(N__71536),
            .I(N__71518));
    InMux I__17688 (
            .O(N__71535),
            .I(N__71513));
    InMux I__17687 (
            .O(N__71534),
            .I(N__71513));
    LocalMux I__17686 (
            .O(N__71531),
            .I(N__71510));
    Span4Mux_v I__17685 (
            .O(N__71528),
            .I(N__71507));
    InMux I__17684 (
            .O(N__71527),
            .I(N__71500));
    InMux I__17683 (
            .O(N__71526),
            .I(N__71497));
    CascadeMux I__17682 (
            .O(N__71525),
            .I(N__71493));
    InMux I__17681 (
            .O(N__71524),
            .I(N__71489));
    Span4Mux_h I__17680 (
            .O(N__71521),
            .I(N__71480));
    LocalMux I__17679 (
            .O(N__71518),
            .I(N__71480));
    LocalMux I__17678 (
            .O(N__71513),
            .I(N__71473));
    Span4Mux_v I__17677 (
            .O(N__71510),
            .I(N__71473));
    Span4Mux_h I__17676 (
            .O(N__71507),
            .I(N__71473));
    InMux I__17675 (
            .O(N__71506),
            .I(N__71470));
    InMux I__17674 (
            .O(N__71505),
            .I(N__71467));
    InMux I__17673 (
            .O(N__71504),
            .I(N__71459));
    InMux I__17672 (
            .O(N__71503),
            .I(N__71459));
    LocalMux I__17671 (
            .O(N__71500),
            .I(N__71456));
    LocalMux I__17670 (
            .O(N__71497),
            .I(N__71453));
    InMux I__17669 (
            .O(N__71496),
            .I(N__71450));
    InMux I__17668 (
            .O(N__71493),
            .I(N__71445));
    InMux I__17667 (
            .O(N__71492),
            .I(N__71445));
    LocalMux I__17666 (
            .O(N__71489),
            .I(N__71442));
    InMux I__17665 (
            .O(N__71488),
            .I(N__71437));
    InMux I__17664 (
            .O(N__71487),
            .I(N__71437));
    InMux I__17663 (
            .O(N__71486),
            .I(N__71433));
    InMux I__17662 (
            .O(N__71485),
            .I(N__71430));
    Span4Mux_v I__17661 (
            .O(N__71480),
            .I(N__71427));
    Span4Mux_h I__17660 (
            .O(N__71473),
            .I(N__71420));
    LocalMux I__17659 (
            .O(N__71470),
            .I(N__71420));
    LocalMux I__17658 (
            .O(N__71467),
            .I(N__71420));
    InMux I__17657 (
            .O(N__71466),
            .I(N__71412));
    InMux I__17656 (
            .O(N__71465),
            .I(N__71412));
    InMux I__17655 (
            .O(N__71464),
            .I(N__71412));
    LocalMux I__17654 (
            .O(N__71459),
            .I(N__71409));
    Span4Mux_v I__17653 (
            .O(N__71456),
            .I(N__71404));
    Span4Mux_v I__17652 (
            .O(N__71453),
            .I(N__71404));
    LocalMux I__17651 (
            .O(N__71450),
            .I(N__71399));
    LocalMux I__17650 (
            .O(N__71445),
            .I(N__71399));
    Span4Mux_v I__17649 (
            .O(N__71442),
            .I(N__71394));
    LocalMux I__17648 (
            .O(N__71437),
            .I(N__71394));
    InMux I__17647 (
            .O(N__71436),
            .I(N__71390));
    LocalMux I__17646 (
            .O(N__71433),
            .I(N__71385));
    LocalMux I__17645 (
            .O(N__71430),
            .I(N__71385));
    Sp12to4 I__17644 (
            .O(N__71427),
            .I(N__71380));
    Sp12to4 I__17643 (
            .O(N__71420),
            .I(N__71380));
    InMux I__17642 (
            .O(N__71419),
            .I(N__71377));
    LocalMux I__17641 (
            .O(N__71412),
            .I(N__71369));
    Span12Mux_v I__17640 (
            .O(N__71409),
            .I(N__71369));
    Span4Mux_h I__17639 (
            .O(N__71404),
            .I(N__71362));
    Span4Mux_h I__17638 (
            .O(N__71399),
            .I(N__71362));
    Span4Mux_v I__17637 (
            .O(N__71394),
            .I(N__71362));
    InMux I__17636 (
            .O(N__71393),
            .I(N__71359));
    LocalMux I__17635 (
            .O(N__71390),
            .I(N__71356));
    Span4Mux_h I__17634 (
            .O(N__71385),
            .I(N__71353));
    Span12Mux_h I__17633 (
            .O(N__71380),
            .I(N__71350));
    LocalMux I__17632 (
            .O(N__71377),
            .I(N__71344));
    InMux I__17631 (
            .O(N__71376),
            .I(N__71341));
    InMux I__17630 (
            .O(N__71375),
            .I(N__71336));
    InMux I__17629 (
            .O(N__71374),
            .I(N__71336));
    Span12Mux_h I__17628 (
            .O(N__71369),
            .I(N__71333));
    Sp12to4 I__17627 (
            .O(N__71362),
            .I(N__71330));
    LocalMux I__17626 (
            .O(N__71359),
            .I(N__71323));
    Span4Mux_h I__17625 (
            .O(N__71356),
            .I(N__71323));
    Span4Mux_v I__17624 (
            .O(N__71353),
            .I(N__71323));
    Span12Mux_v I__17623 (
            .O(N__71350),
            .I(N__71320));
    InMux I__17622 (
            .O(N__71349),
            .I(N__71315));
    InMux I__17621 (
            .O(N__71348),
            .I(N__71315));
    InMux I__17620 (
            .O(N__71347),
            .I(N__71312));
    Span4Mux_h I__17619 (
            .O(N__71344),
            .I(N__71307));
    LocalMux I__17618 (
            .O(N__71341),
            .I(N__71307));
    LocalMux I__17617 (
            .O(N__71336),
            .I(N__71302));
    Span12Mux_v I__17616 (
            .O(N__71333),
            .I(N__71302));
    Span12Mux_h I__17615 (
            .O(N__71330),
            .I(N__71295));
    Sp12to4 I__17614 (
            .O(N__71323),
            .I(N__71295));
    Span12Mux_h I__17613 (
            .O(N__71320),
            .I(N__71295));
    LocalMux I__17612 (
            .O(N__71315),
            .I(rx_data_1));
    LocalMux I__17611 (
            .O(N__71312),
            .I(rx_data_1));
    Odrv4 I__17610 (
            .O(N__71307),
            .I(rx_data_1));
    Odrv12 I__17609 (
            .O(N__71302),
            .I(rx_data_1));
    Odrv12 I__17608 (
            .O(N__71295),
            .I(rx_data_1));
    CascadeMux I__17607 (
            .O(N__71284),
            .I(N__71280));
    InMux I__17606 (
            .O(N__71283),
            .I(N__71277));
    InMux I__17605 (
            .O(N__71280),
            .I(N__71274));
    LocalMux I__17604 (
            .O(N__71277),
            .I(N__71270));
    LocalMux I__17603 (
            .O(N__71274),
            .I(N__71267));
    CascadeMux I__17602 (
            .O(N__71273),
            .I(N__71262));
    Span4Mux_h I__17601 (
            .O(N__71270),
            .I(N__71259));
    Span4Mux_h I__17600 (
            .O(N__71267),
            .I(N__71256));
    InMux I__17599 (
            .O(N__71266),
            .I(N__71251));
    InMux I__17598 (
            .O(N__71265),
            .I(N__71251));
    InMux I__17597 (
            .O(N__71262),
            .I(N__71248));
    Span4Mux_h I__17596 (
            .O(N__71259),
            .I(N__71245));
    Span4Mux_h I__17595 (
            .O(N__71256),
            .I(N__71240));
    LocalMux I__17594 (
            .O(N__71251),
            .I(N__71240));
    LocalMux I__17593 (
            .O(N__71248),
            .I(\c0.data_in_frame_21_1 ));
    Odrv4 I__17592 (
            .O(N__71245),
            .I(\c0.data_in_frame_21_1 ));
    Odrv4 I__17591 (
            .O(N__71240),
            .I(\c0.data_in_frame_21_1 ));
    ClkMux I__17590 (
            .O(N__71233),
            .I(N__70504));
    ClkMux I__17589 (
            .O(N__71232),
            .I(N__70504));
    ClkMux I__17588 (
            .O(N__71231),
            .I(N__70504));
    ClkMux I__17587 (
            .O(N__71230),
            .I(N__70504));
    ClkMux I__17586 (
            .O(N__71229),
            .I(N__70504));
    ClkMux I__17585 (
            .O(N__71228),
            .I(N__70504));
    ClkMux I__17584 (
            .O(N__71227),
            .I(N__70504));
    ClkMux I__17583 (
            .O(N__71226),
            .I(N__70504));
    ClkMux I__17582 (
            .O(N__71225),
            .I(N__70504));
    ClkMux I__17581 (
            .O(N__71224),
            .I(N__70504));
    ClkMux I__17580 (
            .O(N__71223),
            .I(N__70504));
    ClkMux I__17579 (
            .O(N__71222),
            .I(N__70504));
    ClkMux I__17578 (
            .O(N__71221),
            .I(N__70504));
    ClkMux I__17577 (
            .O(N__71220),
            .I(N__70504));
    ClkMux I__17576 (
            .O(N__71219),
            .I(N__70504));
    ClkMux I__17575 (
            .O(N__71218),
            .I(N__70504));
    ClkMux I__17574 (
            .O(N__71217),
            .I(N__70504));
    ClkMux I__17573 (
            .O(N__71216),
            .I(N__70504));
    ClkMux I__17572 (
            .O(N__71215),
            .I(N__70504));
    ClkMux I__17571 (
            .O(N__71214),
            .I(N__70504));
    ClkMux I__17570 (
            .O(N__71213),
            .I(N__70504));
    ClkMux I__17569 (
            .O(N__71212),
            .I(N__70504));
    ClkMux I__17568 (
            .O(N__71211),
            .I(N__70504));
    ClkMux I__17567 (
            .O(N__71210),
            .I(N__70504));
    ClkMux I__17566 (
            .O(N__71209),
            .I(N__70504));
    ClkMux I__17565 (
            .O(N__71208),
            .I(N__70504));
    ClkMux I__17564 (
            .O(N__71207),
            .I(N__70504));
    ClkMux I__17563 (
            .O(N__71206),
            .I(N__70504));
    ClkMux I__17562 (
            .O(N__71205),
            .I(N__70504));
    ClkMux I__17561 (
            .O(N__71204),
            .I(N__70504));
    ClkMux I__17560 (
            .O(N__71203),
            .I(N__70504));
    ClkMux I__17559 (
            .O(N__71202),
            .I(N__70504));
    ClkMux I__17558 (
            .O(N__71201),
            .I(N__70504));
    ClkMux I__17557 (
            .O(N__71200),
            .I(N__70504));
    ClkMux I__17556 (
            .O(N__71199),
            .I(N__70504));
    ClkMux I__17555 (
            .O(N__71198),
            .I(N__70504));
    ClkMux I__17554 (
            .O(N__71197),
            .I(N__70504));
    ClkMux I__17553 (
            .O(N__71196),
            .I(N__70504));
    ClkMux I__17552 (
            .O(N__71195),
            .I(N__70504));
    ClkMux I__17551 (
            .O(N__71194),
            .I(N__70504));
    ClkMux I__17550 (
            .O(N__71193),
            .I(N__70504));
    ClkMux I__17549 (
            .O(N__71192),
            .I(N__70504));
    ClkMux I__17548 (
            .O(N__71191),
            .I(N__70504));
    ClkMux I__17547 (
            .O(N__71190),
            .I(N__70504));
    ClkMux I__17546 (
            .O(N__71189),
            .I(N__70504));
    ClkMux I__17545 (
            .O(N__71188),
            .I(N__70504));
    ClkMux I__17544 (
            .O(N__71187),
            .I(N__70504));
    ClkMux I__17543 (
            .O(N__71186),
            .I(N__70504));
    ClkMux I__17542 (
            .O(N__71185),
            .I(N__70504));
    ClkMux I__17541 (
            .O(N__71184),
            .I(N__70504));
    ClkMux I__17540 (
            .O(N__71183),
            .I(N__70504));
    ClkMux I__17539 (
            .O(N__71182),
            .I(N__70504));
    ClkMux I__17538 (
            .O(N__71181),
            .I(N__70504));
    ClkMux I__17537 (
            .O(N__71180),
            .I(N__70504));
    ClkMux I__17536 (
            .O(N__71179),
            .I(N__70504));
    ClkMux I__17535 (
            .O(N__71178),
            .I(N__70504));
    ClkMux I__17534 (
            .O(N__71177),
            .I(N__70504));
    ClkMux I__17533 (
            .O(N__71176),
            .I(N__70504));
    ClkMux I__17532 (
            .O(N__71175),
            .I(N__70504));
    ClkMux I__17531 (
            .O(N__71174),
            .I(N__70504));
    ClkMux I__17530 (
            .O(N__71173),
            .I(N__70504));
    ClkMux I__17529 (
            .O(N__71172),
            .I(N__70504));
    ClkMux I__17528 (
            .O(N__71171),
            .I(N__70504));
    ClkMux I__17527 (
            .O(N__71170),
            .I(N__70504));
    ClkMux I__17526 (
            .O(N__71169),
            .I(N__70504));
    ClkMux I__17525 (
            .O(N__71168),
            .I(N__70504));
    ClkMux I__17524 (
            .O(N__71167),
            .I(N__70504));
    ClkMux I__17523 (
            .O(N__71166),
            .I(N__70504));
    ClkMux I__17522 (
            .O(N__71165),
            .I(N__70504));
    ClkMux I__17521 (
            .O(N__71164),
            .I(N__70504));
    ClkMux I__17520 (
            .O(N__71163),
            .I(N__70504));
    ClkMux I__17519 (
            .O(N__71162),
            .I(N__70504));
    ClkMux I__17518 (
            .O(N__71161),
            .I(N__70504));
    ClkMux I__17517 (
            .O(N__71160),
            .I(N__70504));
    ClkMux I__17516 (
            .O(N__71159),
            .I(N__70504));
    ClkMux I__17515 (
            .O(N__71158),
            .I(N__70504));
    ClkMux I__17514 (
            .O(N__71157),
            .I(N__70504));
    ClkMux I__17513 (
            .O(N__71156),
            .I(N__70504));
    ClkMux I__17512 (
            .O(N__71155),
            .I(N__70504));
    ClkMux I__17511 (
            .O(N__71154),
            .I(N__70504));
    ClkMux I__17510 (
            .O(N__71153),
            .I(N__70504));
    ClkMux I__17509 (
            .O(N__71152),
            .I(N__70504));
    ClkMux I__17508 (
            .O(N__71151),
            .I(N__70504));
    ClkMux I__17507 (
            .O(N__71150),
            .I(N__70504));
    ClkMux I__17506 (
            .O(N__71149),
            .I(N__70504));
    ClkMux I__17505 (
            .O(N__71148),
            .I(N__70504));
    ClkMux I__17504 (
            .O(N__71147),
            .I(N__70504));
    ClkMux I__17503 (
            .O(N__71146),
            .I(N__70504));
    ClkMux I__17502 (
            .O(N__71145),
            .I(N__70504));
    ClkMux I__17501 (
            .O(N__71144),
            .I(N__70504));
    ClkMux I__17500 (
            .O(N__71143),
            .I(N__70504));
    ClkMux I__17499 (
            .O(N__71142),
            .I(N__70504));
    ClkMux I__17498 (
            .O(N__71141),
            .I(N__70504));
    ClkMux I__17497 (
            .O(N__71140),
            .I(N__70504));
    ClkMux I__17496 (
            .O(N__71139),
            .I(N__70504));
    ClkMux I__17495 (
            .O(N__71138),
            .I(N__70504));
    ClkMux I__17494 (
            .O(N__71137),
            .I(N__70504));
    ClkMux I__17493 (
            .O(N__71136),
            .I(N__70504));
    ClkMux I__17492 (
            .O(N__71135),
            .I(N__70504));
    ClkMux I__17491 (
            .O(N__71134),
            .I(N__70504));
    ClkMux I__17490 (
            .O(N__71133),
            .I(N__70504));
    ClkMux I__17489 (
            .O(N__71132),
            .I(N__70504));
    ClkMux I__17488 (
            .O(N__71131),
            .I(N__70504));
    ClkMux I__17487 (
            .O(N__71130),
            .I(N__70504));
    ClkMux I__17486 (
            .O(N__71129),
            .I(N__70504));
    ClkMux I__17485 (
            .O(N__71128),
            .I(N__70504));
    ClkMux I__17484 (
            .O(N__71127),
            .I(N__70504));
    ClkMux I__17483 (
            .O(N__71126),
            .I(N__70504));
    ClkMux I__17482 (
            .O(N__71125),
            .I(N__70504));
    ClkMux I__17481 (
            .O(N__71124),
            .I(N__70504));
    ClkMux I__17480 (
            .O(N__71123),
            .I(N__70504));
    ClkMux I__17479 (
            .O(N__71122),
            .I(N__70504));
    ClkMux I__17478 (
            .O(N__71121),
            .I(N__70504));
    ClkMux I__17477 (
            .O(N__71120),
            .I(N__70504));
    ClkMux I__17476 (
            .O(N__71119),
            .I(N__70504));
    ClkMux I__17475 (
            .O(N__71118),
            .I(N__70504));
    ClkMux I__17474 (
            .O(N__71117),
            .I(N__70504));
    ClkMux I__17473 (
            .O(N__71116),
            .I(N__70504));
    ClkMux I__17472 (
            .O(N__71115),
            .I(N__70504));
    ClkMux I__17471 (
            .O(N__71114),
            .I(N__70504));
    ClkMux I__17470 (
            .O(N__71113),
            .I(N__70504));
    ClkMux I__17469 (
            .O(N__71112),
            .I(N__70504));
    ClkMux I__17468 (
            .O(N__71111),
            .I(N__70504));
    ClkMux I__17467 (
            .O(N__71110),
            .I(N__70504));
    ClkMux I__17466 (
            .O(N__71109),
            .I(N__70504));
    ClkMux I__17465 (
            .O(N__71108),
            .I(N__70504));
    ClkMux I__17464 (
            .O(N__71107),
            .I(N__70504));
    ClkMux I__17463 (
            .O(N__71106),
            .I(N__70504));
    ClkMux I__17462 (
            .O(N__71105),
            .I(N__70504));
    ClkMux I__17461 (
            .O(N__71104),
            .I(N__70504));
    ClkMux I__17460 (
            .O(N__71103),
            .I(N__70504));
    ClkMux I__17459 (
            .O(N__71102),
            .I(N__70504));
    ClkMux I__17458 (
            .O(N__71101),
            .I(N__70504));
    ClkMux I__17457 (
            .O(N__71100),
            .I(N__70504));
    ClkMux I__17456 (
            .O(N__71099),
            .I(N__70504));
    ClkMux I__17455 (
            .O(N__71098),
            .I(N__70504));
    ClkMux I__17454 (
            .O(N__71097),
            .I(N__70504));
    ClkMux I__17453 (
            .O(N__71096),
            .I(N__70504));
    ClkMux I__17452 (
            .O(N__71095),
            .I(N__70504));
    ClkMux I__17451 (
            .O(N__71094),
            .I(N__70504));
    ClkMux I__17450 (
            .O(N__71093),
            .I(N__70504));
    ClkMux I__17449 (
            .O(N__71092),
            .I(N__70504));
    ClkMux I__17448 (
            .O(N__71091),
            .I(N__70504));
    ClkMux I__17447 (
            .O(N__71090),
            .I(N__70504));
    ClkMux I__17446 (
            .O(N__71089),
            .I(N__70504));
    ClkMux I__17445 (
            .O(N__71088),
            .I(N__70504));
    ClkMux I__17444 (
            .O(N__71087),
            .I(N__70504));
    ClkMux I__17443 (
            .O(N__71086),
            .I(N__70504));
    ClkMux I__17442 (
            .O(N__71085),
            .I(N__70504));
    ClkMux I__17441 (
            .O(N__71084),
            .I(N__70504));
    ClkMux I__17440 (
            .O(N__71083),
            .I(N__70504));
    ClkMux I__17439 (
            .O(N__71082),
            .I(N__70504));
    ClkMux I__17438 (
            .O(N__71081),
            .I(N__70504));
    ClkMux I__17437 (
            .O(N__71080),
            .I(N__70504));
    ClkMux I__17436 (
            .O(N__71079),
            .I(N__70504));
    ClkMux I__17435 (
            .O(N__71078),
            .I(N__70504));
    ClkMux I__17434 (
            .O(N__71077),
            .I(N__70504));
    ClkMux I__17433 (
            .O(N__71076),
            .I(N__70504));
    ClkMux I__17432 (
            .O(N__71075),
            .I(N__70504));
    ClkMux I__17431 (
            .O(N__71074),
            .I(N__70504));
    ClkMux I__17430 (
            .O(N__71073),
            .I(N__70504));
    ClkMux I__17429 (
            .O(N__71072),
            .I(N__70504));
    ClkMux I__17428 (
            .O(N__71071),
            .I(N__70504));
    ClkMux I__17427 (
            .O(N__71070),
            .I(N__70504));
    ClkMux I__17426 (
            .O(N__71069),
            .I(N__70504));
    ClkMux I__17425 (
            .O(N__71068),
            .I(N__70504));
    ClkMux I__17424 (
            .O(N__71067),
            .I(N__70504));
    ClkMux I__17423 (
            .O(N__71066),
            .I(N__70504));
    ClkMux I__17422 (
            .O(N__71065),
            .I(N__70504));
    ClkMux I__17421 (
            .O(N__71064),
            .I(N__70504));
    ClkMux I__17420 (
            .O(N__71063),
            .I(N__70504));
    ClkMux I__17419 (
            .O(N__71062),
            .I(N__70504));
    ClkMux I__17418 (
            .O(N__71061),
            .I(N__70504));
    ClkMux I__17417 (
            .O(N__71060),
            .I(N__70504));
    ClkMux I__17416 (
            .O(N__71059),
            .I(N__70504));
    ClkMux I__17415 (
            .O(N__71058),
            .I(N__70504));
    ClkMux I__17414 (
            .O(N__71057),
            .I(N__70504));
    ClkMux I__17413 (
            .O(N__71056),
            .I(N__70504));
    ClkMux I__17412 (
            .O(N__71055),
            .I(N__70504));
    ClkMux I__17411 (
            .O(N__71054),
            .I(N__70504));
    ClkMux I__17410 (
            .O(N__71053),
            .I(N__70504));
    ClkMux I__17409 (
            .O(N__71052),
            .I(N__70504));
    ClkMux I__17408 (
            .O(N__71051),
            .I(N__70504));
    ClkMux I__17407 (
            .O(N__71050),
            .I(N__70504));
    ClkMux I__17406 (
            .O(N__71049),
            .I(N__70504));
    ClkMux I__17405 (
            .O(N__71048),
            .I(N__70504));
    ClkMux I__17404 (
            .O(N__71047),
            .I(N__70504));
    ClkMux I__17403 (
            .O(N__71046),
            .I(N__70504));
    ClkMux I__17402 (
            .O(N__71045),
            .I(N__70504));
    ClkMux I__17401 (
            .O(N__71044),
            .I(N__70504));
    ClkMux I__17400 (
            .O(N__71043),
            .I(N__70504));
    ClkMux I__17399 (
            .O(N__71042),
            .I(N__70504));
    ClkMux I__17398 (
            .O(N__71041),
            .I(N__70504));
    ClkMux I__17397 (
            .O(N__71040),
            .I(N__70504));
    ClkMux I__17396 (
            .O(N__71039),
            .I(N__70504));
    ClkMux I__17395 (
            .O(N__71038),
            .I(N__70504));
    ClkMux I__17394 (
            .O(N__71037),
            .I(N__70504));
    ClkMux I__17393 (
            .O(N__71036),
            .I(N__70504));
    ClkMux I__17392 (
            .O(N__71035),
            .I(N__70504));
    ClkMux I__17391 (
            .O(N__71034),
            .I(N__70504));
    ClkMux I__17390 (
            .O(N__71033),
            .I(N__70504));
    ClkMux I__17389 (
            .O(N__71032),
            .I(N__70504));
    ClkMux I__17388 (
            .O(N__71031),
            .I(N__70504));
    ClkMux I__17387 (
            .O(N__71030),
            .I(N__70504));
    ClkMux I__17386 (
            .O(N__71029),
            .I(N__70504));
    ClkMux I__17385 (
            .O(N__71028),
            .I(N__70504));
    ClkMux I__17384 (
            .O(N__71027),
            .I(N__70504));
    ClkMux I__17383 (
            .O(N__71026),
            .I(N__70504));
    ClkMux I__17382 (
            .O(N__71025),
            .I(N__70504));
    ClkMux I__17381 (
            .O(N__71024),
            .I(N__70504));
    ClkMux I__17380 (
            .O(N__71023),
            .I(N__70504));
    ClkMux I__17379 (
            .O(N__71022),
            .I(N__70504));
    ClkMux I__17378 (
            .O(N__71021),
            .I(N__70504));
    ClkMux I__17377 (
            .O(N__71020),
            .I(N__70504));
    ClkMux I__17376 (
            .O(N__71019),
            .I(N__70504));
    ClkMux I__17375 (
            .O(N__71018),
            .I(N__70504));
    ClkMux I__17374 (
            .O(N__71017),
            .I(N__70504));
    ClkMux I__17373 (
            .O(N__71016),
            .I(N__70504));
    ClkMux I__17372 (
            .O(N__71015),
            .I(N__70504));
    ClkMux I__17371 (
            .O(N__71014),
            .I(N__70504));
    ClkMux I__17370 (
            .O(N__71013),
            .I(N__70504));
    ClkMux I__17369 (
            .O(N__71012),
            .I(N__70504));
    ClkMux I__17368 (
            .O(N__71011),
            .I(N__70504));
    ClkMux I__17367 (
            .O(N__71010),
            .I(N__70504));
    ClkMux I__17366 (
            .O(N__71009),
            .I(N__70504));
    ClkMux I__17365 (
            .O(N__71008),
            .I(N__70504));
    ClkMux I__17364 (
            .O(N__71007),
            .I(N__70504));
    ClkMux I__17363 (
            .O(N__71006),
            .I(N__70504));
    ClkMux I__17362 (
            .O(N__71005),
            .I(N__70504));
    ClkMux I__17361 (
            .O(N__71004),
            .I(N__70504));
    ClkMux I__17360 (
            .O(N__71003),
            .I(N__70504));
    ClkMux I__17359 (
            .O(N__71002),
            .I(N__70504));
    ClkMux I__17358 (
            .O(N__71001),
            .I(N__70504));
    ClkMux I__17357 (
            .O(N__71000),
            .I(N__70504));
    ClkMux I__17356 (
            .O(N__70999),
            .I(N__70504));
    ClkMux I__17355 (
            .O(N__70998),
            .I(N__70504));
    ClkMux I__17354 (
            .O(N__70997),
            .I(N__70504));
    ClkMux I__17353 (
            .O(N__70996),
            .I(N__70504));
    ClkMux I__17352 (
            .O(N__70995),
            .I(N__70504));
    ClkMux I__17351 (
            .O(N__70994),
            .I(N__70504));
    ClkMux I__17350 (
            .O(N__70993),
            .I(N__70504));
    ClkMux I__17349 (
            .O(N__70992),
            .I(N__70504));
    ClkMux I__17348 (
            .O(N__70991),
            .I(N__70504));
    GlobalMux I__17347 (
            .O(N__70504),
            .I(N__70501));
    gio2CtrlBuf I__17346 (
            .O(N__70501),
            .I(CLK_c));
    CascadeMux I__17345 (
            .O(N__70498),
            .I(N__70495));
    InMux I__17344 (
            .O(N__70495),
            .I(N__70491));
    InMux I__17343 (
            .O(N__70494),
            .I(N__70488));
    LocalMux I__17342 (
            .O(N__70491),
            .I(N__70485));
    LocalMux I__17341 (
            .O(N__70488),
            .I(N__70482));
    Span4Mux_v I__17340 (
            .O(N__70485),
            .I(N__70478));
    Span4Mux_h I__17339 (
            .O(N__70482),
            .I(N__70475));
    InMux I__17338 (
            .O(N__70481),
            .I(N__70472));
    Odrv4 I__17337 (
            .O(N__70478),
            .I(\c0.n19162 ));
    Odrv4 I__17336 (
            .O(N__70475),
            .I(\c0.n19162 ));
    LocalMux I__17335 (
            .O(N__70472),
            .I(\c0.n19162 ));
    CascadeMux I__17334 (
            .O(N__70465),
            .I(N__70461));
    InMux I__17333 (
            .O(N__70464),
            .I(N__70457));
    InMux I__17332 (
            .O(N__70461),
            .I(N__70451));
    InMux I__17331 (
            .O(N__70460),
            .I(N__70451));
    LocalMux I__17330 (
            .O(N__70457),
            .I(N__70448));
    InMux I__17329 (
            .O(N__70456),
            .I(N__70445));
    LocalMux I__17328 (
            .O(N__70451),
            .I(N__70442));
    Span4Mux_v I__17327 (
            .O(N__70448),
            .I(N__70439));
    LocalMux I__17326 (
            .O(N__70445),
            .I(N__70435));
    Span4Mux_v I__17325 (
            .O(N__70442),
            .I(N__70432));
    Span4Mux_h I__17324 (
            .O(N__70439),
            .I(N__70429));
    InMux I__17323 (
            .O(N__70438),
            .I(N__70425));
    Span4Mux_v I__17322 (
            .O(N__70435),
            .I(N__70420));
    Span4Mux_h I__17321 (
            .O(N__70432),
            .I(N__70420));
    Span4Mux_h I__17320 (
            .O(N__70429),
            .I(N__70417));
    InMux I__17319 (
            .O(N__70428),
            .I(N__70414));
    LocalMux I__17318 (
            .O(N__70425),
            .I(data_in_frame_22_1));
    Odrv4 I__17317 (
            .O(N__70420),
            .I(data_in_frame_22_1));
    Odrv4 I__17316 (
            .O(N__70417),
            .I(data_in_frame_22_1));
    LocalMux I__17315 (
            .O(N__70414),
            .I(data_in_frame_22_1));
    InMux I__17314 (
            .O(N__70405),
            .I(N__70402));
    LocalMux I__17313 (
            .O(N__70402),
            .I(N__70399));
    Span4Mux_v I__17312 (
            .O(N__70399),
            .I(N__70396));
    Span4Mux_h I__17311 (
            .O(N__70396),
            .I(N__70393));
    Odrv4 I__17310 (
            .O(N__70393),
            .I(\c0.n20332 ));
    InMux I__17309 (
            .O(N__70390),
            .I(N__70386));
    InMux I__17308 (
            .O(N__70389),
            .I(N__70383));
    LocalMux I__17307 (
            .O(N__70386),
            .I(N__70379));
    LocalMux I__17306 (
            .O(N__70383),
            .I(N__70376));
    InMux I__17305 (
            .O(N__70382),
            .I(N__70371));
    Span4Mux_v I__17304 (
            .O(N__70379),
            .I(N__70368));
    Span4Mux_h I__17303 (
            .O(N__70376),
            .I(N__70365));
    InMux I__17302 (
            .O(N__70375),
            .I(N__70362));
    InMux I__17301 (
            .O(N__70374),
            .I(N__70359));
    LocalMux I__17300 (
            .O(N__70371),
            .I(N__70354));
    Span4Mux_v I__17299 (
            .O(N__70368),
            .I(N__70354));
    Span4Mux_h I__17298 (
            .O(N__70365),
            .I(N__70351));
    LocalMux I__17297 (
            .O(N__70362),
            .I(N__70348));
    LocalMux I__17296 (
            .O(N__70359),
            .I(data_in_frame_24_1));
    Odrv4 I__17295 (
            .O(N__70354),
            .I(data_in_frame_24_1));
    Odrv4 I__17294 (
            .O(N__70351),
            .I(data_in_frame_24_1));
    Odrv4 I__17293 (
            .O(N__70348),
            .I(data_in_frame_24_1));
    InMux I__17292 (
            .O(N__70339),
            .I(N__70334));
    CascadeMux I__17291 (
            .O(N__70338),
            .I(N__70331));
    InMux I__17290 (
            .O(N__70337),
            .I(N__70328));
    LocalMux I__17289 (
            .O(N__70334),
            .I(N__70325));
    InMux I__17288 (
            .O(N__70331),
            .I(N__70321));
    LocalMux I__17287 (
            .O(N__70328),
            .I(N__70318));
    Span4Mux_h I__17286 (
            .O(N__70325),
            .I(N__70315));
    InMux I__17285 (
            .O(N__70324),
            .I(N__70311));
    LocalMux I__17284 (
            .O(N__70321),
            .I(N__70308));
    Span4Mux_v I__17283 (
            .O(N__70318),
            .I(N__70303));
    Span4Mux_v I__17282 (
            .O(N__70315),
            .I(N__70303));
    InMux I__17281 (
            .O(N__70314),
            .I(N__70300));
    LocalMux I__17280 (
            .O(N__70311),
            .I(data_in_frame_24_3));
    Odrv12 I__17279 (
            .O(N__70308),
            .I(data_in_frame_24_3));
    Odrv4 I__17278 (
            .O(N__70303),
            .I(data_in_frame_24_3));
    LocalMux I__17277 (
            .O(N__70300),
            .I(data_in_frame_24_3));
    CascadeMux I__17276 (
            .O(N__70291),
            .I(\c0.n20332_cascade_ ));
    InMux I__17275 (
            .O(N__70288),
            .I(N__70285));
    LocalMux I__17274 (
            .O(N__70285),
            .I(N__70282));
    Odrv4 I__17273 (
            .O(N__70282),
            .I(\c0.n18413 ));
    InMux I__17272 (
            .O(N__70279),
            .I(N__70276));
    LocalMux I__17271 (
            .O(N__70276),
            .I(N__70273));
    Span4Mux_v I__17270 (
            .O(N__70273),
            .I(N__70270));
    Span4Mux_h I__17269 (
            .O(N__70270),
            .I(N__70267));
    Odrv4 I__17268 (
            .O(N__70267),
            .I(\c0.n36 ));
    InMux I__17267 (
            .O(N__70264),
            .I(N__70261));
    LocalMux I__17266 (
            .O(N__70261),
            .I(N__70258));
    Span4Mux_h I__17265 (
            .O(N__70258),
            .I(N__70254));
    InMux I__17264 (
            .O(N__70257),
            .I(N__70251));
    Span4Mux_v I__17263 (
            .O(N__70254),
            .I(N__70248));
    LocalMux I__17262 (
            .O(N__70251),
            .I(\c0.n20642 ));
    Odrv4 I__17261 (
            .O(N__70248),
            .I(\c0.n20642 ));
    InMux I__17260 (
            .O(N__70243),
            .I(N__70239));
    InMux I__17259 (
            .O(N__70242),
            .I(N__70236));
    LocalMux I__17258 (
            .O(N__70239),
            .I(N__70233));
    LocalMux I__17257 (
            .O(N__70236),
            .I(N__70230));
    Odrv4 I__17256 (
            .O(N__70233),
            .I(\c0.n18525 ));
    Odrv4 I__17255 (
            .O(N__70230),
            .I(\c0.n18525 ));
    CascadeMux I__17254 (
            .O(N__70225),
            .I(N__70221));
    CascadeMux I__17253 (
            .O(N__70224),
            .I(N__70218));
    InMux I__17252 (
            .O(N__70221),
            .I(N__70213));
    InMux I__17251 (
            .O(N__70218),
            .I(N__70213));
    LocalMux I__17250 (
            .O(N__70213),
            .I(N__70210));
    Span4Mux_h I__17249 (
            .O(N__70210),
            .I(N__70205));
    InMux I__17248 (
            .O(N__70209),
            .I(N__70202));
    InMux I__17247 (
            .O(N__70208),
            .I(N__70199));
    Span4Mux_h I__17246 (
            .O(N__70205),
            .I(N__70196));
    LocalMux I__17245 (
            .O(N__70202),
            .I(data_in_frame_24_2));
    LocalMux I__17244 (
            .O(N__70199),
            .I(data_in_frame_24_2));
    Odrv4 I__17243 (
            .O(N__70196),
            .I(data_in_frame_24_2));
    InMux I__17242 (
            .O(N__70189),
            .I(N__70183));
    InMux I__17241 (
            .O(N__70188),
            .I(N__70183));
    LocalMux I__17240 (
            .O(N__70183),
            .I(\c0.n18498 ));
    InMux I__17239 (
            .O(N__70180),
            .I(N__70177));
    LocalMux I__17238 (
            .O(N__70177),
            .I(N__70174));
    Span4Mux_h I__17237 (
            .O(N__70174),
            .I(N__70171));
    Span4Mux_h I__17236 (
            .O(N__70171),
            .I(N__70168));
    Odrv4 I__17235 (
            .O(N__70168),
            .I(\c0.n10_adj_3410 ));
    CascadeMux I__17234 (
            .O(N__70165),
            .I(N__70162));
    InMux I__17233 (
            .O(N__70162),
            .I(N__70158));
    InMux I__17232 (
            .O(N__70161),
            .I(N__70155));
    LocalMux I__17231 (
            .O(N__70158),
            .I(N__70151));
    LocalMux I__17230 (
            .O(N__70155),
            .I(N__70148));
    CascadeMux I__17229 (
            .O(N__70154),
            .I(N__70144));
    Span4Mux_v I__17228 (
            .O(N__70151),
            .I(N__70139));
    Span4Mux_v I__17227 (
            .O(N__70148),
            .I(N__70139));
    InMux I__17226 (
            .O(N__70147),
            .I(N__70134));
    InMux I__17225 (
            .O(N__70144),
            .I(N__70134));
    Span4Mux_h I__17224 (
            .O(N__70139),
            .I(N__70131));
    LocalMux I__17223 (
            .O(N__70134),
            .I(\c0.data_in_frame_20_7 ));
    Odrv4 I__17222 (
            .O(N__70131),
            .I(\c0.data_in_frame_20_7 ));
    InMux I__17221 (
            .O(N__70126),
            .I(N__70120));
    CascadeMux I__17220 (
            .O(N__70125),
            .I(N__70117));
    InMux I__17219 (
            .O(N__70124),
            .I(N__70114));
    InMux I__17218 (
            .O(N__70123),
            .I(N__70111));
    LocalMux I__17217 (
            .O(N__70120),
            .I(N__70108));
    InMux I__17216 (
            .O(N__70117),
            .I(N__70105));
    LocalMux I__17215 (
            .O(N__70114),
            .I(N__70102));
    LocalMux I__17214 (
            .O(N__70111),
            .I(N__70099));
    Span12Mux_h I__17213 (
            .O(N__70108),
            .I(N__70096));
    LocalMux I__17212 (
            .O(N__70105),
            .I(N__70091));
    Span12Mux_v I__17211 (
            .O(N__70102),
            .I(N__70091));
    Odrv4 I__17210 (
            .O(N__70099),
            .I(\c0.data_in_frame_20_6 ));
    Odrv12 I__17209 (
            .O(N__70096),
            .I(\c0.data_in_frame_20_6 ));
    Odrv12 I__17208 (
            .O(N__70091),
            .I(\c0.data_in_frame_20_6 ));
    InMux I__17207 (
            .O(N__70084),
            .I(N__70080));
    InMux I__17206 (
            .O(N__70083),
            .I(N__70077));
    LocalMux I__17205 (
            .O(N__70080),
            .I(N__70074));
    LocalMux I__17204 (
            .O(N__70077),
            .I(\c0.n20576 ));
    Odrv12 I__17203 (
            .O(N__70074),
            .I(\c0.n20576 ));
    InMux I__17202 (
            .O(N__70069),
            .I(N__70066));
    LocalMux I__17201 (
            .O(N__70066),
            .I(\c0.n12_adj_3439 ));
    InMux I__17200 (
            .O(N__70063),
            .I(N__70060));
    LocalMux I__17199 (
            .O(N__70060),
            .I(N__70057));
    Span4Mux_v I__17198 (
            .O(N__70057),
            .I(N__70053));
    InMux I__17197 (
            .O(N__70056),
            .I(N__70050));
    Span4Mux_h I__17196 (
            .O(N__70053),
            .I(N__70045));
    LocalMux I__17195 (
            .O(N__70050),
            .I(N__70045));
    Span4Mux_v I__17194 (
            .O(N__70045),
            .I(N__70041));
    InMux I__17193 (
            .O(N__70044),
            .I(N__70038));
    Sp12to4 I__17192 (
            .O(N__70041),
            .I(N__70032));
    LocalMux I__17191 (
            .O(N__70038),
            .I(N__70032));
    InMux I__17190 (
            .O(N__70037),
            .I(N__70029));
    Span12Mux_h I__17189 (
            .O(N__70032),
            .I(N__70026));
    LocalMux I__17188 (
            .O(N__70029),
            .I(data_in_frame_22_0));
    Odrv12 I__17187 (
            .O(N__70026),
            .I(data_in_frame_22_0));
    InMux I__17186 (
            .O(N__70021),
            .I(N__70018));
    LocalMux I__17185 (
            .O(N__70018),
            .I(N__70013));
    InMux I__17184 (
            .O(N__70017),
            .I(N__70010));
    InMux I__17183 (
            .O(N__70016),
            .I(N__70007));
    Span4Mux_h I__17182 (
            .O(N__70013),
            .I(N__70004));
    LocalMux I__17181 (
            .O(N__70010),
            .I(N__70001));
    LocalMux I__17180 (
            .O(N__70007),
            .I(N__69998));
    Odrv4 I__17179 (
            .O(N__70004),
            .I(\c0.n18415 ));
    Odrv4 I__17178 (
            .O(N__70001),
            .I(\c0.n18415 ));
    Odrv4 I__17177 (
            .O(N__69998),
            .I(\c0.n18415 ));
    CascadeMux I__17176 (
            .O(N__69991),
            .I(\c0.n4_adj_3067_cascade_ ));
    InMux I__17175 (
            .O(N__69988),
            .I(N__69983));
    InMux I__17174 (
            .O(N__69987),
            .I(N__69980));
    InMux I__17173 (
            .O(N__69986),
            .I(N__69977));
    LocalMux I__17172 (
            .O(N__69983),
            .I(N__69974));
    LocalMux I__17171 (
            .O(N__69980),
            .I(N__69971));
    LocalMux I__17170 (
            .O(N__69977),
            .I(N__69968));
    Span4Mux_v I__17169 (
            .O(N__69974),
            .I(N__69961));
    Span4Mux_h I__17168 (
            .O(N__69971),
            .I(N__69958));
    Span4Mux_h I__17167 (
            .O(N__69968),
            .I(N__69955));
    InMux I__17166 (
            .O(N__69967),
            .I(N__69946));
    InMux I__17165 (
            .O(N__69966),
            .I(N__69946));
    InMux I__17164 (
            .O(N__69965),
            .I(N__69946));
    InMux I__17163 (
            .O(N__69964),
            .I(N__69946));
    Odrv4 I__17162 (
            .O(N__69961),
            .I(\c0.n6009 ));
    Odrv4 I__17161 (
            .O(N__69958),
            .I(\c0.n6009 ));
    Odrv4 I__17160 (
            .O(N__69955),
            .I(\c0.n6009 ));
    LocalMux I__17159 (
            .O(N__69946),
            .I(\c0.n6009 ));
    InMux I__17158 (
            .O(N__69937),
            .I(N__69934));
    LocalMux I__17157 (
            .O(N__69934),
            .I(N__69930));
    InMux I__17156 (
            .O(N__69933),
            .I(N__69927));
    Odrv12 I__17155 (
            .O(N__69930),
            .I(\c0.n19369 ));
    LocalMux I__17154 (
            .O(N__69927),
            .I(\c0.n19369 ));
    CascadeMux I__17153 (
            .O(N__69922),
            .I(\c0.n22_adj_3322_cascade_ ));
    InMux I__17152 (
            .O(N__69919),
            .I(N__69913));
    InMux I__17151 (
            .O(N__69918),
            .I(N__69913));
    LocalMux I__17150 (
            .O(N__69913),
            .I(N__69910));
    Odrv4 I__17149 (
            .O(N__69910),
            .I(\c0.n36_adj_3090 ));
    CascadeMux I__17148 (
            .O(N__69907),
            .I(N__69904));
    InMux I__17147 (
            .O(N__69904),
            .I(N__69900));
    InMux I__17146 (
            .O(N__69903),
            .I(N__69897));
    LocalMux I__17145 (
            .O(N__69900),
            .I(N__69893));
    LocalMux I__17144 (
            .O(N__69897),
            .I(N__69890));
    CascadeMux I__17143 (
            .O(N__69896),
            .I(N__69886));
    Span4Mux_h I__17142 (
            .O(N__69893),
            .I(N__69883));
    Span4Mux_v I__17141 (
            .O(N__69890),
            .I(N__69880));
    CascadeMux I__17140 (
            .O(N__69889),
            .I(N__69876));
    InMux I__17139 (
            .O(N__69886),
            .I(N__69873));
    Span4Mux_h I__17138 (
            .O(N__69883),
            .I(N__69870));
    Sp12to4 I__17137 (
            .O(N__69880),
            .I(N__69867));
    InMux I__17136 (
            .O(N__69879),
            .I(N__69862));
    InMux I__17135 (
            .O(N__69876),
            .I(N__69862));
    LocalMux I__17134 (
            .O(N__69873),
            .I(\c0.data_in_frame_21_2 ));
    Odrv4 I__17133 (
            .O(N__69870),
            .I(\c0.data_in_frame_21_2 ));
    Odrv12 I__17132 (
            .O(N__69867),
            .I(\c0.data_in_frame_21_2 ));
    LocalMux I__17131 (
            .O(N__69862),
            .I(\c0.data_in_frame_21_2 ));
    InMux I__17130 (
            .O(N__69853),
            .I(N__69850));
    LocalMux I__17129 (
            .O(N__69850),
            .I(N__69845));
    InMux I__17128 (
            .O(N__69849),
            .I(N__69840));
    InMux I__17127 (
            .O(N__69848),
            .I(N__69840));
    Odrv4 I__17126 (
            .O(N__69845),
            .I(\c0.n29_adj_3383 ));
    LocalMux I__17125 (
            .O(N__69840),
            .I(\c0.n29_adj_3383 ));
    InMux I__17124 (
            .O(N__69835),
            .I(N__69831));
    InMux I__17123 (
            .O(N__69834),
            .I(N__69828));
    LocalMux I__17122 (
            .O(N__69831),
            .I(N__69822));
    LocalMux I__17121 (
            .O(N__69828),
            .I(N__69819));
    InMux I__17120 (
            .O(N__69827),
            .I(N__69812));
    InMux I__17119 (
            .O(N__69826),
            .I(N__69812));
    InMux I__17118 (
            .O(N__69825),
            .I(N__69809));
    Span4Mux_h I__17117 (
            .O(N__69822),
            .I(N__69804));
    Span4Mux_h I__17116 (
            .O(N__69819),
            .I(N__69804));
    InMux I__17115 (
            .O(N__69818),
            .I(N__69801));
    InMux I__17114 (
            .O(N__69817),
            .I(N__69798));
    LocalMux I__17113 (
            .O(N__69812),
            .I(\c0.n20917 ));
    LocalMux I__17112 (
            .O(N__69809),
            .I(\c0.n20917 ));
    Odrv4 I__17111 (
            .O(N__69804),
            .I(\c0.n20917 ));
    LocalMux I__17110 (
            .O(N__69801),
            .I(\c0.n20917 ));
    LocalMux I__17109 (
            .O(N__69798),
            .I(\c0.n20917 ));
    InMux I__17108 (
            .O(N__69787),
            .I(N__69784));
    LocalMux I__17107 (
            .O(N__69784),
            .I(N__69781));
    Span4Mux_h I__17106 (
            .O(N__69781),
            .I(N__69778));
    Span4Mux_v I__17105 (
            .O(N__69778),
            .I(N__69774));
    CascadeMux I__17104 (
            .O(N__69777),
            .I(N__69769));
    Sp12to4 I__17103 (
            .O(N__69774),
            .I(N__69766));
    InMux I__17102 (
            .O(N__69773),
            .I(N__69761));
    InMux I__17101 (
            .O(N__69772),
            .I(N__69761));
    InMux I__17100 (
            .O(N__69769),
            .I(N__69758));
    Span12Mux_s8_h I__17099 (
            .O(N__69766),
            .I(N__69753));
    LocalMux I__17098 (
            .O(N__69761),
            .I(N__69753));
    LocalMux I__17097 (
            .O(N__69758),
            .I(\c0.data_in_frame_20_0 ));
    Odrv12 I__17096 (
            .O(N__69753),
            .I(\c0.data_in_frame_20_0 ));
    InMux I__17095 (
            .O(N__69748),
            .I(N__69739));
    InMux I__17094 (
            .O(N__69747),
            .I(N__69739));
    InMux I__17093 (
            .O(N__69746),
            .I(N__69734));
    InMux I__17092 (
            .O(N__69745),
            .I(N__69734));
    InMux I__17091 (
            .O(N__69744),
            .I(N__69731));
    LocalMux I__17090 (
            .O(N__69739),
            .I(N__69726));
    LocalMux I__17089 (
            .O(N__69734),
            .I(N__69726));
    LocalMux I__17088 (
            .O(N__69731),
            .I(N__69723));
    Span4Mux_v I__17087 (
            .O(N__69726),
            .I(N__69718));
    Span4Mux_v I__17086 (
            .O(N__69723),
            .I(N__69718));
    Odrv4 I__17085 (
            .O(N__69718),
            .I(\c0.n4_adj_3435 ));
    CascadeMux I__17084 (
            .O(N__69715),
            .I(N__69711));
    InMux I__17083 (
            .O(N__69714),
            .I(N__69708));
    InMux I__17082 (
            .O(N__69711),
            .I(N__69704));
    LocalMux I__17081 (
            .O(N__69708),
            .I(N__69701));
    InMux I__17080 (
            .O(N__69707),
            .I(N__69698));
    LocalMux I__17079 (
            .O(N__69704),
            .I(N__69695));
    Odrv4 I__17078 (
            .O(N__69701),
            .I(\c0.n6_adj_3091 ));
    LocalMux I__17077 (
            .O(N__69698),
            .I(\c0.n6_adj_3091 ));
    Odrv12 I__17076 (
            .O(N__69695),
            .I(\c0.n6_adj_3091 ));
    InMux I__17075 (
            .O(N__69688),
            .I(N__69685));
    LocalMux I__17074 (
            .O(N__69685),
            .I(N__69679));
    InMux I__17073 (
            .O(N__69684),
            .I(N__69676));
    InMux I__17072 (
            .O(N__69683),
            .I(N__69673));
    InMux I__17071 (
            .O(N__69682),
            .I(N__69670));
    Odrv12 I__17070 (
            .O(N__69679),
            .I(\c0.n18375 ));
    LocalMux I__17069 (
            .O(N__69676),
            .I(\c0.n18375 ));
    LocalMux I__17068 (
            .O(N__69673),
            .I(\c0.n18375 ));
    LocalMux I__17067 (
            .O(N__69670),
            .I(\c0.n18375 ));
    CascadeMux I__17066 (
            .O(N__69661),
            .I(\c0.n6_adj_3091_cascade_ ));
    InMux I__17065 (
            .O(N__69658),
            .I(N__69653));
    CascadeMux I__17064 (
            .O(N__69657),
            .I(N__69649));
    InMux I__17063 (
            .O(N__69656),
            .I(N__69645));
    LocalMux I__17062 (
            .O(N__69653),
            .I(N__69642));
    InMux I__17061 (
            .O(N__69652),
            .I(N__69637));
    InMux I__17060 (
            .O(N__69649),
            .I(N__69637));
    InMux I__17059 (
            .O(N__69648),
            .I(N__69633));
    LocalMux I__17058 (
            .O(N__69645),
            .I(N__69630));
    Span4Mux_v I__17057 (
            .O(N__69642),
            .I(N__69625));
    LocalMux I__17056 (
            .O(N__69637),
            .I(N__69625));
    InMux I__17055 (
            .O(N__69636),
            .I(N__69622));
    LocalMux I__17054 (
            .O(N__69633),
            .I(N__69619));
    Span4Mux_h I__17053 (
            .O(N__69630),
            .I(N__69614));
    Span4Mux_h I__17052 (
            .O(N__69625),
            .I(N__69614));
    LocalMux I__17051 (
            .O(N__69622),
            .I(\c0.n17900 ));
    Odrv12 I__17050 (
            .O(N__69619),
            .I(\c0.n17900 ));
    Odrv4 I__17049 (
            .O(N__69614),
            .I(\c0.n17900 ));
    CascadeMux I__17048 (
            .O(N__69607),
            .I(N__69603));
    CascadeMux I__17047 (
            .O(N__69606),
            .I(N__69599));
    InMux I__17046 (
            .O(N__69603),
            .I(N__69596));
    CascadeMux I__17045 (
            .O(N__69602),
            .I(N__69592));
    InMux I__17044 (
            .O(N__69599),
            .I(N__69589));
    LocalMux I__17043 (
            .O(N__69596),
            .I(N__69586));
    InMux I__17042 (
            .O(N__69595),
            .I(N__69583));
    InMux I__17041 (
            .O(N__69592),
            .I(N__69580));
    LocalMux I__17040 (
            .O(N__69589),
            .I(N__69577));
    Span4Mux_h I__17039 (
            .O(N__69586),
            .I(N__69572));
    LocalMux I__17038 (
            .O(N__69583),
            .I(N__69572));
    LocalMux I__17037 (
            .O(N__69580),
            .I(\c0.data_in_frame_21_3 ));
    Odrv4 I__17036 (
            .O(N__69577),
            .I(\c0.data_in_frame_21_3 ));
    Odrv4 I__17035 (
            .O(N__69572),
            .I(\c0.data_in_frame_21_3 ));
    InMux I__17034 (
            .O(N__69565),
            .I(N__69561));
    CascadeMux I__17033 (
            .O(N__69564),
            .I(N__69558));
    LocalMux I__17032 (
            .O(N__69561),
            .I(N__69552));
    InMux I__17031 (
            .O(N__69558),
            .I(N__69547));
    InMux I__17030 (
            .O(N__69557),
            .I(N__69547));
    CascadeMux I__17029 (
            .O(N__69556),
            .I(N__69544));
    CascadeMux I__17028 (
            .O(N__69555),
            .I(N__69540));
    Span4Mux_v I__17027 (
            .O(N__69552),
            .I(N__69537));
    LocalMux I__17026 (
            .O(N__69547),
            .I(N__69534));
    InMux I__17025 (
            .O(N__69544),
            .I(N__69529));
    InMux I__17024 (
            .O(N__69543),
            .I(N__69529));
    InMux I__17023 (
            .O(N__69540),
            .I(N__69526));
    Odrv4 I__17022 (
            .O(N__69537),
            .I(\c0.data_in_frame_21_5 ));
    Odrv4 I__17021 (
            .O(N__69534),
            .I(\c0.data_in_frame_21_5 ));
    LocalMux I__17020 (
            .O(N__69529),
            .I(\c0.data_in_frame_21_5 ));
    LocalMux I__17019 (
            .O(N__69526),
            .I(\c0.data_in_frame_21_5 ));
    InMux I__17018 (
            .O(N__69517),
            .I(N__69514));
    LocalMux I__17017 (
            .O(N__69514),
            .I(N__69511));
    Span4Mux_h I__17016 (
            .O(N__69511),
            .I(N__69506));
    InMux I__17015 (
            .O(N__69510),
            .I(N__69501));
    InMux I__17014 (
            .O(N__69509),
            .I(N__69501));
    Odrv4 I__17013 (
            .O(N__69506),
            .I(\c0.n19321 ));
    LocalMux I__17012 (
            .O(N__69501),
            .I(\c0.n19321 ));
    InMux I__17011 (
            .O(N__69496),
            .I(N__69493));
    LocalMux I__17010 (
            .O(N__69493),
            .I(N__69489));
    InMux I__17009 (
            .O(N__69492),
            .I(N__69486));
    Span4Mux_h I__17008 (
            .O(N__69489),
            .I(N__69483));
    LocalMux I__17007 (
            .O(N__69486),
            .I(N__69480));
    Odrv4 I__17006 (
            .O(N__69483),
            .I(\c0.n12037 ));
    Odrv12 I__17005 (
            .O(N__69480),
            .I(\c0.n12037 ));
    CascadeMux I__17004 (
            .O(N__69475),
            .I(N__69472));
    InMux I__17003 (
            .O(N__69472),
            .I(N__69469));
    LocalMux I__17002 (
            .O(N__69469),
            .I(N__69466));
    Span4Mux_h I__17001 (
            .O(N__69466),
            .I(N__69462));
    CascadeMux I__17000 (
            .O(N__69465),
            .I(N__69459));
    Span4Mux_v I__16999 (
            .O(N__69462),
            .I(N__69455));
    InMux I__16998 (
            .O(N__69459),
            .I(N__69450));
    InMux I__16997 (
            .O(N__69458),
            .I(N__69450));
    Odrv4 I__16996 (
            .O(N__69455),
            .I(data_in_frame_19_7));
    LocalMux I__16995 (
            .O(N__69450),
            .I(data_in_frame_19_7));
    InMux I__16994 (
            .O(N__69445),
            .I(N__69439));
    CascadeMux I__16993 (
            .O(N__69444),
            .I(N__69432));
    InMux I__16992 (
            .O(N__69443),
            .I(N__69429));
    InMux I__16991 (
            .O(N__69442),
            .I(N__69426));
    LocalMux I__16990 (
            .O(N__69439),
            .I(N__69418));
    InMux I__16989 (
            .O(N__69438),
            .I(N__69415));
    CascadeMux I__16988 (
            .O(N__69437),
            .I(N__69411));
    InMux I__16987 (
            .O(N__69436),
            .I(N__69405));
    InMux I__16986 (
            .O(N__69435),
            .I(N__69402));
    InMux I__16985 (
            .O(N__69432),
            .I(N__69399));
    LocalMux I__16984 (
            .O(N__69429),
            .I(N__69396));
    LocalMux I__16983 (
            .O(N__69426),
            .I(N__69393));
    InMux I__16982 (
            .O(N__69425),
            .I(N__69390));
    InMux I__16981 (
            .O(N__69424),
            .I(N__69385));
    InMux I__16980 (
            .O(N__69423),
            .I(N__69385));
    InMux I__16979 (
            .O(N__69422),
            .I(N__69382));
    InMux I__16978 (
            .O(N__69421),
            .I(N__69377));
    Span4Mux_h I__16977 (
            .O(N__69418),
            .I(N__69371));
    LocalMux I__16976 (
            .O(N__69415),
            .I(N__69371));
    InMux I__16975 (
            .O(N__69414),
            .I(N__69364));
    InMux I__16974 (
            .O(N__69411),
            .I(N__69364));
    InMux I__16973 (
            .O(N__69410),
            .I(N__69364));
    InMux I__16972 (
            .O(N__69409),
            .I(N__69360));
    InMux I__16971 (
            .O(N__69408),
            .I(N__69357));
    LocalMux I__16970 (
            .O(N__69405),
            .I(N__69352));
    LocalMux I__16969 (
            .O(N__69402),
            .I(N__69352));
    LocalMux I__16968 (
            .O(N__69399),
            .I(N__69349));
    Span4Mux_v I__16967 (
            .O(N__69396),
            .I(N__69342));
    Span4Mux_v I__16966 (
            .O(N__69393),
            .I(N__69342));
    LocalMux I__16965 (
            .O(N__69390),
            .I(N__69342));
    LocalMux I__16964 (
            .O(N__69385),
            .I(N__69339));
    LocalMux I__16963 (
            .O(N__69382),
            .I(N__69336));
    InMux I__16962 (
            .O(N__69381),
            .I(N__69331));
    InMux I__16961 (
            .O(N__69380),
            .I(N__69331));
    LocalMux I__16960 (
            .O(N__69377),
            .I(N__69328));
    InMux I__16959 (
            .O(N__69376),
            .I(N__69325));
    Span4Mux_v I__16958 (
            .O(N__69371),
            .I(N__69320));
    LocalMux I__16957 (
            .O(N__69364),
            .I(N__69320));
    CascadeMux I__16956 (
            .O(N__69363),
            .I(N__69317));
    LocalMux I__16955 (
            .O(N__69360),
            .I(N__69311));
    LocalMux I__16954 (
            .O(N__69357),
            .I(N__69308));
    Span4Mux_v I__16953 (
            .O(N__69352),
            .I(N__69301));
    Span4Mux_h I__16952 (
            .O(N__69349),
            .I(N__69301));
    Span4Mux_h I__16951 (
            .O(N__69342),
            .I(N__69301));
    Span4Mux_v I__16950 (
            .O(N__69339),
            .I(N__69298));
    Span4Mux_h I__16949 (
            .O(N__69336),
            .I(N__69293));
    LocalMux I__16948 (
            .O(N__69331),
            .I(N__69293));
    Span4Mux_h I__16947 (
            .O(N__69328),
            .I(N__69288));
    LocalMux I__16946 (
            .O(N__69325),
            .I(N__69288));
    Span4Mux_h I__16945 (
            .O(N__69320),
            .I(N__69284));
    InMux I__16944 (
            .O(N__69317),
            .I(N__69279));
    InMux I__16943 (
            .O(N__69316),
            .I(N__69279));
    InMux I__16942 (
            .O(N__69315),
            .I(N__69274));
    InMux I__16941 (
            .O(N__69314),
            .I(N__69271));
    Span4Mux_h I__16940 (
            .O(N__69311),
            .I(N__69264));
    Span4Mux_v I__16939 (
            .O(N__69308),
            .I(N__69264));
    Span4Mux_v I__16938 (
            .O(N__69301),
            .I(N__69264));
    Span4Mux_v I__16937 (
            .O(N__69298),
            .I(N__69261));
    Span4Mux_h I__16936 (
            .O(N__69293),
            .I(N__69256));
    Span4Mux_v I__16935 (
            .O(N__69288),
            .I(N__69256));
    InMux I__16934 (
            .O(N__69287),
            .I(N__69253));
    Span4Mux_v I__16933 (
            .O(N__69284),
            .I(N__69248));
    LocalMux I__16932 (
            .O(N__69279),
            .I(N__69248));
    InMux I__16931 (
            .O(N__69278),
            .I(N__69242));
    InMux I__16930 (
            .O(N__69277),
            .I(N__69242));
    LocalMux I__16929 (
            .O(N__69274),
            .I(N__69239));
    LocalMux I__16928 (
            .O(N__69271),
            .I(N__69236));
    Span4Mux_v I__16927 (
            .O(N__69264),
            .I(N__69233));
    Span4Mux_v I__16926 (
            .O(N__69261),
            .I(N__69228));
    Span4Mux_h I__16925 (
            .O(N__69256),
            .I(N__69228));
    LocalMux I__16924 (
            .O(N__69253),
            .I(N__69225));
    Span4Mux_h I__16923 (
            .O(N__69248),
            .I(N__69222));
    InMux I__16922 (
            .O(N__69247),
            .I(N__69219));
    LocalMux I__16921 (
            .O(N__69242),
            .I(N__69212));
    Span4Mux_h I__16920 (
            .O(N__69239),
            .I(N__69207));
    Span4Mux_h I__16919 (
            .O(N__69236),
            .I(N__69207));
    Span4Mux_h I__16918 (
            .O(N__69233),
            .I(N__69204));
    Span4Mux_v I__16917 (
            .O(N__69228),
            .I(N__69201));
    Span4Mux_h I__16916 (
            .O(N__69225),
            .I(N__69194));
    Span4Mux_h I__16915 (
            .O(N__69222),
            .I(N__69194));
    LocalMux I__16914 (
            .O(N__69219),
            .I(N__69194));
    InMux I__16913 (
            .O(N__69218),
            .I(N__69189));
    InMux I__16912 (
            .O(N__69217),
            .I(N__69189));
    InMux I__16911 (
            .O(N__69216),
            .I(N__69184));
    InMux I__16910 (
            .O(N__69215),
            .I(N__69184));
    Odrv12 I__16909 (
            .O(N__69212),
            .I(rx_data_3));
    Odrv4 I__16908 (
            .O(N__69207),
            .I(rx_data_3));
    Odrv4 I__16907 (
            .O(N__69204),
            .I(rx_data_3));
    Odrv4 I__16906 (
            .O(N__69201),
            .I(rx_data_3));
    Odrv4 I__16905 (
            .O(N__69194),
            .I(rx_data_3));
    LocalMux I__16904 (
            .O(N__69189),
            .I(rx_data_3));
    LocalMux I__16903 (
            .O(N__69184),
            .I(rx_data_3));
    InMux I__16902 (
            .O(N__69169),
            .I(N__69164));
    InMux I__16901 (
            .O(N__69168),
            .I(N__69161));
    InMux I__16900 (
            .O(N__69167),
            .I(N__69158));
    LocalMux I__16899 (
            .O(N__69164),
            .I(N__69155));
    LocalMux I__16898 (
            .O(N__69161),
            .I(N__69152));
    LocalMux I__16897 (
            .O(N__69158),
            .I(N__69147));
    Span4Mux_h I__16896 (
            .O(N__69155),
            .I(N__69143));
    Span4Mux_v I__16895 (
            .O(N__69152),
            .I(N__69140));
    InMux I__16894 (
            .O(N__69151),
            .I(N__69133));
    InMux I__16893 (
            .O(N__69150),
            .I(N__69133));
    Span4Mux_h I__16892 (
            .O(N__69147),
            .I(N__69130));
    InMux I__16891 (
            .O(N__69146),
            .I(N__69127));
    Span4Mux_v I__16890 (
            .O(N__69143),
            .I(N__69124));
    Sp12to4 I__16889 (
            .O(N__69140),
            .I(N__69121));
    InMux I__16888 (
            .O(N__69139),
            .I(N__69116));
    InMux I__16887 (
            .O(N__69138),
            .I(N__69116));
    LocalMux I__16886 (
            .O(N__69133),
            .I(N__69111));
    Span4Mux_v I__16885 (
            .O(N__69130),
            .I(N__69111));
    LocalMux I__16884 (
            .O(N__69127),
            .I(N__69108));
    Span4Mux_v I__16883 (
            .O(N__69124),
            .I(N__69105));
    Span12Mux_s10_v I__16882 (
            .O(N__69121),
            .I(N__69102));
    LocalMux I__16881 (
            .O(N__69116),
            .I(N__69097));
    Span4Mux_h I__16880 (
            .O(N__69111),
            .I(N__69097));
    Span4Mux_h I__16879 (
            .O(N__69108),
            .I(N__69092));
    Span4Mux_h I__16878 (
            .O(N__69105),
            .I(N__69092));
    Span12Mux_v I__16877 (
            .O(N__69102),
            .I(N__69089));
    Odrv4 I__16876 (
            .O(N__69097),
            .I(n19128));
    Odrv4 I__16875 (
            .O(N__69092),
            .I(n19128));
    Odrv12 I__16874 (
            .O(N__69089),
            .I(n19128));
    InMux I__16873 (
            .O(N__69082),
            .I(N__69071));
    InMux I__16872 (
            .O(N__69081),
            .I(N__69071));
    InMux I__16871 (
            .O(N__69080),
            .I(N__69071));
    InMux I__16870 (
            .O(N__69079),
            .I(N__69066));
    InMux I__16869 (
            .O(N__69078),
            .I(N__69066));
    LocalMux I__16868 (
            .O(N__69071),
            .I(N__69063));
    LocalMux I__16867 (
            .O(N__69066),
            .I(N__69060));
    Span4Mux_v I__16866 (
            .O(N__69063),
            .I(N__69057));
    Span4Mux_v I__16865 (
            .O(N__69060),
            .I(N__69050));
    Span4Mux_v I__16864 (
            .O(N__69057),
            .I(N__69050));
    InMux I__16863 (
            .O(N__69056),
            .I(N__69045));
    InMux I__16862 (
            .O(N__69055),
            .I(N__69045));
    Odrv4 I__16861 (
            .O(N__69050),
            .I(data_in_frame_19_3));
    LocalMux I__16860 (
            .O(N__69045),
            .I(data_in_frame_19_3));
    InMux I__16859 (
            .O(N__69040),
            .I(N__69037));
    LocalMux I__16858 (
            .O(N__69037),
            .I(N__69032));
    InMux I__16857 (
            .O(N__69036),
            .I(N__69026));
    InMux I__16856 (
            .O(N__69035),
            .I(N__69026));
    Span4Mux_v I__16855 (
            .O(N__69032),
            .I(N__69019));
    InMux I__16854 (
            .O(N__69031),
            .I(N__69016));
    LocalMux I__16853 (
            .O(N__69026),
            .I(N__69008));
    CascadeMux I__16852 (
            .O(N__69025),
            .I(N__69003));
    InMux I__16851 (
            .O(N__69024),
            .I(N__68998));
    CascadeMux I__16850 (
            .O(N__69023),
            .I(N__68995));
    InMux I__16849 (
            .O(N__69022),
            .I(N__68991));
    Span4Mux_h I__16848 (
            .O(N__69019),
            .I(N__68986));
    LocalMux I__16847 (
            .O(N__69016),
            .I(N__68986));
    InMux I__16846 (
            .O(N__69015),
            .I(N__68981));
    InMux I__16845 (
            .O(N__69014),
            .I(N__68981));
    InMux I__16844 (
            .O(N__69013),
            .I(N__68977));
    InMux I__16843 (
            .O(N__69012),
            .I(N__68974));
    InMux I__16842 (
            .O(N__69011),
            .I(N__68970));
    Span4Mux_v I__16841 (
            .O(N__69008),
            .I(N__68967));
    InMux I__16840 (
            .O(N__69007),
            .I(N__68964));
    InMux I__16839 (
            .O(N__69006),
            .I(N__68961));
    InMux I__16838 (
            .O(N__69003),
            .I(N__68956));
    InMux I__16837 (
            .O(N__69002),
            .I(N__68956));
    InMux I__16836 (
            .O(N__69001),
            .I(N__68953));
    LocalMux I__16835 (
            .O(N__68998),
            .I(N__68950));
    InMux I__16834 (
            .O(N__68995),
            .I(N__68945));
    InMux I__16833 (
            .O(N__68994),
            .I(N__68945));
    LocalMux I__16832 (
            .O(N__68991),
            .I(N__68938));
    Span4Mux_v I__16831 (
            .O(N__68986),
            .I(N__68938));
    LocalMux I__16830 (
            .O(N__68981),
            .I(N__68938));
    InMux I__16829 (
            .O(N__68980),
            .I(N__68935));
    LocalMux I__16828 (
            .O(N__68977),
            .I(N__68932));
    LocalMux I__16827 (
            .O(N__68974),
            .I(N__68929));
    CascadeMux I__16826 (
            .O(N__68973),
            .I(N__68924));
    LocalMux I__16825 (
            .O(N__68970),
            .I(N__68920));
    Span4Mux_h I__16824 (
            .O(N__68967),
            .I(N__68917));
    LocalMux I__16823 (
            .O(N__68964),
            .I(N__68912));
    LocalMux I__16822 (
            .O(N__68961),
            .I(N__68912));
    LocalMux I__16821 (
            .O(N__68956),
            .I(N__68909));
    LocalMux I__16820 (
            .O(N__68953),
            .I(N__68904));
    Span4Mux_v I__16819 (
            .O(N__68950),
            .I(N__68904));
    LocalMux I__16818 (
            .O(N__68945),
            .I(N__68898));
    Span4Mux_v I__16817 (
            .O(N__68938),
            .I(N__68898));
    LocalMux I__16816 (
            .O(N__68935),
            .I(N__68895));
    Span4Mux_v I__16815 (
            .O(N__68932),
            .I(N__68890));
    Span4Mux_h I__16814 (
            .O(N__68929),
            .I(N__68890));
    InMux I__16813 (
            .O(N__68928),
            .I(N__68887));
    InMux I__16812 (
            .O(N__68927),
            .I(N__68882));
    InMux I__16811 (
            .O(N__68924),
            .I(N__68882));
    InMux I__16810 (
            .O(N__68923),
            .I(N__68879));
    Span4Mux_h I__16809 (
            .O(N__68920),
            .I(N__68872));
    Span4Mux_v I__16808 (
            .O(N__68917),
            .I(N__68872));
    Span4Mux_v I__16807 (
            .O(N__68912),
            .I(N__68872));
    Span4Mux_h I__16806 (
            .O(N__68909),
            .I(N__68867));
    Span4Mux_v I__16805 (
            .O(N__68904),
            .I(N__68867));
    InMux I__16804 (
            .O(N__68903),
            .I(N__68863));
    Span4Mux_h I__16803 (
            .O(N__68898),
            .I(N__68860));
    Span4Mux_v I__16802 (
            .O(N__68895),
            .I(N__68855));
    Span4Mux_v I__16801 (
            .O(N__68890),
            .I(N__68855));
    LocalMux I__16800 (
            .O(N__68887),
            .I(N__68850));
    LocalMux I__16799 (
            .O(N__68882),
            .I(N__68845));
    LocalMux I__16798 (
            .O(N__68879),
            .I(N__68845));
    Span4Mux_v I__16797 (
            .O(N__68872),
            .I(N__68840));
    Span4Mux_v I__16796 (
            .O(N__68867),
            .I(N__68837));
    InMux I__16795 (
            .O(N__68866),
            .I(N__68834));
    LocalMux I__16794 (
            .O(N__68863),
            .I(N__68827));
    Span4Mux_v I__16793 (
            .O(N__68860),
            .I(N__68827));
    Span4Mux_v I__16792 (
            .O(N__68855),
            .I(N__68827));
    CascadeMux I__16791 (
            .O(N__68854),
            .I(N__68821));
    InMux I__16790 (
            .O(N__68853),
            .I(N__68818));
    Span4Mux_v I__16789 (
            .O(N__68850),
            .I(N__68813));
    Span4Mux_v I__16788 (
            .O(N__68845),
            .I(N__68813));
    InMux I__16787 (
            .O(N__68844),
            .I(N__68808));
    InMux I__16786 (
            .O(N__68843),
            .I(N__68808));
    Span4Mux_h I__16785 (
            .O(N__68840),
            .I(N__68803));
    Span4Mux_h I__16784 (
            .O(N__68837),
            .I(N__68803));
    LocalMux I__16783 (
            .O(N__68834),
            .I(N__68800));
    Span4Mux_h I__16782 (
            .O(N__68827),
            .I(N__68797));
    InMux I__16781 (
            .O(N__68826),
            .I(N__68794));
    InMux I__16780 (
            .O(N__68825),
            .I(N__68789));
    InMux I__16779 (
            .O(N__68824),
            .I(N__68789));
    InMux I__16778 (
            .O(N__68821),
            .I(N__68786));
    LocalMux I__16777 (
            .O(N__68818),
            .I(N__68781));
    Span4Mux_h I__16776 (
            .O(N__68813),
            .I(N__68781));
    LocalMux I__16775 (
            .O(N__68808),
            .I(N__68776));
    Span4Mux_h I__16774 (
            .O(N__68803),
            .I(N__68776));
    Span4Mux_v I__16773 (
            .O(N__68800),
            .I(N__68771));
    Span4Mux_h I__16772 (
            .O(N__68797),
            .I(N__68771));
    LocalMux I__16771 (
            .O(N__68794),
            .I(rx_data_6));
    LocalMux I__16770 (
            .O(N__68789),
            .I(rx_data_6));
    LocalMux I__16769 (
            .O(N__68786),
            .I(rx_data_6));
    Odrv4 I__16768 (
            .O(N__68781),
            .I(rx_data_6));
    Odrv4 I__16767 (
            .O(N__68776),
            .I(rx_data_6));
    Odrv4 I__16766 (
            .O(N__68771),
            .I(rx_data_6));
    CascadeMux I__16765 (
            .O(N__68758),
            .I(N__68755));
    InMux I__16764 (
            .O(N__68755),
            .I(N__68752));
    LocalMux I__16763 (
            .O(N__68752),
            .I(N__68747));
    CascadeMux I__16762 (
            .O(N__68751),
            .I(N__68741));
    InMux I__16761 (
            .O(N__68750),
            .I(N__68737));
    Span4Mux_v I__16760 (
            .O(N__68747),
            .I(N__68734));
    InMux I__16759 (
            .O(N__68746),
            .I(N__68731));
    InMux I__16758 (
            .O(N__68745),
            .I(N__68728));
    InMux I__16757 (
            .O(N__68744),
            .I(N__68719));
    InMux I__16756 (
            .O(N__68741),
            .I(N__68716));
    InMux I__16755 (
            .O(N__68740),
            .I(N__68713));
    LocalMux I__16754 (
            .O(N__68737),
            .I(N__68708));
    Span4Mux_h I__16753 (
            .O(N__68734),
            .I(N__68701));
    LocalMux I__16752 (
            .O(N__68731),
            .I(N__68701));
    LocalMux I__16751 (
            .O(N__68728),
            .I(N__68701));
    InMux I__16750 (
            .O(N__68727),
            .I(N__68698));
    InMux I__16749 (
            .O(N__68726),
            .I(N__68695));
    InMux I__16748 (
            .O(N__68725),
            .I(N__68692));
    CascadeMux I__16747 (
            .O(N__68724),
            .I(N__68688));
    InMux I__16746 (
            .O(N__68723),
            .I(N__68683));
    InMux I__16745 (
            .O(N__68722),
            .I(N__68683));
    LocalMux I__16744 (
            .O(N__68719),
            .I(N__68675));
    LocalMux I__16743 (
            .O(N__68716),
            .I(N__68675));
    LocalMux I__16742 (
            .O(N__68713),
            .I(N__68675));
    InMux I__16741 (
            .O(N__68712),
            .I(N__68671));
    InMux I__16740 (
            .O(N__68711),
            .I(N__68668));
    Span4Mux_v I__16739 (
            .O(N__68708),
            .I(N__68657));
    Span4Mux_v I__16738 (
            .O(N__68701),
            .I(N__68657));
    LocalMux I__16737 (
            .O(N__68698),
            .I(N__68657));
    LocalMux I__16736 (
            .O(N__68695),
            .I(N__68657));
    LocalMux I__16735 (
            .O(N__68692),
            .I(N__68657));
    InMux I__16734 (
            .O(N__68691),
            .I(N__68652));
    InMux I__16733 (
            .O(N__68688),
            .I(N__68649));
    LocalMux I__16732 (
            .O(N__68683),
            .I(N__68641));
    InMux I__16731 (
            .O(N__68682),
            .I(N__68638));
    Span4Mux_v I__16730 (
            .O(N__68675),
            .I(N__68635));
    InMux I__16729 (
            .O(N__68674),
            .I(N__68632));
    LocalMux I__16728 (
            .O(N__68671),
            .I(N__68629));
    LocalMux I__16727 (
            .O(N__68668),
            .I(N__68626));
    Span4Mux_v I__16726 (
            .O(N__68657),
            .I(N__68623));
    InMux I__16725 (
            .O(N__68656),
            .I(N__68619));
    InMux I__16724 (
            .O(N__68655),
            .I(N__68616));
    LocalMux I__16723 (
            .O(N__68652),
            .I(N__68613));
    LocalMux I__16722 (
            .O(N__68649),
            .I(N__68609));
    InMux I__16721 (
            .O(N__68648),
            .I(N__68604));
    InMux I__16720 (
            .O(N__68647),
            .I(N__68604));
    InMux I__16719 (
            .O(N__68646),
            .I(N__68601));
    InMux I__16718 (
            .O(N__68645),
            .I(N__68598));
    InMux I__16717 (
            .O(N__68644),
            .I(N__68595));
    Span4Mux_h I__16716 (
            .O(N__68641),
            .I(N__68590));
    LocalMux I__16715 (
            .O(N__68638),
            .I(N__68587));
    Span4Mux_h I__16714 (
            .O(N__68635),
            .I(N__68584));
    LocalMux I__16713 (
            .O(N__68632),
            .I(N__68581));
    Span4Mux_h I__16712 (
            .O(N__68629),
            .I(N__68576));
    Span4Mux_h I__16711 (
            .O(N__68626),
            .I(N__68576));
    Span4Mux_h I__16710 (
            .O(N__68623),
            .I(N__68573));
    InMux I__16709 (
            .O(N__68622),
            .I(N__68570));
    LocalMux I__16708 (
            .O(N__68619),
            .I(N__68565));
    LocalMux I__16707 (
            .O(N__68616),
            .I(N__68565));
    Span4Mux_h I__16706 (
            .O(N__68613),
            .I(N__68562));
    InMux I__16705 (
            .O(N__68612),
            .I(N__68559));
    Span4Mux_h I__16704 (
            .O(N__68609),
            .I(N__68554));
    LocalMux I__16703 (
            .O(N__68604),
            .I(N__68554));
    LocalMux I__16702 (
            .O(N__68601),
            .I(N__68546));
    LocalMux I__16701 (
            .O(N__68598),
            .I(N__68546));
    LocalMux I__16700 (
            .O(N__68595),
            .I(N__68546));
    InMux I__16699 (
            .O(N__68594),
            .I(N__68543));
    InMux I__16698 (
            .O(N__68593),
            .I(N__68540));
    Span4Mux_v I__16697 (
            .O(N__68590),
            .I(N__68535));
    Span4Mux_h I__16696 (
            .O(N__68587),
            .I(N__68535));
    Sp12to4 I__16695 (
            .O(N__68584),
            .I(N__68532));
    Span4Mux_h I__16694 (
            .O(N__68581),
            .I(N__68529));
    Span4Mux_v I__16693 (
            .O(N__68576),
            .I(N__68526));
    Span4Mux_v I__16692 (
            .O(N__68573),
            .I(N__68523));
    LocalMux I__16691 (
            .O(N__68570),
            .I(N__68518));
    Sp12to4 I__16690 (
            .O(N__68565),
            .I(N__68515));
    Span4Mux_h I__16689 (
            .O(N__68562),
            .I(N__68512));
    LocalMux I__16688 (
            .O(N__68559),
            .I(N__68509));
    Span4Mux_v I__16687 (
            .O(N__68554),
            .I(N__68506));
    InMux I__16686 (
            .O(N__68553),
            .I(N__68503));
    Span4Mux_v I__16685 (
            .O(N__68546),
            .I(N__68500));
    LocalMux I__16684 (
            .O(N__68543),
            .I(N__68495));
    LocalMux I__16683 (
            .O(N__68540),
            .I(N__68495));
    Sp12to4 I__16682 (
            .O(N__68535),
            .I(N__68492));
    Span12Mux_h I__16681 (
            .O(N__68532),
            .I(N__68489));
    Span4Mux_v I__16680 (
            .O(N__68529),
            .I(N__68484));
    Span4Mux_v I__16679 (
            .O(N__68526),
            .I(N__68484));
    Sp12to4 I__16678 (
            .O(N__68523),
            .I(N__68481));
    InMux I__16677 (
            .O(N__68522),
            .I(N__68476));
    InMux I__16676 (
            .O(N__68521),
            .I(N__68476));
    Span4Mux_v I__16675 (
            .O(N__68518),
            .I(N__68473));
    Span12Mux_v I__16674 (
            .O(N__68515),
            .I(N__68470));
    Span4Mux_v I__16673 (
            .O(N__68512),
            .I(N__68463));
    Span4Mux_v I__16672 (
            .O(N__68509),
            .I(N__68463));
    Span4Mux_v I__16671 (
            .O(N__68506),
            .I(N__68463));
    LocalMux I__16670 (
            .O(N__68503),
            .I(N__68456));
    Span4Mux_v I__16669 (
            .O(N__68500),
            .I(N__68456));
    Span4Mux_h I__16668 (
            .O(N__68495),
            .I(N__68456));
    Span12Mux_v I__16667 (
            .O(N__68492),
            .I(N__68447));
    Span12Mux_v I__16666 (
            .O(N__68489),
            .I(N__68447));
    Sp12to4 I__16665 (
            .O(N__68484),
            .I(N__68447));
    Span12Mux_s6_h I__16664 (
            .O(N__68481),
            .I(N__68447));
    LocalMux I__16663 (
            .O(N__68476),
            .I(rx_data_2));
    Odrv4 I__16662 (
            .O(N__68473),
            .I(rx_data_2));
    Odrv12 I__16661 (
            .O(N__68470),
            .I(rx_data_2));
    Odrv4 I__16660 (
            .O(N__68463),
            .I(rx_data_2));
    Odrv4 I__16659 (
            .O(N__68456),
            .I(rx_data_2));
    Odrv12 I__16658 (
            .O(N__68447),
            .I(rx_data_2));
    InMux I__16657 (
            .O(N__68434),
            .I(N__68431));
    LocalMux I__16656 (
            .O(N__68431),
            .I(N__68425));
    InMux I__16655 (
            .O(N__68430),
            .I(N__68422));
    InMux I__16654 (
            .O(N__68429),
            .I(N__68419));
    InMux I__16653 (
            .O(N__68428),
            .I(N__68416));
    Span4Mux_v I__16652 (
            .O(N__68425),
            .I(N__68413));
    LocalMux I__16651 (
            .O(N__68422),
            .I(N__68410));
    LocalMux I__16650 (
            .O(N__68419),
            .I(N__68405));
    LocalMux I__16649 (
            .O(N__68416),
            .I(N__68405));
    Span4Mux_h I__16648 (
            .O(N__68413),
            .I(N__68398));
    Span4Mux_v I__16647 (
            .O(N__68410),
            .I(N__68398));
    Span4Mux_h I__16646 (
            .O(N__68405),
            .I(N__68398));
    Span4Mux_v I__16645 (
            .O(N__68398),
            .I(N__68395));
    Odrv4 I__16644 (
            .O(N__68395),
            .I(\c0.n19474 ));
    CascadeMux I__16643 (
            .O(N__68392),
            .I(N__68388));
    CascadeMux I__16642 (
            .O(N__68391),
            .I(N__68385));
    InMux I__16641 (
            .O(N__68388),
            .I(N__68378));
    InMux I__16640 (
            .O(N__68385),
            .I(N__68378));
    InMux I__16639 (
            .O(N__68384),
            .I(N__68375));
    InMux I__16638 (
            .O(N__68383),
            .I(N__68371));
    LocalMux I__16637 (
            .O(N__68378),
            .I(N__68368));
    LocalMux I__16636 (
            .O(N__68375),
            .I(N__68365));
    InMux I__16635 (
            .O(N__68374),
            .I(N__68361));
    LocalMux I__16634 (
            .O(N__68371),
            .I(N__68356));
    Span4Mux_v I__16633 (
            .O(N__68368),
            .I(N__68356));
    Span4Mux_v I__16632 (
            .O(N__68365),
            .I(N__68352));
    CascadeMux I__16631 (
            .O(N__68364),
            .I(N__68349));
    LocalMux I__16630 (
            .O(N__68361),
            .I(N__68345));
    Span4Mux_v I__16629 (
            .O(N__68356),
            .I(N__68342));
    InMux I__16628 (
            .O(N__68355),
            .I(N__68339));
    Span4Mux_h I__16627 (
            .O(N__68352),
            .I(N__68336));
    InMux I__16626 (
            .O(N__68349),
            .I(N__68333));
    InMux I__16625 (
            .O(N__68348),
            .I(N__68330));
    Span12Mux_h I__16624 (
            .O(N__68345),
            .I(N__68327));
    Span4Mux_h I__16623 (
            .O(N__68342),
            .I(N__68324));
    LocalMux I__16622 (
            .O(N__68339),
            .I(N__68317));
    Span4Mux_h I__16621 (
            .O(N__68336),
            .I(N__68317));
    LocalMux I__16620 (
            .O(N__68333),
            .I(N__68317));
    LocalMux I__16619 (
            .O(N__68330),
            .I(\c0.data_in_frame_17_2 ));
    Odrv12 I__16618 (
            .O(N__68327),
            .I(\c0.data_in_frame_17_2 ));
    Odrv4 I__16617 (
            .O(N__68324),
            .I(\c0.data_in_frame_17_2 ));
    Odrv4 I__16616 (
            .O(N__68317),
            .I(\c0.data_in_frame_17_2 ));
    InMux I__16615 (
            .O(N__68308),
            .I(N__68304));
    InMux I__16614 (
            .O(N__68307),
            .I(N__68301));
    LocalMux I__16613 (
            .O(N__68304),
            .I(N__68296));
    LocalMux I__16612 (
            .O(N__68301),
            .I(N__68293));
    InMux I__16611 (
            .O(N__68300),
            .I(N__68290));
    InMux I__16610 (
            .O(N__68299),
            .I(N__68286));
    Span4Mux_h I__16609 (
            .O(N__68296),
            .I(N__68283));
    Span4Mux_h I__16608 (
            .O(N__68293),
            .I(N__68278));
    LocalMux I__16607 (
            .O(N__68290),
            .I(N__68278));
    InMux I__16606 (
            .O(N__68289),
            .I(N__68275));
    LocalMux I__16605 (
            .O(N__68286),
            .I(N__68271));
    Span4Mux_h I__16604 (
            .O(N__68283),
            .I(N__68266));
    Span4Mux_h I__16603 (
            .O(N__68278),
            .I(N__68266));
    LocalMux I__16602 (
            .O(N__68275),
            .I(N__68263));
    InMux I__16601 (
            .O(N__68274),
            .I(N__68260));
    Span4Mux_v I__16600 (
            .O(N__68271),
            .I(N__68257));
    Span4Mux_v I__16599 (
            .O(N__68266),
            .I(N__68252));
    Span4Mux_h I__16598 (
            .O(N__68263),
            .I(N__68252));
    LocalMux I__16597 (
            .O(N__68260),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__16596 (
            .O(N__68257),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__16595 (
            .O(N__68252),
            .I(\c0.data_in_frame_17_3 ));
    InMux I__16594 (
            .O(N__68245),
            .I(N__68242));
    LocalMux I__16593 (
            .O(N__68242),
            .I(N__68239));
    Odrv4 I__16592 (
            .O(N__68239),
            .I(\c0.n14_adj_3436 ));
    InMux I__16591 (
            .O(N__68236),
            .I(N__68229));
    InMux I__16590 (
            .O(N__68235),
            .I(N__68229));
    InMux I__16589 (
            .O(N__68234),
            .I(N__68224));
    LocalMux I__16588 (
            .O(N__68229),
            .I(N__68221));
    CascadeMux I__16587 (
            .O(N__68228),
            .I(N__68218));
    InMux I__16586 (
            .O(N__68227),
            .I(N__68214));
    LocalMux I__16585 (
            .O(N__68224),
            .I(N__68208));
    Span4Mux_h I__16584 (
            .O(N__68221),
            .I(N__68208));
    InMux I__16583 (
            .O(N__68218),
            .I(N__68203));
    InMux I__16582 (
            .O(N__68217),
            .I(N__68203));
    LocalMux I__16581 (
            .O(N__68214),
            .I(N__68200));
    InMux I__16580 (
            .O(N__68213),
            .I(N__68197));
    Span4Mux_v I__16579 (
            .O(N__68208),
            .I(N__68192));
    LocalMux I__16578 (
            .O(N__68203),
            .I(N__68185));
    Span4Mux_h I__16577 (
            .O(N__68200),
            .I(N__68185));
    LocalMux I__16576 (
            .O(N__68197),
            .I(N__68185));
    InMux I__16575 (
            .O(N__68196),
            .I(N__68180));
    InMux I__16574 (
            .O(N__68195),
            .I(N__68180));
    Odrv4 I__16573 (
            .O(N__68192),
            .I(\c0.data_in_frame_20_4 ));
    Odrv4 I__16572 (
            .O(N__68185),
            .I(\c0.data_in_frame_20_4 ));
    LocalMux I__16571 (
            .O(N__68180),
            .I(\c0.data_in_frame_20_4 ));
    CascadeMux I__16570 (
            .O(N__68173),
            .I(N__68170));
    InMux I__16569 (
            .O(N__68170),
            .I(N__68166));
    InMux I__16568 (
            .O(N__68169),
            .I(N__68162));
    LocalMux I__16567 (
            .O(N__68166),
            .I(N__68159));
    InMux I__16566 (
            .O(N__68165),
            .I(N__68154));
    LocalMux I__16565 (
            .O(N__68162),
            .I(N__68151));
    Span4Mux_v I__16564 (
            .O(N__68159),
            .I(N__68148));
    InMux I__16563 (
            .O(N__68158),
            .I(N__68143));
    InMux I__16562 (
            .O(N__68157),
            .I(N__68143));
    LocalMux I__16561 (
            .O(N__68154),
            .I(N__68140));
    Span4Mux_v I__16560 (
            .O(N__68151),
            .I(N__68133));
    Span4Mux_h I__16559 (
            .O(N__68148),
            .I(N__68133));
    LocalMux I__16558 (
            .O(N__68143),
            .I(N__68133));
    Span12Mux_v I__16557 (
            .O(N__68140),
            .I(N__68130));
    Odrv4 I__16556 (
            .O(N__68133),
            .I(\c0.n19274 ));
    Odrv12 I__16555 (
            .O(N__68130),
            .I(\c0.n19274 ));
    CascadeMux I__16554 (
            .O(N__68125),
            .I(N__68121));
    InMux I__16553 (
            .O(N__68124),
            .I(N__68114));
    InMux I__16552 (
            .O(N__68121),
            .I(N__68114));
    InMux I__16551 (
            .O(N__68120),
            .I(N__68109));
    InMux I__16550 (
            .O(N__68119),
            .I(N__68106));
    LocalMux I__16549 (
            .O(N__68114),
            .I(N__68101));
    InMux I__16548 (
            .O(N__68113),
            .I(N__68096));
    InMux I__16547 (
            .O(N__68112),
            .I(N__68096));
    LocalMux I__16546 (
            .O(N__68109),
            .I(N__68093));
    LocalMux I__16545 (
            .O(N__68106),
            .I(N__68090));
    InMux I__16544 (
            .O(N__68105),
            .I(N__68085));
    InMux I__16543 (
            .O(N__68104),
            .I(N__68085));
    Span4Mux_h I__16542 (
            .O(N__68101),
            .I(N__68081));
    LocalMux I__16541 (
            .O(N__68096),
            .I(N__68076));
    Span4Mux_v I__16540 (
            .O(N__68093),
            .I(N__68076));
    Span4Mux_h I__16539 (
            .O(N__68090),
            .I(N__68071));
    LocalMux I__16538 (
            .O(N__68085),
            .I(N__68071));
    InMux I__16537 (
            .O(N__68084),
            .I(N__68067));
    Span4Mux_v I__16536 (
            .O(N__68081),
            .I(N__68064));
    Span4Mux_h I__16535 (
            .O(N__68076),
            .I(N__68059));
    Span4Mux_v I__16534 (
            .O(N__68071),
            .I(N__68059));
    InMux I__16533 (
            .O(N__68070),
            .I(N__68056));
    LocalMux I__16532 (
            .O(N__68067),
            .I(\c0.data_in_frame_20_3 ));
    Odrv4 I__16531 (
            .O(N__68064),
            .I(\c0.data_in_frame_20_3 ));
    Odrv4 I__16530 (
            .O(N__68059),
            .I(\c0.data_in_frame_20_3 ));
    LocalMux I__16529 (
            .O(N__68056),
            .I(\c0.data_in_frame_20_3 ));
    CascadeMux I__16528 (
            .O(N__68047),
            .I(N__68044));
    InMux I__16527 (
            .O(N__68044),
            .I(N__68040));
    InMux I__16526 (
            .O(N__68043),
            .I(N__68037));
    LocalMux I__16525 (
            .O(N__68040),
            .I(N__68034));
    LocalMux I__16524 (
            .O(N__68037),
            .I(N__68031));
    Span4Mux_h I__16523 (
            .O(N__68034),
            .I(N__68026));
    Span4Mux_v I__16522 (
            .O(N__68031),
            .I(N__68026));
    Odrv4 I__16521 (
            .O(N__68026),
            .I(\c0.n54_adj_3388 ));
    InMux I__16520 (
            .O(N__68023),
            .I(N__68019));
    InMux I__16519 (
            .O(N__68022),
            .I(N__68014));
    LocalMux I__16518 (
            .O(N__68019),
            .I(N__68011));
    InMux I__16517 (
            .O(N__68018),
            .I(N__68008));
    InMux I__16516 (
            .O(N__68017),
            .I(N__68005));
    LocalMux I__16515 (
            .O(N__68014),
            .I(N__68002));
    Odrv12 I__16514 (
            .O(N__68011),
            .I(\c0.n32_adj_3310 ));
    LocalMux I__16513 (
            .O(N__68008),
            .I(\c0.n32_adj_3310 ));
    LocalMux I__16512 (
            .O(N__68005),
            .I(\c0.n32_adj_3310 ));
    Odrv4 I__16511 (
            .O(N__68002),
            .I(\c0.n32_adj_3310 ));
    InMux I__16510 (
            .O(N__67993),
            .I(N__67990));
    LocalMux I__16509 (
            .O(N__67990),
            .I(\c0.n43_adj_3131 ));
    InMux I__16508 (
            .O(N__67987),
            .I(N__67984));
    LocalMux I__16507 (
            .O(N__67984),
            .I(N__67976));
    InMux I__16506 (
            .O(N__67983),
            .I(N__67973));
    InMux I__16505 (
            .O(N__67982),
            .I(N__67968));
    InMux I__16504 (
            .O(N__67981),
            .I(N__67965));
    InMux I__16503 (
            .O(N__67980),
            .I(N__67961));
    InMux I__16502 (
            .O(N__67979),
            .I(N__67958));
    Span4Mux_h I__16501 (
            .O(N__67976),
            .I(N__67953));
    LocalMux I__16500 (
            .O(N__67973),
            .I(N__67953));
    InMux I__16499 (
            .O(N__67972),
            .I(N__67941));
    InMux I__16498 (
            .O(N__67971),
            .I(N__67936));
    LocalMux I__16497 (
            .O(N__67968),
            .I(N__67933));
    LocalMux I__16496 (
            .O(N__67965),
            .I(N__67929));
    InMux I__16495 (
            .O(N__67964),
            .I(N__67926));
    LocalMux I__16494 (
            .O(N__67961),
            .I(N__67923));
    LocalMux I__16493 (
            .O(N__67958),
            .I(N__67916));
    Span4Mux_v I__16492 (
            .O(N__67953),
            .I(N__67913));
    InMux I__16491 (
            .O(N__67952),
            .I(N__67908));
    InMux I__16490 (
            .O(N__67951),
            .I(N__67905));
    InMux I__16489 (
            .O(N__67950),
            .I(N__67900));
    InMux I__16488 (
            .O(N__67949),
            .I(N__67900));
    InMux I__16487 (
            .O(N__67948),
            .I(N__67897));
    InMux I__16486 (
            .O(N__67947),
            .I(N__67890));
    InMux I__16485 (
            .O(N__67946),
            .I(N__67890));
    InMux I__16484 (
            .O(N__67945),
            .I(N__67890));
    CascadeMux I__16483 (
            .O(N__67944),
            .I(N__67886));
    LocalMux I__16482 (
            .O(N__67941),
            .I(N__67883));
    InMux I__16481 (
            .O(N__67940),
            .I(N__67880));
    InMux I__16480 (
            .O(N__67939),
            .I(N__67877));
    LocalMux I__16479 (
            .O(N__67936),
            .I(N__67872));
    Span4Mux_h I__16478 (
            .O(N__67933),
            .I(N__67872));
    InMux I__16477 (
            .O(N__67932),
            .I(N__67869));
    Span4Mux_h I__16476 (
            .O(N__67929),
            .I(N__67866));
    LocalMux I__16475 (
            .O(N__67926),
            .I(N__67861));
    Span4Mux_h I__16474 (
            .O(N__67923),
            .I(N__67861));
    InMux I__16473 (
            .O(N__67922),
            .I(N__67858));
    InMux I__16472 (
            .O(N__67921),
            .I(N__67855));
    InMux I__16471 (
            .O(N__67920),
            .I(N__67849));
    InMux I__16470 (
            .O(N__67919),
            .I(N__67849));
    Span4Mux_h I__16469 (
            .O(N__67916),
            .I(N__67846));
    Span4Mux_v I__16468 (
            .O(N__67913),
            .I(N__67843));
    InMux I__16467 (
            .O(N__67912),
            .I(N__67840));
    InMux I__16466 (
            .O(N__67911),
            .I(N__67837));
    LocalMux I__16465 (
            .O(N__67908),
            .I(N__67826));
    LocalMux I__16464 (
            .O(N__67905),
            .I(N__67826));
    LocalMux I__16463 (
            .O(N__67900),
            .I(N__67826));
    LocalMux I__16462 (
            .O(N__67897),
            .I(N__67826));
    LocalMux I__16461 (
            .O(N__67890),
            .I(N__67826));
    InMux I__16460 (
            .O(N__67889),
            .I(N__67821));
    InMux I__16459 (
            .O(N__67886),
            .I(N__67821));
    Span4Mux_v I__16458 (
            .O(N__67883),
            .I(N__67818));
    LocalMux I__16457 (
            .O(N__67880),
            .I(N__67813));
    LocalMux I__16456 (
            .O(N__67877),
            .I(N__67813));
    Span4Mux_h I__16455 (
            .O(N__67872),
            .I(N__67808));
    LocalMux I__16454 (
            .O(N__67869),
            .I(N__67808));
    Span4Mux_h I__16453 (
            .O(N__67866),
            .I(N__67803));
    Span4Mux_v I__16452 (
            .O(N__67861),
            .I(N__67803));
    LocalMux I__16451 (
            .O(N__67858),
            .I(N__67799));
    LocalMux I__16450 (
            .O(N__67855),
            .I(N__67796));
    InMux I__16449 (
            .O(N__67854),
            .I(N__67793));
    LocalMux I__16448 (
            .O(N__67849),
            .I(N__67790));
    Span4Mux_h I__16447 (
            .O(N__67846),
            .I(N__67785));
    Span4Mux_v I__16446 (
            .O(N__67843),
            .I(N__67785));
    LocalMux I__16445 (
            .O(N__67840),
            .I(N__67778));
    LocalMux I__16444 (
            .O(N__67837),
            .I(N__67778));
    Span4Mux_v I__16443 (
            .O(N__67826),
            .I(N__67778));
    LocalMux I__16442 (
            .O(N__67821),
            .I(N__67773));
    Sp12to4 I__16441 (
            .O(N__67818),
            .I(N__67770));
    Span12Mux_h I__16440 (
            .O(N__67813),
            .I(N__67763));
    Sp12to4 I__16439 (
            .O(N__67808),
            .I(N__67763));
    Sp12to4 I__16438 (
            .O(N__67803),
            .I(N__67763));
    InMux I__16437 (
            .O(N__67802),
            .I(N__67760));
    Span4Mux_v I__16436 (
            .O(N__67799),
            .I(N__67757));
    Span4Mux_h I__16435 (
            .O(N__67796),
            .I(N__67750));
    LocalMux I__16434 (
            .O(N__67793),
            .I(N__67750));
    Span4Mux_h I__16433 (
            .O(N__67790),
            .I(N__67750));
    Span4Mux_h I__16432 (
            .O(N__67785),
            .I(N__67747));
    Span4Mux_v I__16431 (
            .O(N__67778),
            .I(N__67744));
    InMux I__16430 (
            .O(N__67777),
            .I(N__67741));
    InMux I__16429 (
            .O(N__67776),
            .I(N__67738));
    Span12Mux_h I__16428 (
            .O(N__67773),
            .I(N__67733));
    Span12Mux_v I__16427 (
            .O(N__67770),
            .I(N__67733));
    Span12Mux_v I__16426 (
            .O(N__67763),
            .I(N__67730));
    LocalMux I__16425 (
            .O(N__67760),
            .I(N__67723));
    Span4Mux_h I__16424 (
            .O(N__67757),
            .I(N__67723));
    Span4Mux_v I__16423 (
            .O(N__67750),
            .I(N__67723));
    Span4Mux_v I__16422 (
            .O(N__67747),
            .I(N__67718));
    Span4Mux_h I__16421 (
            .O(N__67744),
            .I(N__67718));
    LocalMux I__16420 (
            .O(N__67741),
            .I(rx_data_5));
    LocalMux I__16419 (
            .O(N__67738),
            .I(rx_data_5));
    Odrv12 I__16418 (
            .O(N__67733),
            .I(rx_data_5));
    Odrv12 I__16417 (
            .O(N__67730),
            .I(rx_data_5));
    Odrv4 I__16416 (
            .O(N__67723),
            .I(rx_data_5));
    Odrv4 I__16415 (
            .O(N__67718),
            .I(rx_data_5));
    CascadeMux I__16414 (
            .O(N__67705),
            .I(N__67701));
    CascadeMux I__16413 (
            .O(N__67704),
            .I(N__67698));
    InMux I__16412 (
            .O(N__67701),
            .I(N__67693));
    InMux I__16411 (
            .O(N__67698),
            .I(N__67690));
    InMux I__16410 (
            .O(N__67697),
            .I(N__67685));
    InMux I__16409 (
            .O(N__67696),
            .I(N__67685));
    LocalMux I__16408 (
            .O(N__67693),
            .I(N__67682));
    LocalMux I__16407 (
            .O(N__67690),
            .I(\c0.data_in_frame_20_2 ));
    LocalMux I__16406 (
            .O(N__67685),
            .I(\c0.data_in_frame_20_2 ));
    Odrv4 I__16405 (
            .O(N__67682),
            .I(\c0.data_in_frame_20_2 ));
    InMux I__16404 (
            .O(N__67675),
            .I(N__67670));
    InMux I__16403 (
            .O(N__67674),
            .I(N__67667));
    InMux I__16402 (
            .O(N__67673),
            .I(N__67663));
    LocalMux I__16401 (
            .O(N__67670),
            .I(N__67658));
    LocalMux I__16400 (
            .O(N__67667),
            .I(N__67658));
    InMux I__16399 (
            .O(N__67666),
            .I(N__67654));
    LocalMux I__16398 (
            .O(N__67663),
            .I(N__67649));
    Span4Mux_v I__16397 (
            .O(N__67658),
            .I(N__67649));
    InMux I__16396 (
            .O(N__67657),
            .I(N__67646));
    LocalMux I__16395 (
            .O(N__67654),
            .I(\c0.n20840 ));
    Odrv4 I__16394 (
            .O(N__67649),
            .I(\c0.n20840 ));
    LocalMux I__16393 (
            .O(N__67646),
            .I(\c0.n20840 ));
    InMux I__16392 (
            .O(N__67639),
            .I(N__67636));
    LocalMux I__16391 (
            .O(N__67636),
            .I(N__67633));
    Span4Mux_v I__16390 (
            .O(N__67633),
            .I(N__67630));
    Span4Mux_h I__16389 (
            .O(N__67630),
            .I(N__67626));
    InMux I__16388 (
            .O(N__67629),
            .I(N__67623));
    Odrv4 I__16387 (
            .O(N__67626),
            .I(\c0.n22_adj_3322 ));
    LocalMux I__16386 (
            .O(N__67623),
            .I(\c0.n22_adj_3322 ));
    InMux I__16385 (
            .O(N__67618),
            .I(N__67615));
    LocalMux I__16384 (
            .O(N__67615),
            .I(N__67610));
    InMux I__16383 (
            .O(N__67614),
            .I(N__67607));
    InMux I__16382 (
            .O(N__67613),
            .I(N__67604));
    Span4Mux_h I__16381 (
            .O(N__67610),
            .I(N__67601));
    LocalMux I__16380 (
            .O(N__67607),
            .I(N__67598));
    LocalMux I__16379 (
            .O(N__67604),
            .I(N__67595));
    Span4Mux_v I__16378 (
            .O(N__67601),
            .I(N__67590));
    Span4Mux_v I__16377 (
            .O(N__67598),
            .I(N__67590));
    Span4Mux_h I__16376 (
            .O(N__67595),
            .I(N__67587));
    Odrv4 I__16375 (
            .O(N__67590),
            .I(\c0.n11971 ));
    Odrv4 I__16374 (
            .O(N__67587),
            .I(\c0.n11971 ));
    InMux I__16373 (
            .O(N__67582),
            .I(N__67579));
    LocalMux I__16372 (
            .O(N__67579),
            .I(\c0.n19484 ));
    CascadeMux I__16371 (
            .O(N__67576),
            .I(\c0.n7_adj_3072_cascade_ ));
    CascadeMux I__16370 (
            .O(N__67573),
            .I(\c0.n18413_cascade_ ));
    InMux I__16369 (
            .O(N__67570),
            .I(N__67567));
    LocalMux I__16368 (
            .O(N__67567),
            .I(N__67563));
    InMux I__16367 (
            .O(N__67566),
            .I(N__67559));
    Span4Mux_v I__16366 (
            .O(N__67563),
            .I(N__67556));
    CascadeMux I__16365 (
            .O(N__67562),
            .I(N__67553));
    LocalMux I__16364 (
            .O(N__67559),
            .I(N__67550));
    Span4Mux_h I__16363 (
            .O(N__67556),
            .I(N__67547));
    InMux I__16362 (
            .O(N__67553),
            .I(N__67544));
    Span4Mux_h I__16361 (
            .O(N__67550),
            .I(N__67541));
    Span4Mux_h I__16360 (
            .O(N__67547),
            .I(N__67538));
    LocalMux I__16359 (
            .O(N__67544),
            .I(\c0.data_in_frame_26_3 ));
    Odrv4 I__16358 (
            .O(N__67541),
            .I(\c0.data_in_frame_26_3 ));
    Odrv4 I__16357 (
            .O(N__67538),
            .I(\c0.data_in_frame_26_3 ));
    InMux I__16356 (
            .O(N__67531),
            .I(N__67523));
    InMux I__16355 (
            .O(N__67530),
            .I(N__67519));
    InMux I__16354 (
            .O(N__67529),
            .I(N__67516));
    InMux I__16353 (
            .O(N__67528),
            .I(N__67511));
    InMux I__16352 (
            .O(N__67527),
            .I(N__67511));
    InMux I__16351 (
            .O(N__67526),
            .I(N__67508));
    LocalMux I__16350 (
            .O(N__67523),
            .I(N__67505));
    InMux I__16349 (
            .O(N__67522),
            .I(N__67501));
    LocalMux I__16348 (
            .O(N__67519),
            .I(N__67498));
    LocalMux I__16347 (
            .O(N__67516),
            .I(N__67495));
    LocalMux I__16346 (
            .O(N__67511),
            .I(N__67492));
    LocalMux I__16345 (
            .O(N__67508),
            .I(N__67489));
    Span4Mux_h I__16344 (
            .O(N__67505),
            .I(N__67486));
    InMux I__16343 (
            .O(N__67504),
            .I(N__67483));
    LocalMux I__16342 (
            .O(N__67501),
            .I(N__67478));
    Span4Mux_v I__16341 (
            .O(N__67498),
            .I(N__67478));
    Span4Mux_v I__16340 (
            .O(N__67495),
            .I(N__67475));
    Span4Mux_h I__16339 (
            .O(N__67492),
            .I(N__67472));
    Span4Mux_h I__16338 (
            .O(N__67489),
            .I(N__67467));
    Span4Mux_h I__16337 (
            .O(N__67486),
            .I(N__67467));
    LocalMux I__16336 (
            .O(N__67483),
            .I(N__67462));
    Span4Mux_v I__16335 (
            .O(N__67478),
            .I(N__67462));
    Span4Mux_h I__16334 (
            .O(N__67475),
            .I(N__67459));
    Span4Mux_h I__16333 (
            .O(N__67472),
            .I(N__67456));
    Span4Mux_v I__16332 (
            .O(N__67467),
            .I(N__67453));
    Span4Mux_h I__16331 (
            .O(N__67462),
            .I(N__67450));
    Sp12to4 I__16330 (
            .O(N__67459),
            .I(N__67447));
    Odrv4 I__16329 (
            .O(N__67456),
            .I(n19127));
    Odrv4 I__16328 (
            .O(N__67453),
            .I(n19127));
    Odrv4 I__16327 (
            .O(N__67450),
            .I(n19127));
    Odrv12 I__16326 (
            .O(N__67447),
            .I(n19127));
    InMux I__16325 (
            .O(N__67438),
            .I(N__67435));
    LocalMux I__16324 (
            .O(N__67435),
            .I(N__67431));
    CascadeMux I__16323 (
            .O(N__67434),
            .I(N__67428));
    Span4Mux_v I__16322 (
            .O(N__67431),
            .I(N__67424));
    InMux I__16321 (
            .O(N__67428),
            .I(N__67421));
    InMux I__16320 (
            .O(N__67427),
            .I(N__67418));
    Sp12to4 I__16319 (
            .O(N__67424),
            .I(N__67413));
    LocalMux I__16318 (
            .O(N__67421),
            .I(N__67413));
    LocalMux I__16317 (
            .O(N__67418),
            .I(data_in_frame_22_5));
    Odrv12 I__16316 (
            .O(N__67413),
            .I(data_in_frame_22_5));
    InMux I__16315 (
            .O(N__67408),
            .I(N__67405));
    LocalMux I__16314 (
            .O(N__67405),
            .I(N__67401));
    InMux I__16313 (
            .O(N__67404),
            .I(N__67398));
    Span4Mux_v I__16312 (
            .O(N__67401),
            .I(N__67393));
    LocalMux I__16311 (
            .O(N__67398),
            .I(N__67393));
    Span4Mux_h I__16310 (
            .O(N__67393),
            .I(N__67390));
    Odrv4 I__16309 (
            .O(N__67390),
            .I(\c0.n9_adj_3069 ));
    InMux I__16308 (
            .O(N__67387),
            .I(N__67383));
    InMux I__16307 (
            .O(N__67386),
            .I(N__67380));
    LocalMux I__16306 (
            .O(N__67383),
            .I(N__67373));
    LocalMux I__16305 (
            .O(N__67380),
            .I(N__67373));
    InMux I__16304 (
            .O(N__67379),
            .I(N__67368));
    InMux I__16303 (
            .O(N__67378),
            .I(N__67368));
    Span4Mux_v I__16302 (
            .O(N__67373),
            .I(N__67365));
    LocalMux I__16301 (
            .O(N__67368),
            .I(\c0.n20451 ));
    Odrv4 I__16300 (
            .O(N__67365),
            .I(\c0.n20451 ));
    InMux I__16299 (
            .O(N__67360),
            .I(N__67357));
    LocalMux I__16298 (
            .O(N__67357),
            .I(\c0.n8_adj_3070 ));
    InMux I__16297 (
            .O(N__67354),
            .I(N__67351));
    LocalMux I__16296 (
            .O(N__67351),
            .I(\c0.n19315 ));
    InMux I__16295 (
            .O(N__67348),
            .I(N__67345));
    LocalMux I__16294 (
            .O(N__67345),
            .I(N__67342));
    Span4Mux_v I__16293 (
            .O(N__67342),
            .I(N__67339));
    Span4Mux_h I__16292 (
            .O(N__67339),
            .I(N__67336));
    Span4Mux_v I__16291 (
            .O(N__67336),
            .I(N__67333));
    Odrv4 I__16290 (
            .O(N__67333),
            .I(\c0.n26_adj_3550 ));
    InMux I__16289 (
            .O(N__67330),
            .I(N__67327));
    LocalMux I__16288 (
            .O(N__67327),
            .I(N__67324));
    Span4Mux_h I__16287 (
            .O(N__67324),
            .I(N__67321));
    Span4Mux_v I__16286 (
            .O(N__67321),
            .I(N__67318));
    Odrv4 I__16285 (
            .O(N__67318),
            .I(\c0.n27_adj_3551 ));
    CascadeMux I__16284 (
            .O(N__67315),
            .I(N__67312));
    InMux I__16283 (
            .O(N__67312),
            .I(N__67309));
    LocalMux I__16282 (
            .O(N__67309),
            .I(N__67306));
    Odrv12 I__16281 (
            .O(N__67306),
            .I(\c0.n25_adj_3553 ));
    InMux I__16280 (
            .O(N__67303),
            .I(N__67299));
    InMux I__16279 (
            .O(N__67302),
            .I(N__67296));
    LocalMux I__16278 (
            .O(N__67299),
            .I(N__67293));
    LocalMux I__16277 (
            .O(N__67296),
            .I(N__67290));
    Span4Mux_h I__16276 (
            .O(N__67293),
            .I(N__67285));
    Span4Mux_h I__16275 (
            .O(N__67290),
            .I(N__67282));
    InMux I__16274 (
            .O(N__67289),
            .I(N__67277));
    InMux I__16273 (
            .O(N__67288),
            .I(N__67277));
    Odrv4 I__16272 (
            .O(N__67285),
            .I(\c0.n49_adj_3358 ));
    Odrv4 I__16271 (
            .O(N__67282),
            .I(\c0.n49_adj_3358 ));
    LocalMux I__16270 (
            .O(N__67277),
            .I(\c0.n49_adj_3358 ));
    CascadeMux I__16269 (
            .O(N__67270),
            .I(N__67267));
    InMux I__16268 (
            .O(N__67267),
            .I(N__67260));
    InMux I__16267 (
            .O(N__67266),
            .I(N__67255));
    InMux I__16266 (
            .O(N__67265),
            .I(N__67255));
    InMux I__16265 (
            .O(N__67264),
            .I(N__67250));
    InMux I__16264 (
            .O(N__67263),
            .I(N__67250));
    LocalMux I__16263 (
            .O(N__67260),
            .I(\c0.n17832 ));
    LocalMux I__16262 (
            .O(N__67255),
            .I(\c0.n17832 ));
    LocalMux I__16261 (
            .O(N__67250),
            .I(\c0.n17832 ));
    InMux I__16260 (
            .O(N__67243),
            .I(N__67234));
    InMux I__16259 (
            .O(N__67242),
            .I(N__67234));
    InMux I__16258 (
            .O(N__67241),
            .I(N__67234));
    LocalMux I__16257 (
            .O(N__67234),
            .I(\c0.n40_adj_3271 ));
    CascadeMux I__16256 (
            .O(N__67231),
            .I(N__67228));
    InMux I__16255 (
            .O(N__67228),
            .I(N__67213));
    InMux I__16254 (
            .O(N__67227),
            .I(N__67213));
    InMux I__16253 (
            .O(N__67226),
            .I(N__67204));
    InMux I__16252 (
            .O(N__67225),
            .I(N__67204));
    InMux I__16251 (
            .O(N__67224),
            .I(N__67204));
    InMux I__16250 (
            .O(N__67223),
            .I(N__67204));
    CascadeMux I__16249 (
            .O(N__67222),
            .I(N__67201));
    InMux I__16248 (
            .O(N__67221),
            .I(N__67191));
    InMux I__16247 (
            .O(N__67220),
            .I(N__67191));
    CascadeMux I__16246 (
            .O(N__67219),
            .I(N__67188));
    InMux I__16245 (
            .O(N__67218),
            .I(N__67184));
    LocalMux I__16244 (
            .O(N__67213),
            .I(N__67179));
    LocalMux I__16243 (
            .O(N__67204),
            .I(N__67179));
    InMux I__16242 (
            .O(N__67201),
            .I(N__67173));
    InMux I__16241 (
            .O(N__67200),
            .I(N__67173));
    InMux I__16240 (
            .O(N__67199),
            .I(N__67170));
    InMux I__16239 (
            .O(N__67198),
            .I(N__67167));
    InMux I__16238 (
            .O(N__67197),
            .I(N__67163));
    InMux I__16237 (
            .O(N__67196),
            .I(N__67160));
    LocalMux I__16236 (
            .O(N__67191),
            .I(N__67157));
    InMux I__16235 (
            .O(N__67188),
            .I(N__67154));
    InMux I__16234 (
            .O(N__67187),
            .I(N__67151));
    LocalMux I__16233 (
            .O(N__67184),
            .I(N__67148));
    Span4Mux_v I__16232 (
            .O(N__67179),
            .I(N__67145));
    InMux I__16231 (
            .O(N__67178),
            .I(N__67141));
    LocalMux I__16230 (
            .O(N__67173),
            .I(N__67138));
    LocalMux I__16229 (
            .O(N__67170),
            .I(N__67135));
    LocalMux I__16228 (
            .O(N__67167),
            .I(N__67132));
    InMux I__16227 (
            .O(N__67166),
            .I(N__67127));
    LocalMux I__16226 (
            .O(N__67163),
            .I(N__67122));
    LocalMux I__16225 (
            .O(N__67160),
            .I(N__67122));
    Span4Mux_h I__16224 (
            .O(N__67157),
            .I(N__67119));
    LocalMux I__16223 (
            .O(N__67154),
            .I(N__67113));
    LocalMux I__16222 (
            .O(N__67151),
            .I(N__67113));
    Span4Mux_v I__16221 (
            .O(N__67148),
            .I(N__67108));
    Span4Mux_h I__16220 (
            .O(N__67145),
            .I(N__67108));
    InMux I__16219 (
            .O(N__67144),
            .I(N__67105));
    LocalMux I__16218 (
            .O(N__67141),
            .I(N__67102));
    Span4Mux_v I__16217 (
            .O(N__67138),
            .I(N__67095));
    Span4Mux_v I__16216 (
            .O(N__67135),
            .I(N__67095));
    Span4Mux_h I__16215 (
            .O(N__67132),
            .I(N__67095));
    InMux I__16214 (
            .O(N__67131),
            .I(N__67092));
    InMux I__16213 (
            .O(N__67130),
            .I(N__67089));
    LocalMux I__16212 (
            .O(N__67127),
            .I(N__67086));
    Span4Mux_v I__16211 (
            .O(N__67122),
            .I(N__67081));
    Span4Mux_v I__16210 (
            .O(N__67119),
            .I(N__67081));
    InMux I__16209 (
            .O(N__67118),
            .I(N__67078));
    Span4Mux_h I__16208 (
            .O(N__67113),
            .I(N__67075));
    Span4Mux_h I__16207 (
            .O(N__67108),
            .I(N__67072));
    LocalMux I__16206 (
            .O(N__67105),
            .I(N__67065));
    Span4Mux_h I__16205 (
            .O(N__67102),
            .I(N__67065));
    Span4Mux_h I__16204 (
            .O(N__67095),
            .I(N__67065));
    LocalMux I__16203 (
            .O(N__67092),
            .I(N__67062));
    LocalMux I__16202 (
            .O(N__67089),
            .I(N__67057));
    Span4Mux_v I__16201 (
            .O(N__67086),
            .I(N__67057));
    Span4Mux_h I__16200 (
            .O(N__67081),
            .I(N__67054));
    LocalMux I__16199 (
            .O(N__67078),
            .I(N__67051));
    Span4Mux_h I__16198 (
            .O(N__67075),
            .I(N__67044));
    Span4Mux_h I__16197 (
            .O(N__67072),
            .I(N__67044));
    Span4Mux_v I__16196 (
            .O(N__67065),
            .I(N__67044));
    Span4Mux_h I__16195 (
            .O(N__67062),
            .I(N__67041));
    Span4Mux_v I__16194 (
            .O(N__67057),
            .I(N__67038));
    Sp12to4 I__16193 (
            .O(N__67054),
            .I(N__67035));
    Span4Mux_v I__16192 (
            .O(N__67051),
            .I(N__67030));
    Span4Mux_v I__16191 (
            .O(N__67044),
            .I(N__67030));
    Odrv4 I__16190 (
            .O(N__67041),
            .I(\c0.n19111 ));
    Odrv4 I__16189 (
            .O(N__67038),
            .I(\c0.n19111 ));
    Odrv12 I__16188 (
            .O(N__67035),
            .I(\c0.n19111 ));
    Odrv4 I__16187 (
            .O(N__67030),
            .I(\c0.n19111 ));
    CascadeMux I__16186 (
            .O(N__67021),
            .I(N__67017));
    CascadeMux I__16185 (
            .O(N__67020),
            .I(N__67014));
    InMux I__16184 (
            .O(N__67017),
            .I(N__67011));
    InMux I__16183 (
            .O(N__67014),
            .I(N__67008));
    LocalMux I__16182 (
            .O(N__67011),
            .I(N__67005));
    LocalMux I__16181 (
            .O(N__67008),
            .I(N__67002));
    Span4Mux_v I__16180 (
            .O(N__67005),
            .I(N__66999));
    Span4Mux_h I__16179 (
            .O(N__67002),
            .I(N__66994));
    Span4Mux_v I__16178 (
            .O(N__66999),
            .I(N__66994));
    Span4Mux_h I__16177 (
            .O(N__66994),
            .I(N__66991));
    Odrv4 I__16176 (
            .O(N__66991),
            .I(\c0.data_in_frame_29_3 ));
    CascadeMux I__16175 (
            .O(N__66988),
            .I(N__66984));
    CascadeMux I__16174 (
            .O(N__66987),
            .I(N__66981));
    InMux I__16173 (
            .O(N__66984),
            .I(N__66963));
    InMux I__16172 (
            .O(N__66981),
            .I(N__66963));
    InMux I__16171 (
            .O(N__66980),
            .I(N__66963));
    InMux I__16170 (
            .O(N__66979),
            .I(N__66963));
    CascadeMux I__16169 (
            .O(N__66978),
            .I(N__66959));
    CascadeMux I__16168 (
            .O(N__66977),
            .I(N__66949));
    CascadeMux I__16167 (
            .O(N__66976),
            .I(N__66944));
    CascadeMux I__16166 (
            .O(N__66975),
            .I(N__66938));
    CascadeMux I__16165 (
            .O(N__66974),
            .I(N__66935));
    InMux I__16164 (
            .O(N__66973),
            .I(N__66928));
    InMux I__16163 (
            .O(N__66972),
            .I(N__66928));
    LocalMux I__16162 (
            .O(N__66963),
            .I(N__66925));
    InMux I__16161 (
            .O(N__66962),
            .I(N__66918));
    InMux I__16160 (
            .O(N__66959),
            .I(N__66918));
    CascadeMux I__16159 (
            .O(N__66958),
            .I(N__66913));
    InMux I__16158 (
            .O(N__66957),
            .I(N__66909));
    InMux I__16157 (
            .O(N__66956),
            .I(N__66900));
    InMux I__16156 (
            .O(N__66955),
            .I(N__66900));
    InMux I__16155 (
            .O(N__66954),
            .I(N__66900));
    InMux I__16154 (
            .O(N__66953),
            .I(N__66900));
    InMux I__16153 (
            .O(N__66952),
            .I(N__66889));
    InMux I__16152 (
            .O(N__66949),
            .I(N__66889));
    InMux I__16151 (
            .O(N__66948),
            .I(N__66889));
    InMux I__16150 (
            .O(N__66947),
            .I(N__66882));
    InMux I__16149 (
            .O(N__66944),
            .I(N__66882));
    InMux I__16148 (
            .O(N__66943),
            .I(N__66882));
    InMux I__16147 (
            .O(N__66942),
            .I(N__66868));
    InMux I__16146 (
            .O(N__66941),
            .I(N__66868));
    InMux I__16145 (
            .O(N__66938),
            .I(N__66868));
    InMux I__16144 (
            .O(N__66935),
            .I(N__66868));
    InMux I__16143 (
            .O(N__66934),
            .I(N__66868));
    InMux I__16142 (
            .O(N__66933),
            .I(N__66865));
    LocalMux I__16141 (
            .O(N__66928),
            .I(N__66860));
    Span4Mux_v I__16140 (
            .O(N__66925),
            .I(N__66860));
    InMux I__16139 (
            .O(N__66924),
            .I(N__66857));
    InMux I__16138 (
            .O(N__66923),
            .I(N__66854));
    LocalMux I__16137 (
            .O(N__66918),
            .I(N__66851));
    InMux I__16136 (
            .O(N__66917),
            .I(N__66846));
    InMux I__16135 (
            .O(N__66916),
            .I(N__66841));
    InMux I__16134 (
            .O(N__66913),
            .I(N__66841));
    InMux I__16133 (
            .O(N__66912),
            .I(N__66838));
    LocalMux I__16132 (
            .O(N__66909),
            .I(N__66835));
    LocalMux I__16131 (
            .O(N__66900),
            .I(N__66832));
    InMux I__16130 (
            .O(N__66899),
            .I(N__66829));
    InMux I__16129 (
            .O(N__66898),
            .I(N__66826));
    InMux I__16128 (
            .O(N__66897),
            .I(N__66821));
    InMux I__16127 (
            .O(N__66896),
            .I(N__66821));
    LocalMux I__16126 (
            .O(N__66889),
            .I(N__66816));
    LocalMux I__16125 (
            .O(N__66882),
            .I(N__66816));
    InMux I__16124 (
            .O(N__66881),
            .I(N__66809));
    InMux I__16123 (
            .O(N__66880),
            .I(N__66809));
    InMux I__16122 (
            .O(N__66879),
            .I(N__66809));
    LocalMux I__16121 (
            .O(N__66868),
            .I(N__66806));
    LocalMux I__16120 (
            .O(N__66865),
            .I(N__66799));
    Span4Mux_h I__16119 (
            .O(N__66860),
            .I(N__66799));
    LocalMux I__16118 (
            .O(N__66857),
            .I(N__66799));
    LocalMux I__16117 (
            .O(N__66854),
            .I(N__66794));
    Span4Mux_v I__16116 (
            .O(N__66851),
            .I(N__66794));
    CascadeMux I__16115 (
            .O(N__66850),
            .I(N__66791));
    InMux I__16114 (
            .O(N__66849),
            .I(N__66788));
    LocalMux I__16113 (
            .O(N__66846),
            .I(N__66785));
    LocalMux I__16112 (
            .O(N__66841),
            .I(N__66782));
    LocalMux I__16111 (
            .O(N__66838),
            .I(N__66777));
    Span4Mux_h I__16110 (
            .O(N__66835),
            .I(N__66777));
    Span4Mux_v I__16109 (
            .O(N__66832),
            .I(N__66774));
    LocalMux I__16108 (
            .O(N__66829),
            .I(N__66771));
    LocalMux I__16107 (
            .O(N__66826),
            .I(N__66768));
    LocalMux I__16106 (
            .O(N__66821),
            .I(N__66761));
    Span4Mux_v I__16105 (
            .O(N__66816),
            .I(N__66761));
    LocalMux I__16104 (
            .O(N__66809),
            .I(N__66761));
    Span4Mux_v I__16103 (
            .O(N__66806),
            .I(N__66758));
    Span4Mux_h I__16102 (
            .O(N__66799),
            .I(N__66755));
    Sp12to4 I__16101 (
            .O(N__66794),
            .I(N__66751));
    InMux I__16100 (
            .O(N__66791),
            .I(N__66748));
    LocalMux I__16099 (
            .O(N__66788),
            .I(N__66739));
    Span4Mux_v I__16098 (
            .O(N__66785),
            .I(N__66739));
    Span4Mux_h I__16097 (
            .O(N__66782),
            .I(N__66739));
    Span4Mux_h I__16096 (
            .O(N__66777),
            .I(N__66739));
    Span4Mux_h I__16095 (
            .O(N__66774),
            .I(N__66732));
    Span4Mux_v I__16094 (
            .O(N__66771),
            .I(N__66732));
    Span4Mux_h I__16093 (
            .O(N__66768),
            .I(N__66732));
    Span4Mux_v I__16092 (
            .O(N__66761),
            .I(N__66729));
    Span4Mux_h I__16091 (
            .O(N__66758),
            .I(N__66724));
    Span4Mux_v I__16090 (
            .O(N__66755),
            .I(N__66724));
    InMux I__16089 (
            .O(N__66754),
            .I(N__66721));
    Span12Mux_v I__16088 (
            .O(N__66751),
            .I(N__66718));
    LocalMux I__16087 (
            .O(N__66748),
            .I(N__66711));
    Span4Mux_v I__16086 (
            .O(N__66739),
            .I(N__66711));
    Span4Mux_h I__16085 (
            .O(N__66732),
            .I(N__66711));
    Span4Mux_h I__16084 (
            .O(N__66729),
            .I(N__66708));
    Span4Mux_v I__16083 (
            .O(N__66724),
            .I(N__66705));
    LocalMux I__16082 (
            .O(N__66721),
            .I(\c0.n12_adj_3006 ));
    Odrv12 I__16081 (
            .O(N__66718),
            .I(\c0.n12_adj_3006 ));
    Odrv4 I__16080 (
            .O(N__66711),
            .I(\c0.n12_adj_3006 ));
    Odrv4 I__16079 (
            .O(N__66708),
            .I(\c0.n12_adj_3006 ));
    Odrv4 I__16078 (
            .O(N__66705),
            .I(\c0.n12_adj_3006 ));
    CascadeMux I__16077 (
            .O(N__66694),
            .I(N__66691));
    InMux I__16076 (
            .O(N__66691),
            .I(N__66687));
    InMux I__16075 (
            .O(N__66690),
            .I(N__66684));
    LocalMux I__16074 (
            .O(N__66687),
            .I(N__66681));
    LocalMux I__16073 (
            .O(N__66684),
            .I(N__66676));
    Span12Mux_h I__16072 (
            .O(N__66681),
            .I(N__66676));
    Odrv12 I__16071 (
            .O(N__66676),
            .I(\c0.data_in_frame_29_5 ));
    InMux I__16070 (
            .O(N__66673),
            .I(N__66670));
    LocalMux I__16069 (
            .O(N__66670),
            .I(N__66667));
    Span4Mux_h I__16068 (
            .O(N__66667),
            .I(N__66664));
    Odrv4 I__16067 (
            .O(N__66664),
            .I(\c0.n15_adj_3432 ));
    InMux I__16066 (
            .O(N__66661),
            .I(N__66658));
    LocalMux I__16065 (
            .O(N__66658),
            .I(N__66655));
    Span4Mux_v I__16064 (
            .O(N__66655),
            .I(N__66652));
    Odrv4 I__16063 (
            .O(N__66652),
            .I(\c0.n20503 ));
    CascadeMux I__16062 (
            .O(N__66649),
            .I(N__66644));
    InMux I__16061 (
            .O(N__66648),
            .I(N__66641));
    InMux I__16060 (
            .O(N__66647),
            .I(N__66636));
    InMux I__16059 (
            .O(N__66644),
            .I(N__66636));
    LocalMux I__16058 (
            .O(N__66641),
            .I(N__66633));
    LocalMux I__16057 (
            .O(N__66636),
            .I(N__66628));
    Span4Mux_h I__16056 (
            .O(N__66633),
            .I(N__66625));
    InMux I__16055 (
            .O(N__66632),
            .I(N__66622));
    InMux I__16054 (
            .O(N__66631),
            .I(N__66619));
    Span12Mux_s10_v I__16053 (
            .O(N__66628),
            .I(N__66616));
    Span4Mux_h I__16052 (
            .O(N__66625),
            .I(N__66613));
    LocalMux I__16051 (
            .O(N__66622),
            .I(data_in_frame_23_1));
    LocalMux I__16050 (
            .O(N__66619),
            .I(data_in_frame_23_1));
    Odrv12 I__16049 (
            .O(N__66616),
            .I(data_in_frame_23_1));
    Odrv4 I__16048 (
            .O(N__66613),
            .I(data_in_frame_23_1));
    CascadeMux I__16047 (
            .O(N__66604),
            .I(\c0.n20503_cascade_ ));
    InMux I__16046 (
            .O(N__66601),
            .I(N__66598));
    LocalMux I__16045 (
            .O(N__66598),
            .I(N__66595));
    Span12Mux_h I__16044 (
            .O(N__66595),
            .I(N__66592));
    Odrv12 I__16043 (
            .O(N__66592),
            .I(\c0.n12_adj_3494 ));
    InMux I__16042 (
            .O(N__66589),
            .I(N__66586));
    LocalMux I__16041 (
            .O(N__66586),
            .I(N__66583));
    Span4Mux_v I__16040 (
            .O(N__66583),
            .I(N__66579));
    InMux I__16039 (
            .O(N__66582),
            .I(N__66576));
    Odrv4 I__16038 (
            .O(N__66579),
            .I(\c0.n27_adj_3399 ));
    LocalMux I__16037 (
            .O(N__66576),
            .I(\c0.n27_adj_3399 ));
    InMux I__16036 (
            .O(N__66571),
            .I(N__66567));
    InMux I__16035 (
            .O(N__66570),
            .I(N__66564));
    LocalMux I__16034 (
            .O(N__66567),
            .I(\c0.data_in_frame_28_3 ));
    LocalMux I__16033 (
            .O(N__66564),
            .I(\c0.data_in_frame_28_3 ));
    CascadeMux I__16032 (
            .O(N__66559),
            .I(\c0.n27_adj_3399_cascade_ ));
    InMux I__16031 (
            .O(N__66556),
            .I(N__66553));
    LocalMux I__16030 (
            .O(N__66553),
            .I(N__66550));
    Span4Mux_h I__16029 (
            .O(N__66550),
            .I(N__66547));
    Span4Mux_v I__16028 (
            .O(N__66547),
            .I(N__66542));
    InMux I__16027 (
            .O(N__66546),
            .I(N__66537));
    InMux I__16026 (
            .O(N__66545),
            .I(N__66537));
    Odrv4 I__16025 (
            .O(N__66542),
            .I(\c0.data_in_frame_26_1 ));
    LocalMux I__16024 (
            .O(N__66537),
            .I(\c0.data_in_frame_26_1 ));
    CascadeMux I__16023 (
            .O(N__66532),
            .I(N__66529));
    InMux I__16022 (
            .O(N__66529),
            .I(N__66526));
    LocalMux I__16021 (
            .O(N__66526),
            .I(N__66523));
    Span4Mux_h I__16020 (
            .O(N__66523),
            .I(N__66520));
    Span4Mux_h I__16019 (
            .O(N__66520),
            .I(N__66517));
    Odrv4 I__16018 (
            .O(N__66517),
            .I(\c0.n78_adj_3414 ));
    CascadeMux I__16017 (
            .O(N__66514),
            .I(N__66511));
    InMux I__16016 (
            .O(N__66511),
            .I(N__66507));
    InMux I__16015 (
            .O(N__66510),
            .I(N__66504));
    LocalMux I__16014 (
            .O(N__66507),
            .I(N__66501));
    LocalMux I__16013 (
            .O(N__66504),
            .I(N__66497));
    Span4Mux_h I__16012 (
            .O(N__66501),
            .I(N__66493));
    InMux I__16011 (
            .O(N__66500),
            .I(N__66490));
    Span4Mux_h I__16010 (
            .O(N__66497),
            .I(N__66487));
    InMux I__16009 (
            .O(N__66496),
            .I(N__66484));
    Span4Mux_h I__16008 (
            .O(N__66493),
            .I(N__66481));
    LocalMux I__16007 (
            .O(N__66490),
            .I(N__66476));
    Span4Mux_h I__16006 (
            .O(N__66487),
            .I(N__66476));
    LocalMux I__16005 (
            .O(N__66484),
            .I(data_in_frame_23_6));
    Odrv4 I__16004 (
            .O(N__66481),
            .I(data_in_frame_23_6));
    Odrv4 I__16003 (
            .O(N__66476),
            .I(data_in_frame_23_6));
    InMux I__16002 (
            .O(N__66469),
            .I(N__66466));
    LocalMux I__16001 (
            .O(N__66466),
            .I(N__66461));
    InMux I__16000 (
            .O(N__66465),
            .I(N__66458));
    InMux I__15999 (
            .O(N__66464),
            .I(N__66455));
    Span4Mux_v I__15998 (
            .O(N__66461),
            .I(N__66448));
    LocalMux I__15997 (
            .O(N__66458),
            .I(N__66448));
    LocalMux I__15996 (
            .O(N__66455),
            .I(N__66445));
    InMux I__15995 (
            .O(N__66454),
            .I(N__66440));
    InMux I__15994 (
            .O(N__66453),
            .I(N__66440));
    Span4Mux_h I__15993 (
            .O(N__66448),
            .I(N__66437));
    Span12Mux_s10_h I__15992 (
            .O(N__66445),
            .I(N__66434));
    LocalMux I__15991 (
            .O(N__66440),
            .I(data_in_frame_23_5));
    Odrv4 I__15990 (
            .O(N__66437),
            .I(data_in_frame_23_5));
    Odrv12 I__15989 (
            .O(N__66434),
            .I(data_in_frame_23_5));
    InMux I__15988 (
            .O(N__66427),
            .I(N__66424));
    LocalMux I__15987 (
            .O(N__66424),
            .I(\c0.n19487 ));
    CascadeMux I__15986 (
            .O(N__66421),
            .I(N__66418));
    InMux I__15985 (
            .O(N__66418),
            .I(N__66411));
    InMux I__15984 (
            .O(N__66417),
            .I(N__66411));
    InMux I__15983 (
            .O(N__66416),
            .I(N__66408));
    LocalMux I__15982 (
            .O(N__66411),
            .I(N__66405));
    LocalMux I__15981 (
            .O(N__66408),
            .I(N__66402));
    Span4Mux_h I__15980 (
            .O(N__66405),
            .I(N__66397));
    Span4Mux_h I__15979 (
            .O(N__66402),
            .I(N__66397));
    Span4Mux_v I__15978 (
            .O(N__66397),
            .I(N__66392));
    InMux I__15977 (
            .O(N__66396),
            .I(N__66387));
    InMux I__15976 (
            .O(N__66395),
            .I(N__66387));
    Odrv4 I__15975 (
            .O(N__66392),
            .I(data_in_frame_23_7));
    LocalMux I__15974 (
            .O(N__66387),
            .I(data_in_frame_23_7));
    InMux I__15973 (
            .O(N__66382),
            .I(N__66378));
    InMux I__15972 (
            .O(N__66381),
            .I(N__66375));
    LocalMux I__15971 (
            .O(N__66378),
            .I(N__66370));
    LocalMux I__15970 (
            .O(N__66375),
            .I(N__66370));
    Span4Mux_v I__15969 (
            .O(N__66370),
            .I(N__66367));
    Span4Mux_h I__15968 (
            .O(N__66367),
            .I(N__66364));
    Odrv4 I__15967 (
            .O(N__66364),
            .I(\c0.n19251 ));
    InMux I__15966 (
            .O(N__66361),
            .I(N__66358));
    LocalMux I__15965 (
            .O(N__66358),
            .I(N__66355));
    Span4Mux_v I__15964 (
            .O(N__66355),
            .I(N__66351));
    InMux I__15963 (
            .O(N__66354),
            .I(N__66348));
    Span4Mux_v I__15962 (
            .O(N__66351),
            .I(N__66345));
    LocalMux I__15961 (
            .O(N__66348),
            .I(N__66342));
    Odrv4 I__15960 (
            .O(N__66345),
            .I(\c0.n7_adj_3347 ));
    Odrv12 I__15959 (
            .O(N__66342),
            .I(\c0.n7_adj_3347 ));
    InMux I__15958 (
            .O(N__66337),
            .I(N__66333));
    CascadeMux I__15957 (
            .O(N__66336),
            .I(N__66330));
    LocalMux I__15956 (
            .O(N__66333),
            .I(N__66327));
    InMux I__15955 (
            .O(N__66330),
            .I(N__66323));
    Span4Mux_v I__15954 (
            .O(N__66327),
            .I(N__66320));
    InMux I__15953 (
            .O(N__66326),
            .I(N__66317));
    LocalMux I__15952 (
            .O(N__66323),
            .I(\c0.data_in_frame_10_6 ));
    Odrv4 I__15951 (
            .O(N__66320),
            .I(\c0.data_in_frame_10_6 ));
    LocalMux I__15950 (
            .O(N__66317),
            .I(\c0.data_in_frame_10_6 ));
    CascadeMux I__15949 (
            .O(N__66310),
            .I(N__66307));
    InMux I__15948 (
            .O(N__66307),
            .I(N__66304));
    LocalMux I__15947 (
            .O(N__66304),
            .I(N__66301));
    Odrv4 I__15946 (
            .O(N__66301),
            .I(\c0.n19359 ));
    InMux I__15945 (
            .O(N__66298),
            .I(N__66295));
    LocalMux I__15944 (
            .O(N__66295),
            .I(N__66291));
    InMux I__15943 (
            .O(N__66294),
            .I(N__66288));
    Span4Mux_v I__15942 (
            .O(N__66291),
            .I(N__66281));
    LocalMux I__15941 (
            .O(N__66288),
            .I(N__66281));
    InMux I__15940 (
            .O(N__66287),
            .I(N__66278));
    CascadeMux I__15939 (
            .O(N__66286),
            .I(N__66275));
    Span4Mux_h I__15938 (
            .O(N__66281),
            .I(N__66272));
    LocalMux I__15937 (
            .O(N__66278),
            .I(N__66269));
    InMux I__15936 (
            .O(N__66275),
            .I(N__66266));
    Span4Mux_v I__15935 (
            .O(N__66272),
            .I(N__66261));
    Span4Mux_v I__15934 (
            .O(N__66269),
            .I(N__66261));
    LocalMux I__15933 (
            .O(N__66266),
            .I(\c0.data_in_frame_12_6 ));
    Odrv4 I__15932 (
            .O(N__66261),
            .I(\c0.data_in_frame_12_6 ));
    InMux I__15931 (
            .O(N__66256),
            .I(N__66253));
    LocalMux I__15930 (
            .O(N__66253),
            .I(N__66250));
    Span4Mux_v I__15929 (
            .O(N__66250),
            .I(N__66247));
    Odrv4 I__15928 (
            .O(N__66247),
            .I(\c0.n22_adj_3535 ));
    InMux I__15927 (
            .O(N__66244),
            .I(N__66240));
    InMux I__15926 (
            .O(N__66243),
            .I(N__66236));
    LocalMux I__15925 (
            .O(N__66240),
            .I(N__66233));
    CascadeMux I__15924 (
            .O(N__66239),
            .I(N__66230));
    LocalMux I__15923 (
            .O(N__66236),
            .I(N__66227));
    Span4Mux_h I__15922 (
            .O(N__66233),
            .I(N__66224));
    InMux I__15921 (
            .O(N__66230),
            .I(N__66221));
    Sp12to4 I__15920 (
            .O(N__66227),
            .I(N__66216));
    Sp12to4 I__15919 (
            .O(N__66224),
            .I(N__66216));
    LocalMux I__15918 (
            .O(N__66221),
            .I(\c0.data_in_frame_20_1 ));
    Odrv12 I__15917 (
            .O(N__66216),
            .I(\c0.data_in_frame_20_1 ));
    CascadeMux I__15916 (
            .O(N__66211),
            .I(N__66206));
    InMux I__15915 (
            .O(N__66210),
            .I(N__66198));
    InMux I__15914 (
            .O(N__66209),
            .I(N__66198));
    InMux I__15913 (
            .O(N__66206),
            .I(N__66195));
    CascadeMux I__15912 (
            .O(N__66205),
            .I(N__66190));
    CascadeMux I__15911 (
            .O(N__66204),
            .I(N__66181));
    CascadeMux I__15910 (
            .O(N__66203),
            .I(N__66178));
    LocalMux I__15909 (
            .O(N__66198),
            .I(N__66172));
    LocalMux I__15908 (
            .O(N__66195),
            .I(N__66172));
    InMux I__15907 (
            .O(N__66194),
            .I(N__66169));
    InMux I__15906 (
            .O(N__66193),
            .I(N__66166));
    InMux I__15905 (
            .O(N__66190),
            .I(N__66163));
    CascadeMux I__15904 (
            .O(N__66189),
            .I(N__66159));
    CascadeMux I__15903 (
            .O(N__66188),
            .I(N__66150));
    CascadeMux I__15902 (
            .O(N__66187),
            .I(N__66147));
    CascadeMux I__15901 (
            .O(N__66186),
            .I(N__66141));
    InMux I__15900 (
            .O(N__66185),
            .I(N__66136));
    InMux I__15899 (
            .O(N__66184),
            .I(N__66133));
    InMux I__15898 (
            .O(N__66181),
            .I(N__66126));
    InMux I__15897 (
            .O(N__66178),
            .I(N__66126));
    InMux I__15896 (
            .O(N__66177),
            .I(N__66126));
    Span4Mux_v I__15895 (
            .O(N__66172),
            .I(N__66122));
    LocalMux I__15894 (
            .O(N__66169),
            .I(N__66117));
    LocalMux I__15893 (
            .O(N__66166),
            .I(N__66114));
    LocalMux I__15892 (
            .O(N__66163),
            .I(N__66111));
    InMux I__15891 (
            .O(N__66162),
            .I(N__66102));
    InMux I__15890 (
            .O(N__66159),
            .I(N__66102));
    InMux I__15889 (
            .O(N__66158),
            .I(N__66102));
    InMux I__15888 (
            .O(N__66157),
            .I(N__66102));
    InMux I__15887 (
            .O(N__66156),
            .I(N__66099));
    InMux I__15886 (
            .O(N__66155),
            .I(N__66096));
    InMux I__15885 (
            .O(N__66154),
            .I(N__66093));
    InMux I__15884 (
            .O(N__66153),
            .I(N__66084));
    InMux I__15883 (
            .O(N__66150),
            .I(N__66084));
    InMux I__15882 (
            .O(N__66147),
            .I(N__66084));
    InMux I__15881 (
            .O(N__66146),
            .I(N__66084));
    InMux I__15880 (
            .O(N__66145),
            .I(N__66081));
    InMux I__15879 (
            .O(N__66144),
            .I(N__66078));
    InMux I__15878 (
            .O(N__66141),
            .I(N__66071));
    InMux I__15877 (
            .O(N__66140),
            .I(N__66071));
    InMux I__15876 (
            .O(N__66139),
            .I(N__66071));
    LocalMux I__15875 (
            .O(N__66136),
            .I(N__66068));
    LocalMux I__15874 (
            .O(N__66133),
            .I(N__66061));
    LocalMux I__15873 (
            .O(N__66126),
            .I(N__66061));
    InMux I__15872 (
            .O(N__66125),
            .I(N__66057));
    Span4Mux_h I__15871 (
            .O(N__66122),
            .I(N__66054));
    InMux I__15870 (
            .O(N__66121),
            .I(N__66051));
    CascadeMux I__15869 (
            .O(N__66120),
            .I(N__66047));
    Span4Mux_h I__15868 (
            .O(N__66117),
            .I(N__66040));
    Span4Mux_h I__15867 (
            .O(N__66114),
            .I(N__66040));
    Span4Mux_v I__15866 (
            .O(N__66111),
            .I(N__66033));
    LocalMux I__15865 (
            .O(N__66102),
            .I(N__66033));
    LocalMux I__15864 (
            .O(N__66099),
            .I(N__66026));
    LocalMux I__15863 (
            .O(N__66096),
            .I(N__66026));
    LocalMux I__15862 (
            .O(N__66093),
            .I(N__66026));
    LocalMux I__15861 (
            .O(N__66084),
            .I(N__66023));
    LocalMux I__15860 (
            .O(N__66081),
            .I(N__66020));
    LocalMux I__15859 (
            .O(N__66078),
            .I(N__66013));
    LocalMux I__15858 (
            .O(N__66071),
            .I(N__66013));
    Span4Mux_v I__15857 (
            .O(N__66068),
            .I(N__66013));
    InMux I__15856 (
            .O(N__66067),
            .I(N__66008));
    CascadeMux I__15855 (
            .O(N__66066),
            .I(N__66004));
    Span4Mux_v I__15854 (
            .O(N__66061),
            .I(N__66001));
    InMux I__15853 (
            .O(N__66060),
            .I(N__65998));
    LocalMux I__15852 (
            .O(N__66057),
            .I(N__65995));
    Span4Mux_v I__15851 (
            .O(N__66054),
            .I(N__65992));
    LocalMux I__15850 (
            .O(N__66051),
            .I(N__65989));
    InMux I__15849 (
            .O(N__66050),
            .I(N__65986));
    InMux I__15848 (
            .O(N__66047),
            .I(N__65979));
    InMux I__15847 (
            .O(N__66046),
            .I(N__65979));
    InMux I__15846 (
            .O(N__66045),
            .I(N__65979));
    Span4Mux_h I__15845 (
            .O(N__66040),
            .I(N__65976));
    InMux I__15844 (
            .O(N__66039),
            .I(N__65971));
    InMux I__15843 (
            .O(N__66038),
            .I(N__65971));
    Span4Mux_v I__15842 (
            .O(N__66033),
            .I(N__65968));
    Span4Mux_v I__15841 (
            .O(N__66026),
            .I(N__65965));
    Span4Mux_v I__15840 (
            .O(N__66023),
            .I(N__65958));
    Span4Mux_h I__15839 (
            .O(N__66020),
            .I(N__65958));
    Span4Mux_v I__15838 (
            .O(N__66013),
            .I(N__65958));
    InMux I__15837 (
            .O(N__66012),
            .I(N__65955));
    InMux I__15836 (
            .O(N__66011),
            .I(N__65952));
    LocalMux I__15835 (
            .O(N__66008),
            .I(N__65949));
    InMux I__15834 (
            .O(N__66007),
            .I(N__65944));
    InMux I__15833 (
            .O(N__66004),
            .I(N__65944));
    Span4Mux_v I__15832 (
            .O(N__66001),
            .I(N__65941));
    LocalMux I__15831 (
            .O(N__65998),
            .I(N__65936));
    Span4Mux_h I__15830 (
            .O(N__65995),
            .I(N__65936));
    Sp12to4 I__15829 (
            .O(N__65992),
            .I(N__65933));
    Span4Mux_h I__15828 (
            .O(N__65989),
            .I(N__65930));
    LocalMux I__15827 (
            .O(N__65986),
            .I(N__65921));
    LocalMux I__15826 (
            .O(N__65979),
            .I(N__65921));
    Span4Mux_h I__15825 (
            .O(N__65976),
            .I(N__65921));
    LocalMux I__15824 (
            .O(N__65971),
            .I(N__65921));
    Span4Mux_h I__15823 (
            .O(N__65968),
            .I(N__65918));
    Span4Mux_v I__15822 (
            .O(N__65965),
            .I(N__65913));
    Span4Mux_v I__15821 (
            .O(N__65958),
            .I(N__65913));
    LocalMux I__15820 (
            .O(N__65955),
            .I(N__65904));
    LocalMux I__15819 (
            .O(N__65952),
            .I(N__65904));
    Sp12to4 I__15818 (
            .O(N__65949),
            .I(N__65904));
    LocalMux I__15817 (
            .O(N__65944),
            .I(N__65904));
    Span4Mux_h I__15816 (
            .O(N__65941),
            .I(N__65901));
    Sp12to4 I__15815 (
            .O(N__65936),
            .I(N__65894));
    Span12Mux_h I__15814 (
            .O(N__65933),
            .I(N__65894));
    Sp12to4 I__15813 (
            .O(N__65930),
            .I(N__65894));
    Span4Mux_v I__15812 (
            .O(N__65921),
            .I(N__65891));
    Span4Mux_v I__15811 (
            .O(N__65918),
            .I(N__65888));
    Span4Mux_h I__15810 (
            .O(N__65913),
            .I(N__65885));
    Span12Mux_h I__15809 (
            .O(N__65904),
            .I(N__65878));
    Sp12to4 I__15808 (
            .O(N__65901),
            .I(N__65878));
    Span12Mux_v I__15807 (
            .O(N__65894),
            .I(N__65878));
    Odrv4 I__15806 (
            .O(N__65891),
            .I(\c0.n12_adj_3265 ));
    Odrv4 I__15805 (
            .O(N__65888),
            .I(\c0.n12_adj_3265 ));
    Odrv4 I__15804 (
            .O(N__65885),
            .I(\c0.n12_adj_3265 ));
    Odrv12 I__15803 (
            .O(N__65878),
            .I(\c0.n12_adj_3265 ));
    CascadeMux I__15802 (
            .O(N__65869),
            .I(N__65865));
    InMux I__15801 (
            .O(N__65868),
            .I(N__65860));
    InMux I__15800 (
            .O(N__65865),
            .I(N__65857));
    InMux I__15799 (
            .O(N__65864),
            .I(N__65854));
    CascadeMux I__15798 (
            .O(N__65863),
            .I(N__65850));
    LocalMux I__15797 (
            .O(N__65860),
            .I(N__65846));
    LocalMux I__15796 (
            .O(N__65857),
            .I(N__65843));
    LocalMux I__15795 (
            .O(N__65854),
            .I(N__65840));
    InMux I__15794 (
            .O(N__65853),
            .I(N__65837));
    InMux I__15793 (
            .O(N__65850),
            .I(N__65834));
    InMux I__15792 (
            .O(N__65849),
            .I(N__65831));
    Span4Mux_v I__15791 (
            .O(N__65846),
            .I(N__65828));
    Span4Mux_v I__15790 (
            .O(N__65843),
            .I(N__65823));
    Span4Mux_v I__15789 (
            .O(N__65840),
            .I(N__65823));
    LocalMux I__15788 (
            .O(N__65837),
            .I(N__65818));
    LocalMux I__15787 (
            .O(N__65834),
            .I(N__65818));
    LocalMux I__15786 (
            .O(N__65831),
            .I(N__65815));
    Span4Mux_h I__15785 (
            .O(N__65828),
            .I(N__65812));
    Span4Mux_h I__15784 (
            .O(N__65823),
            .I(N__65809));
    Span4Mux_v I__15783 (
            .O(N__65818),
            .I(N__65806));
    Odrv12 I__15782 (
            .O(N__65815),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__15781 (
            .O(N__65812),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__15780 (
            .O(N__65809),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__15779 (
            .O(N__65806),
            .I(\c0.data_in_frame_12_3 ));
    InMux I__15778 (
            .O(N__65797),
            .I(N__65792));
    InMux I__15777 (
            .O(N__65796),
            .I(N__65789));
    InMux I__15776 (
            .O(N__65795),
            .I(N__65786));
    LocalMux I__15775 (
            .O(N__65792),
            .I(N__65783));
    LocalMux I__15774 (
            .O(N__65789),
            .I(N__65775));
    LocalMux I__15773 (
            .O(N__65786),
            .I(N__65775));
    Span4Mux_v I__15772 (
            .O(N__65783),
            .I(N__65772));
    InMux I__15771 (
            .O(N__65782),
            .I(N__65769));
    InMux I__15770 (
            .O(N__65781),
            .I(N__65766));
    InMux I__15769 (
            .O(N__65780),
            .I(N__65763));
    Span4Mux_v I__15768 (
            .O(N__65775),
            .I(N__65759));
    Sp12to4 I__15767 (
            .O(N__65772),
            .I(N__65752));
    LocalMux I__15766 (
            .O(N__65769),
            .I(N__65752));
    LocalMux I__15765 (
            .O(N__65766),
            .I(N__65752));
    LocalMux I__15764 (
            .O(N__65763),
            .I(N__65749));
    CascadeMux I__15763 (
            .O(N__65762),
            .I(N__65746));
    Span4Mux_h I__15762 (
            .O(N__65759),
            .I(N__65743));
    Span12Mux_h I__15761 (
            .O(N__65752),
            .I(N__65738));
    Sp12to4 I__15760 (
            .O(N__65749),
            .I(N__65738));
    InMux I__15759 (
            .O(N__65746),
            .I(N__65735));
    Span4Mux_v I__15758 (
            .O(N__65743),
            .I(N__65732));
    Span12Mux_v I__15757 (
            .O(N__65738),
            .I(N__65729));
    LocalMux I__15756 (
            .O(N__65735),
            .I(data_in_frame_19_2));
    Odrv4 I__15755 (
            .O(N__65732),
            .I(data_in_frame_19_2));
    Odrv12 I__15754 (
            .O(N__65729),
            .I(data_in_frame_19_2));
    InMux I__15753 (
            .O(N__65722),
            .I(N__65719));
    LocalMux I__15752 (
            .O(N__65719),
            .I(N__65716));
    Span4Mux_h I__15751 (
            .O(N__65716),
            .I(N__65712));
    InMux I__15750 (
            .O(N__65715),
            .I(N__65708));
    Span4Mux_h I__15749 (
            .O(N__65712),
            .I(N__65705));
    InMux I__15748 (
            .O(N__65711),
            .I(N__65702));
    LocalMux I__15747 (
            .O(N__65708),
            .I(data_in_frame_19_5));
    Odrv4 I__15746 (
            .O(N__65705),
            .I(data_in_frame_19_5));
    LocalMux I__15745 (
            .O(N__65702),
            .I(data_in_frame_19_5));
    InMux I__15744 (
            .O(N__65695),
            .I(N__65690));
    InMux I__15743 (
            .O(N__65694),
            .I(N__65687));
    InMux I__15742 (
            .O(N__65693),
            .I(N__65684));
    LocalMux I__15741 (
            .O(N__65690),
            .I(N__65681));
    LocalMux I__15740 (
            .O(N__65687),
            .I(N__65675));
    LocalMux I__15739 (
            .O(N__65684),
            .I(N__65675));
    Span4Mux_h I__15738 (
            .O(N__65681),
            .I(N__65671));
    InMux I__15737 (
            .O(N__65680),
            .I(N__65668));
    Span4Mux_h I__15736 (
            .O(N__65675),
            .I(N__65665));
    CascadeMux I__15735 (
            .O(N__65674),
            .I(N__65662));
    Span4Mux_v I__15734 (
            .O(N__65671),
            .I(N__65658));
    LocalMux I__15733 (
            .O(N__65668),
            .I(N__65655));
    Span4Mux_h I__15732 (
            .O(N__65665),
            .I(N__65652));
    InMux I__15731 (
            .O(N__65662),
            .I(N__65649));
    InMux I__15730 (
            .O(N__65661),
            .I(N__65646));
    Span4Mux_v I__15729 (
            .O(N__65658),
            .I(N__65643));
    Span4Mux_h I__15728 (
            .O(N__65655),
            .I(N__65638));
    Span4Mux_v I__15727 (
            .O(N__65652),
            .I(N__65638));
    LocalMux I__15726 (
            .O(N__65649),
            .I(N__65635));
    LocalMux I__15725 (
            .O(N__65646),
            .I(data_in_frame_19_1));
    Odrv4 I__15724 (
            .O(N__65643),
            .I(data_in_frame_19_1));
    Odrv4 I__15723 (
            .O(N__65638),
            .I(data_in_frame_19_1));
    Odrv12 I__15722 (
            .O(N__65635),
            .I(data_in_frame_19_1));
    InMux I__15721 (
            .O(N__65626),
            .I(N__65623));
    LocalMux I__15720 (
            .O(N__65623),
            .I(N__65620));
    Span4Mux_h I__15719 (
            .O(N__65620),
            .I(N__65615));
    InMux I__15718 (
            .O(N__65619),
            .I(N__65610));
    InMux I__15717 (
            .O(N__65618),
            .I(N__65610));
    Odrv4 I__15716 (
            .O(N__65615),
            .I(\c0.n6166 ));
    LocalMux I__15715 (
            .O(N__65610),
            .I(\c0.n6166 ));
    InMux I__15714 (
            .O(N__65605),
            .I(N__65602));
    LocalMux I__15713 (
            .O(N__65602),
            .I(N__65599));
    Span4Mux_h I__15712 (
            .O(N__65599),
            .I(N__65591));
    InMux I__15711 (
            .O(N__65598),
            .I(N__65587));
    InMux I__15710 (
            .O(N__65597),
            .I(N__65584));
    InMux I__15709 (
            .O(N__65596),
            .I(N__65581));
    InMux I__15708 (
            .O(N__65595),
            .I(N__65575));
    InMux I__15707 (
            .O(N__65594),
            .I(N__65575));
    Span4Mux_h I__15706 (
            .O(N__65591),
            .I(N__65572));
    InMux I__15705 (
            .O(N__65590),
            .I(N__65569));
    LocalMux I__15704 (
            .O(N__65587),
            .I(N__65566));
    LocalMux I__15703 (
            .O(N__65584),
            .I(N__65563));
    LocalMux I__15702 (
            .O(N__65581),
            .I(N__65560));
    InMux I__15701 (
            .O(N__65580),
            .I(N__65557));
    LocalMux I__15700 (
            .O(N__65575),
            .I(N__65554));
    Sp12to4 I__15699 (
            .O(N__65572),
            .I(N__65551));
    LocalMux I__15698 (
            .O(N__65569),
            .I(N__65544));
    Sp12to4 I__15697 (
            .O(N__65566),
            .I(N__65544));
    Sp12to4 I__15696 (
            .O(N__65563),
            .I(N__65544));
    Sp12to4 I__15695 (
            .O(N__65560),
            .I(N__65541));
    LocalMux I__15694 (
            .O(N__65557),
            .I(N__65532));
    Span12Mux_v I__15693 (
            .O(N__65554),
            .I(N__65532));
    Span12Mux_v I__15692 (
            .O(N__65551),
            .I(N__65532));
    Span12Mux_v I__15691 (
            .O(N__65544),
            .I(N__65532));
    Odrv12 I__15690 (
            .O(N__65541),
            .I(n19130));
    Odrv12 I__15689 (
            .O(N__65532),
            .I(n19130));
    InMux I__15688 (
            .O(N__65527),
            .I(N__65522));
    CascadeMux I__15687 (
            .O(N__65526),
            .I(N__65516));
    InMux I__15686 (
            .O(N__65525),
            .I(N__65512));
    LocalMux I__15685 (
            .O(N__65522),
            .I(N__65509));
    InMux I__15684 (
            .O(N__65521),
            .I(N__65504));
    InMux I__15683 (
            .O(N__65520),
            .I(N__65504));
    InMux I__15682 (
            .O(N__65519),
            .I(N__65499));
    InMux I__15681 (
            .O(N__65516),
            .I(N__65499));
    InMux I__15680 (
            .O(N__65515),
            .I(N__65496));
    LocalMux I__15679 (
            .O(N__65512),
            .I(N__65490));
    Span4Mux_h I__15678 (
            .O(N__65509),
            .I(N__65485));
    LocalMux I__15677 (
            .O(N__65504),
            .I(N__65485));
    LocalMux I__15676 (
            .O(N__65499),
            .I(N__65482));
    LocalMux I__15675 (
            .O(N__65496),
            .I(N__65479));
    InMux I__15674 (
            .O(N__65495),
            .I(N__65474));
    InMux I__15673 (
            .O(N__65494),
            .I(N__65474));
    InMux I__15672 (
            .O(N__65493),
            .I(N__65471));
    Span4Mux_h I__15671 (
            .O(N__65490),
            .I(N__65466));
    Span4Mux_v I__15670 (
            .O(N__65485),
            .I(N__65466));
    Span4Mux_h I__15669 (
            .O(N__65482),
            .I(N__65459));
    Span4Mux_h I__15668 (
            .O(N__65479),
            .I(N__65459));
    LocalMux I__15667 (
            .O(N__65474),
            .I(N__65459));
    LocalMux I__15666 (
            .O(N__65471),
            .I(data_in_frame_16_2));
    Odrv4 I__15665 (
            .O(N__65466),
            .I(data_in_frame_16_2));
    Odrv4 I__15664 (
            .O(N__65459),
            .I(data_in_frame_16_2));
    InMux I__15663 (
            .O(N__65452),
            .I(N__65449));
    LocalMux I__15662 (
            .O(N__65449),
            .I(N__65445));
    InMux I__15661 (
            .O(N__65448),
            .I(N__65442));
    Span4Mux_v I__15660 (
            .O(N__65445),
            .I(N__65439));
    LocalMux I__15659 (
            .O(N__65442),
            .I(\c0.data_in_frame_28_5 ));
    Odrv4 I__15658 (
            .O(N__65439),
            .I(\c0.data_in_frame_28_5 ));
    InMux I__15657 (
            .O(N__65434),
            .I(N__65430));
    CascadeMux I__15656 (
            .O(N__65433),
            .I(N__65426));
    LocalMux I__15655 (
            .O(N__65430),
            .I(N__65423));
    InMux I__15654 (
            .O(N__65429),
            .I(N__65420));
    InMux I__15653 (
            .O(N__65426),
            .I(N__65417));
    Span4Mux_h I__15652 (
            .O(N__65423),
            .I(N__65412));
    LocalMux I__15651 (
            .O(N__65420),
            .I(N__65412));
    LocalMux I__15650 (
            .O(N__65417),
            .I(\c0.n19381 ));
    Odrv4 I__15649 (
            .O(N__65412),
            .I(\c0.n19381 ));
    InMux I__15648 (
            .O(N__65407),
            .I(N__65403));
    InMux I__15647 (
            .O(N__65406),
            .I(N__65400));
    LocalMux I__15646 (
            .O(N__65403),
            .I(N__65394));
    LocalMux I__15645 (
            .O(N__65400),
            .I(N__65391));
    InMux I__15644 (
            .O(N__65399),
            .I(N__65388));
    InMux I__15643 (
            .O(N__65398),
            .I(N__65385));
    CascadeMux I__15642 (
            .O(N__65397),
            .I(N__65382));
    Span4Mux_h I__15641 (
            .O(N__65394),
            .I(N__65379));
    Span4Mux_h I__15640 (
            .O(N__65391),
            .I(N__65374));
    LocalMux I__15639 (
            .O(N__65388),
            .I(N__65374));
    LocalMux I__15638 (
            .O(N__65385),
            .I(N__65371));
    InMux I__15637 (
            .O(N__65382),
            .I(N__65368));
    Span4Mux_v I__15636 (
            .O(N__65379),
            .I(N__65365));
    Span4Mux_v I__15635 (
            .O(N__65374),
            .I(N__65362));
    Span4Mux_v I__15634 (
            .O(N__65371),
            .I(N__65359));
    LocalMux I__15633 (
            .O(N__65368),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__15632 (
            .O(N__65365),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__15631 (
            .O(N__65362),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__15630 (
            .O(N__65359),
            .I(\c0.data_in_frame_7_0 ));
    CascadeMux I__15629 (
            .O(N__65350),
            .I(N__65347));
    InMux I__15628 (
            .O(N__65347),
            .I(N__65344));
    LocalMux I__15627 (
            .O(N__65344),
            .I(N__65340));
    InMux I__15626 (
            .O(N__65343),
            .I(N__65337));
    Span4Mux_h I__15625 (
            .O(N__65340),
            .I(N__65334));
    LocalMux I__15624 (
            .O(N__65337),
            .I(N__65331));
    Odrv4 I__15623 (
            .O(N__65334),
            .I(\c0.n7_adj_3355 ));
    Odrv12 I__15622 (
            .O(N__65331),
            .I(\c0.n7_adj_3355 ));
    CascadeMux I__15621 (
            .O(N__65326),
            .I(N__65322));
    InMux I__15620 (
            .O(N__65325),
            .I(N__65317));
    InMux I__15619 (
            .O(N__65322),
            .I(N__65314));
    InMux I__15618 (
            .O(N__65321),
            .I(N__65309));
    InMux I__15617 (
            .O(N__65320),
            .I(N__65309));
    LocalMux I__15616 (
            .O(N__65317),
            .I(N__65306));
    LocalMux I__15615 (
            .O(N__65314),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__15614 (
            .O(N__65309),
            .I(\c0.data_in_frame_17_5 ));
    Odrv4 I__15613 (
            .O(N__65306),
            .I(\c0.data_in_frame_17_5 ));
    InMux I__15612 (
            .O(N__65299),
            .I(N__65293));
    InMux I__15611 (
            .O(N__65298),
            .I(N__65293));
    LocalMux I__15610 (
            .O(N__65293),
            .I(N__65289));
    InMux I__15609 (
            .O(N__65292),
            .I(N__65286));
    Odrv4 I__15608 (
            .O(N__65289),
            .I(\c0.n11590 ));
    LocalMux I__15607 (
            .O(N__65286),
            .I(\c0.n11590 ));
    CascadeMux I__15606 (
            .O(N__65281),
            .I(N__65278));
    InMux I__15605 (
            .O(N__65278),
            .I(N__65275));
    LocalMux I__15604 (
            .O(N__65275),
            .I(N__65272));
    Span4Mux_v I__15603 (
            .O(N__65272),
            .I(N__65269));
    Span4Mux_h I__15602 (
            .O(N__65269),
            .I(N__65266));
    Odrv4 I__15601 (
            .O(N__65266),
            .I(\c0.n14_adj_3449 ));
    InMux I__15600 (
            .O(N__65263),
            .I(N__65253));
    InMux I__15599 (
            .O(N__65262),
            .I(N__65253));
    InMux I__15598 (
            .O(N__65261),
            .I(N__65250));
    InMux I__15597 (
            .O(N__65260),
            .I(N__65243));
    InMux I__15596 (
            .O(N__65259),
            .I(N__65235));
    CascadeMux I__15595 (
            .O(N__65258),
            .I(N__65231));
    LocalMux I__15594 (
            .O(N__65253),
            .I(N__65227));
    LocalMux I__15593 (
            .O(N__65250),
            .I(N__65223));
    InMux I__15592 (
            .O(N__65249),
            .I(N__65218));
    InMux I__15591 (
            .O(N__65248),
            .I(N__65218));
    InMux I__15590 (
            .O(N__65247),
            .I(N__65212));
    InMux I__15589 (
            .O(N__65246),
            .I(N__65212));
    LocalMux I__15588 (
            .O(N__65243),
            .I(N__65209));
    InMux I__15587 (
            .O(N__65242),
            .I(N__65206));
    InMux I__15586 (
            .O(N__65241),
            .I(N__65203));
    InMux I__15585 (
            .O(N__65240),
            .I(N__65199));
    InMux I__15584 (
            .O(N__65239),
            .I(N__65195));
    InMux I__15583 (
            .O(N__65238),
            .I(N__65192));
    LocalMux I__15582 (
            .O(N__65235),
            .I(N__65186));
    InMux I__15581 (
            .O(N__65234),
            .I(N__65179));
    InMux I__15580 (
            .O(N__65231),
            .I(N__65179));
    InMux I__15579 (
            .O(N__65230),
            .I(N__65179));
    Span4Mux_h I__15578 (
            .O(N__65227),
            .I(N__65176));
    InMux I__15577 (
            .O(N__65226),
            .I(N__65173));
    Span4Mux_v I__15576 (
            .O(N__65223),
            .I(N__65169));
    LocalMux I__15575 (
            .O(N__65218),
            .I(N__65166));
    InMux I__15574 (
            .O(N__65217),
            .I(N__65163));
    LocalMux I__15573 (
            .O(N__65212),
            .I(N__65160));
    Span4Mux_h I__15572 (
            .O(N__65209),
            .I(N__65155));
    LocalMux I__15571 (
            .O(N__65206),
            .I(N__65155));
    LocalMux I__15570 (
            .O(N__65203),
            .I(N__65152));
    InMux I__15569 (
            .O(N__65202),
            .I(N__65149));
    LocalMux I__15568 (
            .O(N__65199),
            .I(N__65144));
    InMux I__15567 (
            .O(N__65198),
            .I(N__65141));
    LocalMux I__15566 (
            .O(N__65195),
            .I(N__65136));
    LocalMux I__15565 (
            .O(N__65192),
            .I(N__65136));
    InMux I__15564 (
            .O(N__65191),
            .I(N__65129));
    InMux I__15563 (
            .O(N__65190),
            .I(N__65129));
    InMux I__15562 (
            .O(N__65189),
            .I(N__65129));
    Span4Mux_v I__15561 (
            .O(N__65186),
            .I(N__65124));
    LocalMux I__15560 (
            .O(N__65179),
            .I(N__65124));
    Span4Mux_v I__15559 (
            .O(N__65176),
            .I(N__65119));
    LocalMux I__15558 (
            .O(N__65173),
            .I(N__65119));
    InMux I__15557 (
            .O(N__65172),
            .I(N__65114));
    Span4Mux_h I__15556 (
            .O(N__65169),
            .I(N__65109));
    Span4Mux_h I__15555 (
            .O(N__65166),
            .I(N__65109));
    LocalMux I__15554 (
            .O(N__65163),
            .I(N__65104));
    Span4Mux_h I__15553 (
            .O(N__65160),
            .I(N__65104));
    Span4Mux_v I__15552 (
            .O(N__65155),
            .I(N__65101));
    Span4Mux_v I__15551 (
            .O(N__65152),
            .I(N__65098));
    LocalMux I__15550 (
            .O(N__65149),
            .I(N__65095));
    InMux I__15549 (
            .O(N__65148),
            .I(N__65091));
    InMux I__15548 (
            .O(N__65147),
            .I(N__65088));
    Span4Mux_v I__15547 (
            .O(N__65144),
            .I(N__65085));
    LocalMux I__15546 (
            .O(N__65141),
            .I(N__65082));
    Span4Mux_v I__15545 (
            .O(N__65136),
            .I(N__65079));
    LocalMux I__15544 (
            .O(N__65129),
            .I(N__65074));
    Span4Mux_v I__15543 (
            .O(N__65124),
            .I(N__65074));
    Span4Mux_h I__15542 (
            .O(N__65119),
            .I(N__65071));
    InMux I__15541 (
            .O(N__65118),
            .I(N__65064));
    InMux I__15540 (
            .O(N__65117),
            .I(N__65064));
    LocalMux I__15539 (
            .O(N__65114),
            .I(N__65057));
    Span4Mux_h I__15538 (
            .O(N__65109),
            .I(N__65057));
    Span4Mux_h I__15537 (
            .O(N__65104),
            .I(N__65057));
    Sp12to4 I__15536 (
            .O(N__65101),
            .I(N__65052));
    Sp12to4 I__15535 (
            .O(N__65098),
            .I(N__65052));
    Span4Mux_v I__15534 (
            .O(N__65095),
            .I(N__65049));
    InMux I__15533 (
            .O(N__65094),
            .I(N__65046));
    LocalMux I__15532 (
            .O(N__65091),
            .I(N__65037));
    LocalMux I__15531 (
            .O(N__65088),
            .I(N__65037));
    Span4Mux_h I__15530 (
            .O(N__65085),
            .I(N__65037));
    Span4Mux_v I__15529 (
            .O(N__65082),
            .I(N__65037));
    Span4Mux_v I__15528 (
            .O(N__65079),
            .I(N__65034));
    Span4Mux_v I__15527 (
            .O(N__65074),
            .I(N__65031));
    Sp12to4 I__15526 (
            .O(N__65071),
            .I(N__65028));
    InMux I__15525 (
            .O(N__65070),
            .I(N__65025));
    InMux I__15524 (
            .O(N__65069),
            .I(N__65022));
    LocalMux I__15523 (
            .O(N__65064),
            .I(N__65019));
    Sp12to4 I__15522 (
            .O(N__65057),
            .I(N__65014));
    Span12Mux_h I__15521 (
            .O(N__65052),
            .I(N__65014));
    Span4Mux_h I__15520 (
            .O(N__65049),
            .I(N__65011));
    LocalMux I__15519 (
            .O(N__65046),
            .I(N__65000));
    Sp12to4 I__15518 (
            .O(N__65037),
            .I(N__65000));
    Sp12to4 I__15517 (
            .O(N__65034),
            .I(N__65000));
    Sp12to4 I__15516 (
            .O(N__65031),
            .I(N__65000));
    Span12Mux_v I__15515 (
            .O(N__65028),
            .I(N__65000));
    LocalMux I__15514 (
            .O(N__65025),
            .I(N__64991));
    LocalMux I__15513 (
            .O(N__65022),
            .I(N__64991));
    Span12Mux_h I__15512 (
            .O(N__65019),
            .I(N__64991));
    Span12Mux_v I__15511 (
            .O(N__65014),
            .I(N__64991));
    Odrv4 I__15510 (
            .O(N__65011),
            .I(rx_data_0));
    Odrv12 I__15509 (
            .O(N__65000),
            .I(rx_data_0));
    Odrv12 I__15508 (
            .O(N__64991),
            .I(rx_data_0));
    InMux I__15507 (
            .O(N__64984),
            .I(N__64980));
    InMux I__15506 (
            .O(N__64983),
            .I(N__64976));
    LocalMux I__15505 (
            .O(N__64980),
            .I(N__64973));
    InMux I__15504 (
            .O(N__64979),
            .I(N__64969));
    LocalMux I__15503 (
            .O(N__64976),
            .I(N__64966));
    Span4Mux_v I__15502 (
            .O(N__64973),
            .I(N__64963));
    InMux I__15501 (
            .O(N__64972),
            .I(N__64960));
    LocalMux I__15500 (
            .O(N__64969),
            .I(\c0.data_in_frame_15_1 ));
    Odrv12 I__15499 (
            .O(N__64966),
            .I(\c0.data_in_frame_15_1 ));
    Odrv4 I__15498 (
            .O(N__64963),
            .I(\c0.data_in_frame_15_1 ));
    LocalMux I__15497 (
            .O(N__64960),
            .I(\c0.data_in_frame_15_1 ));
    InMux I__15496 (
            .O(N__64951),
            .I(N__64946));
    InMux I__15495 (
            .O(N__64950),
            .I(N__64943));
    InMux I__15494 (
            .O(N__64949),
            .I(N__64939));
    LocalMux I__15493 (
            .O(N__64946),
            .I(N__64936));
    LocalMux I__15492 (
            .O(N__64943),
            .I(N__64933));
    CascadeMux I__15491 (
            .O(N__64942),
            .I(N__64930));
    LocalMux I__15490 (
            .O(N__64939),
            .I(N__64927));
    Span4Mux_h I__15489 (
            .O(N__64936),
            .I(N__64924));
    Span4Mux_v I__15488 (
            .O(N__64933),
            .I(N__64921));
    InMux I__15487 (
            .O(N__64930),
            .I(N__64917));
    Span4Mux_h I__15486 (
            .O(N__64927),
            .I(N__64910));
    Span4Mux_v I__15485 (
            .O(N__64924),
            .I(N__64910));
    Span4Mux_v I__15484 (
            .O(N__64921),
            .I(N__64910));
    InMux I__15483 (
            .O(N__64920),
            .I(N__64907));
    LocalMux I__15482 (
            .O(N__64917),
            .I(\c0.data_in_frame_14_7 ));
    Odrv4 I__15481 (
            .O(N__64910),
            .I(\c0.data_in_frame_14_7 ));
    LocalMux I__15480 (
            .O(N__64907),
            .I(\c0.data_in_frame_14_7 ));
    InMux I__15479 (
            .O(N__64900),
            .I(N__64896));
    InMux I__15478 (
            .O(N__64899),
            .I(N__64893));
    LocalMux I__15477 (
            .O(N__64896),
            .I(N__64889));
    LocalMux I__15476 (
            .O(N__64893),
            .I(N__64883));
    InMux I__15475 (
            .O(N__64892),
            .I(N__64880));
    Span4Mux_h I__15474 (
            .O(N__64889),
            .I(N__64877));
    InMux I__15473 (
            .O(N__64888),
            .I(N__64874));
    CascadeMux I__15472 (
            .O(N__64887),
            .I(N__64871));
    InMux I__15471 (
            .O(N__64886),
            .I(N__64868));
    Span4Mux_v I__15470 (
            .O(N__64883),
            .I(N__64865));
    LocalMux I__15469 (
            .O(N__64880),
            .I(N__64860));
    Span4Mux_v I__15468 (
            .O(N__64877),
            .I(N__64860));
    LocalMux I__15467 (
            .O(N__64874),
            .I(N__64857));
    InMux I__15466 (
            .O(N__64871),
            .I(N__64854));
    LocalMux I__15465 (
            .O(N__64868),
            .I(N__64849));
    Span4Mux_h I__15464 (
            .O(N__64865),
            .I(N__64849));
    Span4Mux_h I__15463 (
            .O(N__64860),
            .I(N__64846));
    Span12Mux_h I__15462 (
            .O(N__64857),
            .I(N__64843));
    LocalMux I__15461 (
            .O(N__64854),
            .I(\c0.data_in_frame_14_6 ));
    Odrv4 I__15460 (
            .O(N__64849),
            .I(\c0.data_in_frame_14_6 ));
    Odrv4 I__15459 (
            .O(N__64846),
            .I(\c0.data_in_frame_14_6 ));
    Odrv12 I__15458 (
            .O(N__64843),
            .I(\c0.data_in_frame_14_6 ));
    InMux I__15457 (
            .O(N__64834),
            .I(N__64827));
    InMux I__15456 (
            .O(N__64833),
            .I(N__64822));
    InMux I__15455 (
            .O(N__64832),
            .I(N__64822));
    CascadeMux I__15454 (
            .O(N__64831),
            .I(N__64818));
    InMux I__15453 (
            .O(N__64830),
            .I(N__64815));
    LocalMux I__15452 (
            .O(N__64827),
            .I(N__64812));
    LocalMux I__15451 (
            .O(N__64822),
            .I(N__64809));
    CascadeMux I__15450 (
            .O(N__64821),
            .I(N__64806));
    InMux I__15449 (
            .O(N__64818),
            .I(N__64803));
    LocalMux I__15448 (
            .O(N__64815),
            .I(N__64800));
    Span4Mux_v I__15447 (
            .O(N__64812),
            .I(N__64795));
    Span4Mux_v I__15446 (
            .O(N__64809),
            .I(N__64795));
    InMux I__15445 (
            .O(N__64806),
            .I(N__64792));
    LocalMux I__15444 (
            .O(N__64803),
            .I(N__64789));
    Span4Mux_v I__15443 (
            .O(N__64800),
            .I(N__64786));
    Sp12to4 I__15442 (
            .O(N__64795),
            .I(N__64781));
    LocalMux I__15441 (
            .O(N__64792),
            .I(N__64781));
    Span4Mux_h I__15440 (
            .O(N__64789),
            .I(N__64776));
    Span4Mux_h I__15439 (
            .O(N__64786),
            .I(N__64776));
    Odrv12 I__15438 (
            .O(N__64781),
            .I(\c0.n19554 ));
    Odrv4 I__15437 (
            .O(N__64776),
            .I(\c0.n19554 ));
    InMux I__15436 (
            .O(N__64771),
            .I(N__64764));
    InMux I__15435 (
            .O(N__64770),
            .I(N__64764));
    InMux I__15434 (
            .O(N__64769),
            .I(N__64761));
    LocalMux I__15433 (
            .O(N__64764),
            .I(N__64757));
    LocalMux I__15432 (
            .O(N__64761),
            .I(N__64754));
    CascadeMux I__15431 (
            .O(N__64760),
            .I(N__64751));
    Span4Mux_v I__15430 (
            .O(N__64757),
            .I(N__64748));
    Span4Mux_v I__15429 (
            .O(N__64754),
            .I(N__64745));
    InMux I__15428 (
            .O(N__64751),
            .I(N__64742));
    Span4Mux_v I__15427 (
            .O(N__64748),
            .I(N__64739));
    Span4Mux_v I__15426 (
            .O(N__64745),
            .I(N__64736));
    LocalMux I__15425 (
            .O(N__64742),
            .I(N__64731));
    Span4Mux_h I__15424 (
            .O(N__64739),
            .I(N__64731));
    Span4Mux_v I__15423 (
            .O(N__64736),
            .I(N__64728));
    Odrv4 I__15422 (
            .O(N__64731),
            .I(\c0.data_in_frame_17_4 ));
    Odrv4 I__15421 (
            .O(N__64728),
            .I(\c0.data_in_frame_17_4 ));
    CascadeMux I__15420 (
            .O(N__64723),
            .I(N__64720));
    InMux I__15419 (
            .O(N__64720),
            .I(N__64717));
    LocalMux I__15418 (
            .O(N__64717),
            .I(N__64714));
    Sp12to4 I__15417 (
            .O(N__64714),
            .I(N__64711));
    Odrv12 I__15416 (
            .O(N__64711),
            .I(\c0.n18_adj_3235 ));
    CascadeMux I__15415 (
            .O(N__64708),
            .I(N__64704));
    InMux I__15414 (
            .O(N__64707),
            .I(N__64700));
    InMux I__15413 (
            .O(N__64704),
            .I(N__64696));
    InMux I__15412 (
            .O(N__64703),
            .I(N__64693));
    LocalMux I__15411 (
            .O(N__64700),
            .I(N__64690));
    InMux I__15410 (
            .O(N__64699),
            .I(N__64687));
    LocalMux I__15409 (
            .O(N__64696),
            .I(N__64684));
    LocalMux I__15408 (
            .O(N__64693),
            .I(N__64680));
    Span4Mux_v I__15407 (
            .O(N__64690),
            .I(N__64675));
    LocalMux I__15406 (
            .O(N__64687),
            .I(N__64675));
    Span4Mux_h I__15405 (
            .O(N__64684),
            .I(N__64672));
    CascadeMux I__15404 (
            .O(N__64683),
            .I(N__64669));
    Span4Mux_v I__15403 (
            .O(N__64680),
            .I(N__64666));
    Span4Mux_v I__15402 (
            .O(N__64675),
            .I(N__64661));
    Span4Mux_v I__15401 (
            .O(N__64672),
            .I(N__64661));
    InMux I__15400 (
            .O(N__64669),
            .I(N__64658));
    Span4Mux_v I__15399 (
            .O(N__64666),
            .I(N__64655));
    Span4Mux_v I__15398 (
            .O(N__64661),
            .I(N__64652));
    LocalMux I__15397 (
            .O(N__64658),
            .I(\c0.data_in_frame_15_3 ));
    Odrv4 I__15396 (
            .O(N__64655),
            .I(\c0.data_in_frame_15_3 ));
    Odrv4 I__15395 (
            .O(N__64652),
            .I(\c0.data_in_frame_15_3 ));
    InMux I__15394 (
            .O(N__64645),
            .I(N__64642));
    LocalMux I__15393 (
            .O(N__64642),
            .I(N__64639));
    Span4Mux_v I__15392 (
            .O(N__64639),
            .I(N__64636));
    Odrv4 I__15391 (
            .O(N__64636),
            .I(\c0.n10_adj_3483 ));
    InMux I__15390 (
            .O(N__64633),
            .I(N__64629));
    InMux I__15389 (
            .O(N__64632),
            .I(N__64625));
    LocalMux I__15388 (
            .O(N__64629),
            .I(N__64620));
    InMux I__15387 (
            .O(N__64628),
            .I(N__64617));
    LocalMux I__15386 (
            .O(N__64625),
            .I(N__64614));
    InMux I__15385 (
            .O(N__64624),
            .I(N__64609));
    InMux I__15384 (
            .O(N__64623),
            .I(N__64609));
    Span4Mux_v I__15383 (
            .O(N__64620),
            .I(N__64603));
    LocalMux I__15382 (
            .O(N__64617),
            .I(N__64603));
    Span4Mux_v I__15381 (
            .O(N__64614),
            .I(N__64598));
    LocalMux I__15380 (
            .O(N__64609),
            .I(N__64598));
    InMux I__15379 (
            .O(N__64608),
            .I(N__64595));
    Span4Mux_h I__15378 (
            .O(N__64603),
            .I(N__64590));
    Span4Mux_v I__15377 (
            .O(N__64598),
            .I(N__64590));
    LocalMux I__15376 (
            .O(N__64595),
            .I(\c0.n18420 ));
    Odrv4 I__15375 (
            .O(N__64590),
            .I(\c0.n18420 ));
    InMux I__15374 (
            .O(N__64585),
            .I(N__64579));
    InMux I__15373 (
            .O(N__64584),
            .I(N__64574));
    InMux I__15372 (
            .O(N__64583),
            .I(N__64569));
    InMux I__15371 (
            .O(N__64582),
            .I(N__64569));
    LocalMux I__15370 (
            .O(N__64579),
            .I(N__64566));
    CascadeMux I__15369 (
            .O(N__64578),
            .I(N__64561));
    InMux I__15368 (
            .O(N__64577),
            .I(N__64558));
    LocalMux I__15367 (
            .O(N__64574),
            .I(N__64555));
    LocalMux I__15366 (
            .O(N__64569),
            .I(N__64552));
    Span4Mux_v I__15365 (
            .O(N__64566),
            .I(N__64543));
    InMux I__15364 (
            .O(N__64565),
            .I(N__64535));
    InMux I__15363 (
            .O(N__64564),
            .I(N__64535));
    InMux I__15362 (
            .O(N__64561),
            .I(N__64535));
    LocalMux I__15361 (
            .O(N__64558),
            .I(N__64530));
    Span4Mux_v I__15360 (
            .O(N__64555),
            .I(N__64530));
    Span4Mux_v I__15359 (
            .O(N__64552),
            .I(N__64527));
    InMux I__15358 (
            .O(N__64551),
            .I(N__64524));
    InMux I__15357 (
            .O(N__64550),
            .I(N__64519));
    InMux I__15356 (
            .O(N__64549),
            .I(N__64519));
    InMux I__15355 (
            .O(N__64548),
            .I(N__64512));
    InMux I__15354 (
            .O(N__64547),
            .I(N__64512));
    InMux I__15353 (
            .O(N__64546),
            .I(N__64512));
    Span4Mux_h I__15352 (
            .O(N__64543),
            .I(N__64509));
    InMux I__15351 (
            .O(N__64542),
            .I(N__64506));
    LocalMux I__15350 (
            .O(N__64535),
            .I(N__64503));
    Span4Mux_v I__15349 (
            .O(N__64530),
            .I(N__64499));
    Span4Mux_v I__15348 (
            .O(N__64527),
            .I(N__64496));
    LocalMux I__15347 (
            .O(N__64524),
            .I(N__64493));
    LocalMux I__15346 (
            .O(N__64519),
            .I(N__64486));
    LocalMux I__15345 (
            .O(N__64512),
            .I(N__64486));
    Span4Mux_h I__15344 (
            .O(N__64509),
            .I(N__64486));
    LocalMux I__15343 (
            .O(N__64506),
            .I(N__64481));
    Span12Mux_h I__15342 (
            .O(N__64503),
            .I(N__64481));
    InMux I__15341 (
            .O(N__64502),
            .I(N__64478));
    Span4Mux_h I__15340 (
            .O(N__64499),
            .I(N__64475));
    Span4Mux_v I__15339 (
            .O(N__64496),
            .I(N__64472));
    Span4Mux_h I__15338 (
            .O(N__64493),
            .I(N__64467));
    Span4Mux_v I__15337 (
            .O(N__64486),
            .I(N__64467));
    Span12Mux_v I__15336 (
            .O(N__64481),
            .I(N__64464));
    LocalMux I__15335 (
            .O(N__64478),
            .I(\c0.n19131 ));
    Odrv4 I__15334 (
            .O(N__64475),
            .I(\c0.n19131 ));
    Odrv4 I__15333 (
            .O(N__64472),
            .I(\c0.n19131 ));
    Odrv4 I__15332 (
            .O(N__64467),
            .I(\c0.n19131 ));
    Odrv12 I__15331 (
            .O(N__64464),
            .I(\c0.n19131 ));
    CascadeMux I__15330 (
            .O(N__64453),
            .I(N__64450));
    InMux I__15329 (
            .O(N__64450),
            .I(N__64446));
    InMux I__15328 (
            .O(N__64449),
            .I(N__64443));
    LocalMux I__15327 (
            .O(N__64446),
            .I(N__64439));
    LocalMux I__15326 (
            .O(N__64443),
            .I(N__64435));
    InMux I__15325 (
            .O(N__64442),
            .I(N__64432));
    Span12Mux_h I__15324 (
            .O(N__64439),
            .I(N__64429));
    InMux I__15323 (
            .O(N__64438),
            .I(N__64426));
    Span4Mux_h I__15322 (
            .O(N__64435),
            .I(N__64423));
    LocalMux I__15321 (
            .O(N__64432),
            .I(\c0.data_in_frame_11_7 ));
    Odrv12 I__15320 (
            .O(N__64429),
            .I(\c0.data_in_frame_11_7 ));
    LocalMux I__15319 (
            .O(N__64426),
            .I(\c0.data_in_frame_11_7 ));
    Odrv4 I__15318 (
            .O(N__64423),
            .I(\c0.data_in_frame_11_7 ));
    InMux I__15317 (
            .O(N__64414),
            .I(N__64406));
    InMux I__15316 (
            .O(N__64413),
            .I(N__64401));
    InMux I__15315 (
            .O(N__64412),
            .I(N__64401));
    InMux I__15314 (
            .O(N__64411),
            .I(N__64398));
    InMux I__15313 (
            .O(N__64410),
            .I(N__64394));
    InMux I__15312 (
            .O(N__64409),
            .I(N__64390));
    LocalMux I__15311 (
            .O(N__64406),
            .I(N__64379));
    LocalMux I__15310 (
            .O(N__64401),
            .I(N__64379));
    LocalMux I__15309 (
            .O(N__64398),
            .I(N__64379));
    InMux I__15308 (
            .O(N__64397),
            .I(N__64376));
    LocalMux I__15307 (
            .O(N__64394),
            .I(N__64373));
    InMux I__15306 (
            .O(N__64393),
            .I(N__64370));
    LocalMux I__15305 (
            .O(N__64390),
            .I(N__64367));
    CascadeMux I__15304 (
            .O(N__64389),
            .I(N__64363));
    InMux I__15303 (
            .O(N__64388),
            .I(N__64355));
    InMux I__15302 (
            .O(N__64387),
            .I(N__64355));
    InMux I__15301 (
            .O(N__64386),
            .I(N__64355));
    Span4Mux_h I__15300 (
            .O(N__64379),
            .I(N__64352));
    LocalMux I__15299 (
            .O(N__64376),
            .I(N__64349));
    Span4Mux_v I__15298 (
            .O(N__64373),
            .I(N__64346));
    LocalMux I__15297 (
            .O(N__64370),
            .I(N__64341));
    Span4Mux_v I__15296 (
            .O(N__64367),
            .I(N__64337));
    InMux I__15295 (
            .O(N__64366),
            .I(N__64330));
    InMux I__15294 (
            .O(N__64363),
            .I(N__64330));
    InMux I__15293 (
            .O(N__64362),
            .I(N__64330));
    LocalMux I__15292 (
            .O(N__64355),
            .I(N__64327));
    Span4Mux_v I__15291 (
            .O(N__64352),
            .I(N__64322));
    Span4Mux_v I__15290 (
            .O(N__64349),
            .I(N__64322));
    Span4Mux_h I__15289 (
            .O(N__64346),
            .I(N__64319));
    InMux I__15288 (
            .O(N__64345),
            .I(N__64314));
    InMux I__15287 (
            .O(N__64344),
            .I(N__64314));
    Span4Mux_v I__15286 (
            .O(N__64341),
            .I(N__64311));
    InMux I__15285 (
            .O(N__64340),
            .I(N__64308));
    Span4Mux_h I__15284 (
            .O(N__64337),
            .I(N__64305));
    LocalMux I__15283 (
            .O(N__64330),
            .I(N__64302));
    Sp12to4 I__15282 (
            .O(N__64327),
            .I(N__64299));
    Sp12to4 I__15281 (
            .O(N__64322),
            .I(N__64296));
    Sp12to4 I__15280 (
            .O(N__64319),
            .I(N__64293));
    LocalMux I__15279 (
            .O(N__64314),
            .I(N__64290));
    Sp12to4 I__15278 (
            .O(N__64311),
            .I(N__64287));
    LocalMux I__15277 (
            .O(N__64308),
            .I(N__64284));
    Span4Mux_v I__15276 (
            .O(N__64305),
            .I(N__64279));
    Span4Mux_v I__15275 (
            .O(N__64302),
            .I(N__64279));
    Span12Mux_v I__15274 (
            .O(N__64299),
            .I(N__64272));
    Span12Mux_v I__15273 (
            .O(N__64296),
            .I(N__64272));
    Span12Mux_v I__15272 (
            .O(N__64293),
            .I(N__64272));
    Span12Mux_s8_v I__15271 (
            .O(N__64290),
            .I(N__64267));
    Span12Mux_h I__15270 (
            .O(N__64287),
            .I(N__64267));
    Span4Mux_v I__15269 (
            .O(N__64284),
            .I(N__64264));
    Odrv4 I__15268 (
            .O(N__64279),
            .I(\c0.n15489 ));
    Odrv12 I__15267 (
            .O(N__64272),
            .I(\c0.n15489 ));
    Odrv12 I__15266 (
            .O(N__64267),
            .I(\c0.n15489 ));
    Odrv4 I__15265 (
            .O(N__64264),
            .I(\c0.n15489 ));
    InMux I__15264 (
            .O(N__64255),
            .I(N__64239));
    InMux I__15263 (
            .O(N__64254),
            .I(N__64228));
    InMux I__15262 (
            .O(N__64253),
            .I(N__64228));
    InMux I__15261 (
            .O(N__64252),
            .I(N__64228));
    InMux I__15260 (
            .O(N__64251),
            .I(N__64228));
    InMux I__15259 (
            .O(N__64250),
            .I(N__64225));
    CascadeMux I__15258 (
            .O(N__64249),
            .I(N__64222));
    InMux I__15257 (
            .O(N__64248),
            .I(N__64217));
    InMux I__15256 (
            .O(N__64247),
            .I(N__64210));
    InMux I__15255 (
            .O(N__64246),
            .I(N__64210));
    InMux I__15254 (
            .O(N__64245),
            .I(N__64210));
    InMux I__15253 (
            .O(N__64244),
            .I(N__64203));
    InMux I__15252 (
            .O(N__64243),
            .I(N__64203));
    InMux I__15251 (
            .O(N__64242),
            .I(N__64203));
    LocalMux I__15250 (
            .O(N__64239),
            .I(N__64200));
    InMux I__15249 (
            .O(N__64238),
            .I(N__64193));
    InMux I__15248 (
            .O(N__64237),
            .I(N__64193));
    LocalMux I__15247 (
            .O(N__64228),
            .I(N__64188));
    LocalMux I__15246 (
            .O(N__64225),
            .I(N__64188));
    InMux I__15245 (
            .O(N__64222),
            .I(N__64185));
    InMux I__15244 (
            .O(N__64221),
            .I(N__64180));
    InMux I__15243 (
            .O(N__64220),
            .I(N__64177));
    LocalMux I__15242 (
            .O(N__64217),
            .I(N__64174));
    LocalMux I__15241 (
            .O(N__64210),
            .I(N__64167));
    LocalMux I__15240 (
            .O(N__64203),
            .I(N__64167));
    Span4Mux_v I__15239 (
            .O(N__64200),
            .I(N__64167));
    InMux I__15238 (
            .O(N__64199),
            .I(N__64164));
    InMux I__15237 (
            .O(N__64198),
            .I(N__64161));
    LocalMux I__15236 (
            .O(N__64193),
            .I(N__64158));
    Span4Mux_v I__15235 (
            .O(N__64188),
            .I(N__64153));
    LocalMux I__15234 (
            .O(N__64185),
            .I(N__64153));
    InMux I__15233 (
            .O(N__64184),
            .I(N__64148));
    InMux I__15232 (
            .O(N__64183),
            .I(N__64148));
    LocalMux I__15231 (
            .O(N__64180),
            .I(N__64145));
    LocalMux I__15230 (
            .O(N__64177),
            .I(N__64140));
    Span4Mux_v I__15229 (
            .O(N__64174),
            .I(N__64140));
    Span4Mux_v I__15228 (
            .O(N__64167),
            .I(N__64137));
    LocalMux I__15227 (
            .O(N__64164),
            .I(N__64133));
    LocalMux I__15226 (
            .O(N__64161),
            .I(N__64130));
    Span4Mux_v I__15225 (
            .O(N__64158),
            .I(N__64127));
    Span4Mux_h I__15224 (
            .O(N__64153),
            .I(N__64124));
    LocalMux I__15223 (
            .O(N__64148),
            .I(N__64121));
    Span4Mux_h I__15222 (
            .O(N__64145),
            .I(N__64114));
    Span4Mux_v I__15221 (
            .O(N__64140),
            .I(N__64114));
    Span4Mux_h I__15220 (
            .O(N__64137),
            .I(N__64114));
    InMux I__15219 (
            .O(N__64136),
            .I(N__64110));
    Span4Mux_v I__15218 (
            .O(N__64133),
            .I(N__64107));
    Span4Mux_h I__15217 (
            .O(N__64130),
            .I(N__64104));
    Span4Mux_h I__15216 (
            .O(N__64127),
            .I(N__64101));
    Sp12to4 I__15215 (
            .O(N__64124),
            .I(N__64096));
    Span12Mux_s10_v I__15214 (
            .O(N__64121),
            .I(N__64096));
    Span4Mux_v I__15213 (
            .O(N__64114),
            .I(N__64093));
    InMux I__15212 (
            .O(N__64113),
            .I(N__64090));
    LocalMux I__15211 (
            .O(N__64110),
            .I(N__64087));
    Span4Mux_h I__15210 (
            .O(N__64107),
            .I(N__64084));
    Sp12to4 I__15209 (
            .O(N__64104),
            .I(N__64081));
    Span4Mux_v I__15208 (
            .O(N__64101),
            .I(N__64078));
    Span12Mux_v I__15207 (
            .O(N__64096),
            .I(N__64075));
    Span4Mux_v I__15206 (
            .O(N__64093),
            .I(N__64072));
    LocalMux I__15205 (
            .O(N__64090),
            .I(\c0.n19140 ));
    Odrv12 I__15204 (
            .O(N__64087),
            .I(\c0.n19140 ));
    Odrv4 I__15203 (
            .O(N__64084),
            .I(\c0.n19140 ));
    Odrv12 I__15202 (
            .O(N__64081),
            .I(\c0.n19140 ));
    Odrv4 I__15201 (
            .O(N__64078),
            .I(\c0.n19140 ));
    Odrv12 I__15200 (
            .O(N__64075),
            .I(\c0.n19140 ));
    Odrv4 I__15199 (
            .O(N__64072),
            .I(\c0.n19140 ));
    InMux I__15198 (
            .O(N__64057),
            .I(N__64053));
    InMux I__15197 (
            .O(N__64056),
            .I(N__64050));
    LocalMux I__15196 (
            .O(N__64053),
            .I(N__64046));
    LocalMux I__15195 (
            .O(N__64050),
            .I(N__64043));
    CascadeMux I__15194 (
            .O(N__64049),
            .I(N__64040));
    Span4Mux_v I__15193 (
            .O(N__64046),
            .I(N__64036));
    Span4Mux_h I__15192 (
            .O(N__64043),
            .I(N__64033));
    InMux I__15191 (
            .O(N__64040),
            .I(N__64028));
    InMux I__15190 (
            .O(N__64039),
            .I(N__64028));
    Odrv4 I__15189 (
            .O(N__64036),
            .I(\c0.data_in_frame_15_5 ));
    Odrv4 I__15188 (
            .O(N__64033),
            .I(\c0.data_in_frame_15_5 ));
    LocalMux I__15187 (
            .O(N__64028),
            .I(\c0.data_in_frame_15_5 ));
    CascadeMux I__15186 (
            .O(N__64021),
            .I(\c0.n9_adj_3552_cascade_ ));
    CascadeMux I__15185 (
            .O(N__64018),
            .I(N__64015));
    InMux I__15184 (
            .O(N__64015),
            .I(N__64010));
    CascadeMux I__15183 (
            .O(N__64014),
            .I(N__64007));
    InMux I__15182 (
            .O(N__64013),
            .I(N__64004));
    LocalMux I__15181 (
            .O(N__64010),
            .I(N__63999));
    InMux I__15180 (
            .O(N__64007),
            .I(N__63996));
    LocalMux I__15179 (
            .O(N__64004),
            .I(N__63991));
    InMux I__15178 (
            .O(N__64003),
            .I(N__63988));
    InMux I__15177 (
            .O(N__64002),
            .I(N__63985));
    Span4Mux_v I__15176 (
            .O(N__63999),
            .I(N__63982));
    LocalMux I__15175 (
            .O(N__63996),
            .I(N__63979));
    InMux I__15174 (
            .O(N__63995),
            .I(N__63974));
    InMux I__15173 (
            .O(N__63994),
            .I(N__63974));
    Span12Mux_h I__15172 (
            .O(N__63991),
            .I(N__63971));
    LocalMux I__15171 (
            .O(N__63988),
            .I(N__63968));
    LocalMux I__15170 (
            .O(N__63985),
            .I(data_in_frame_18_3));
    Odrv4 I__15169 (
            .O(N__63982),
            .I(data_in_frame_18_3));
    Odrv4 I__15168 (
            .O(N__63979),
            .I(data_in_frame_18_3));
    LocalMux I__15167 (
            .O(N__63974),
            .I(data_in_frame_18_3));
    Odrv12 I__15166 (
            .O(N__63971),
            .I(data_in_frame_18_3));
    Odrv4 I__15165 (
            .O(N__63968),
            .I(data_in_frame_18_3));
    InMux I__15164 (
            .O(N__63955),
            .I(N__63952));
    LocalMux I__15163 (
            .O(N__63952),
            .I(N__63949));
    Span4Mux_v I__15162 (
            .O(N__63949),
            .I(N__63945));
    InMux I__15161 (
            .O(N__63948),
            .I(N__63940));
    Span4Mux_h I__15160 (
            .O(N__63945),
            .I(N__63934));
    InMux I__15159 (
            .O(N__63944),
            .I(N__63931));
    InMux I__15158 (
            .O(N__63943),
            .I(N__63928));
    LocalMux I__15157 (
            .O(N__63940),
            .I(N__63925));
    InMux I__15156 (
            .O(N__63939),
            .I(N__63922));
    InMux I__15155 (
            .O(N__63938),
            .I(N__63919));
    InMux I__15154 (
            .O(N__63937),
            .I(N__63916));
    Span4Mux_h I__15153 (
            .O(N__63934),
            .I(N__63910));
    LocalMux I__15152 (
            .O(N__63931),
            .I(N__63910));
    LocalMux I__15151 (
            .O(N__63928),
            .I(N__63907));
    Span4Mux_h I__15150 (
            .O(N__63925),
            .I(N__63900));
    LocalMux I__15149 (
            .O(N__63922),
            .I(N__63900));
    LocalMux I__15148 (
            .O(N__63919),
            .I(N__63900));
    LocalMux I__15147 (
            .O(N__63916),
            .I(N__63897));
    InMux I__15146 (
            .O(N__63915),
            .I(N__63894));
    Span4Mux_v I__15145 (
            .O(N__63910),
            .I(N__63891));
    Span4Mux_h I__15144 (
            .O(N__63907),
            .I(N__63888));
    Span4Mux_v I__15143 (
            .O(N__63900),
            .I(N__63885));
    Span4Mux_v I__15142 (
            .O(N__63897),
            .I(N__63880));
    LocalMux I__15141 (
            .O(N__63894),
            .I(N__63880));
    Odrv4 I__15140 (
            .O(N__63891),
            .I(n19129));
    Odrv4 I__15139 (
            .O(N__63888),
            .I(n19129));
    Odrv4 I__15138 (
            .O(N__63885),
            .I(n19129));
    Odrv4 I__15137 (
            .O(N__63880),
            .I(n19129));
    InMux I__15136 (
            .O(N__63871),
            .I(N__63865));
    InMux I__15135 (
            .O(N__63870),
            .I(N__63865));
    LocalMux I__15134 (
            .O(N__63865),
            .I(data_in_frame_18_4));
    InMux I__15133 (
            .O(N__63862),
            .I(N__63858));
    InMux I__15132 (
            .O(N__63861),
            .I(N__63855));
    LocalMux I__15131 (
            .O(N__63858),
            .I(N__63850));
    LocalMux I__15130 (
            .O(N__63855),
            .I(N__63847));
    InMux I__15129 (
            .O(N__63854),
            .I(N__63844));
    CascadeMux I__15128 (
            .O(N__63853),
            .I(N__63840));
    Span4Mux_v I__15127 (
            .O(N__63850),
            .I(N__63837));
    Span4Mux_h I__15126 (
            .O(N__63847),
            .I(N__63834));
    LocalMux I__15125 (
            .O(N__63844),
            .I(N__63831));
    InMux I__15124 (
            .O(N__63843),
            .I(N__63828));
    InMux I__15123 (
            .O(N__63840),
            .I(N__63825));
    Span4Mux_v I__15122 (
            .O(N__63837),
            .I(N__63822));
    Span4Mux_h I__15121 (
            .O(N__63834),
            .I(N__63819));
    Span12Mux_h I__15120 (
            .O(N__63831),
            .I(N__63814));
    LocalMux I__15119 (
            .O(N__63828),
            .I(N__63814));
    LocalMux I__15118 (
            .O(N__63825),
            .I(\c0.data_in_frame_12_1 ));
    Odrv4 I__15117 (
            .O(N__63822),
            .I(\c0.data_in_frame_12_1 ));
    Odrv4 I__15116 (
            .O(N__63819),
            .I(\c0.data_in_frame_12_1 ));
    Odrv12 I__15115 (
            .O(N__63814),
            .I(\c0.data_in_frame_12_1 ));
    InMux I__15114 (
            .O(N__63805),
            .I(N__63802));
    LocalMux I__15113 (
            .O(N__63802),
            .I(\c0.n7_adj_3000 ));
    CascadeMux I__15112 (
            .O(N__63799),
            .I(N__63796));
    InMux I__15111 (
            .O(N__63796),
            .I(N__63791));
    InMux I__15110 (
            .O(N__63795),
            .I(N__63786));
    InMux I__15109 (
            .O(N__63794),
            .I(N__63786));
    LocalMux I__15108 (
            .O(N__63791),
            .I(\c0.n19430 ));
    LocalMux I__15107 (
            .O(N__63786),
            .I(\c0.n19430 ));
    CascadeMux I__15106 (
            .O(N__63781),
            .I(\c0.n7_adj_3000_cascade_ ));
    InMux I__15105 (
            .O(N__63778),
            .I(N__63771));
    CascadeMux I__15104 (
            .O(N__63777),
            .I(N__63768));
    InMux I__15103 (
            .O(N__63776),
            .I(N__63762));
    InMux I__15102 (
            .O(N__63775),
            .I(N__63759));
    InMux I__15101 (
            .O(N__63774),
            .I(N__63756));
    LocalMux I__15100 (
            .O(N__63771),
            .I(N__63753));
    InMux I__15099 (
            .O(N__63768),
            .I(N__63748));
    InMux I__15098 (
            .O(N__63767),
            .I(N__63748));
    InMux I__15097 (
            .O(N__63766),
            .I(N__63743));
    InMux I__15096 (
            .O(N__63765),
            .I(N__63743));
    LocalMux I__15095 (
            .O(N__63762),
            .I(N__63736));
    LocalMux I__15094 (
            .O(N__63759),
            .I(N__63736));
    LocalMux I__15093 (
            .O(N__63756),
            .I(N__63733));
    Span4Mux_h I__15092 (
            .O(N__63753),
            .I(N__63728));
    LocalMux I__15091 (
            .O(N__63748),
            .I(N__63728));
    LocalMux I__15090 (
            .O(N__63743),
            .I(N__63725));
    InMux I__15089 (
            .O(N__63742),
            .I(N__63720));
    InMux I__15088 (
            .O(N__63741),
            .I(N__63720));
    Sp12to4 I__15087 (
            .O(N__63736),
            .I(N__63715));
    Span12Mux_h I__15086 (
            .O(N__63733),
            .I(N__63715));
    Span4Mux_h I__15085 (
            .O(N__63728),
            .I(N__63712));
    Span12Mux_v I__15084 (
            .O(N__63725),
            .I(N__63709));
    LocalMux I__15083 (
            .O(N__63720),
            .I(data_in_frame_16_3));
    Odrv12 I__15082 (
            .O(N__63715),
            .I(data_in_frame_16_3));
    Odrv4 I__15081 (
            .O(N__63712),
            .I(data_in_frame_16_3));
    Odrv12 I__15080 (
            .O(N__63709),
            .I(data_in_frame_16_3));
    CascadeMux I__15079 (
            .O(N__63700),
            .I(N__63697));
    InMux I__15078 (
            .O(N__63697),
            .I(N__63694));
    LocalMux I__15077 (
            .O(N__63694),
            .I(N__63691));
    Odrv4 I__15076 (
            .O(N__63691),
            .I(\c0.n6 ));
    CascadeMux I__15075 (
            .O(N__63688),
            .I(N__63684));
    InMux I__15074 (
            .O(N__63687),
            .I(N__63680));
    InMux I__15073 (
            .O(N__63684),
            .I(N__63673));
    InMux I__15072 (
            .O(N__63683),
            .I(N__63673));
    LocalMux I__15071 (
            .O(N__63680),
            .I(N__63670));
    InMux I__15070 (
            .O(N__63679),
            .I(N__63665));
    InMux I__15069 (
            .O(N__63678),
            .I(N__63665));
    LocalMux I__15068 (
            .O(N__63673),
            .I(N__63658));
    Span4Mux_v I__15067 (
            .O(N__63670),
            .I(N__63658));
    LocalMux I__15066 (
            .O(N__63665),
            .I(N__63658));
    Span4Mux_h I__15065 (
            .O(N__63658),
            .I(N__63655));
    Odrv4 I__15064 (
            .O(N__63655),
            .I(\c0.n19187 ));
    CascadeMux I__15063 (
            .O(N__63652),
            .I(N__63648));
    InMux I__15062 (
            .O(N__63651),
            .I(N__63643));
    InMux I__15061 (
            .O(N__63648),
            .I(N__63640));
    InMux I__15060 (
            .O(N__63647),
            .I(N__63637));
    InMux I__15059 (
            .O(N__63646),
            .I(N__63634));
    LocalMux I__15058 (
            .O(N__63643),
            .I(N__63631));
    LocalMux I__15057 (
            .O(N__63640),
            .I(N__63622));
    LocalMux I__15056 (
            .O(N__63637),
            .I(N__63622));
    LocalMux I__15055 (
            .O(N__63634),
            .I(N__63619));
    Span4Mux_v I__15054 (
            .O(N__63631),
            .I(N__63616));
    InMux I__15053 (
            .O(N__63630),
            .I(N__63611));
    InMux I__15052 (
            .O(N__63629),
            .I(N__63611));
    InMux I__15051 (
            .O(N__63628),
            .I(N__63608));
    InMux I__15050 (
            .O(N__63627),
            .I(N__63605));
    Span4Mux_v I__15049 (
            .O(N__63622),
            .I(N__63602));
    Span4Mux_v I__15048 (
            .O(N__63619),
            .I(N__63597));
    Span4Mux_h I__15047 (
            .O(N__63616),
            .I(N__63597));
    LocalMux I__15046 (
            .O(N__63611),
            .I(N__63590));
    LocalMux I__15045 (
            .O(N__63608),
            .I(N__63590));
    LocalMux I__15044 (
            .O(N__63605),
            .I(N__63590));
    Odrv4 I__15043 (
            .O(N__63602),
            .I(\c0.n46_adj_3443 ));
    Odrv4 I__15042 (
            .O(N__63597),
            .I(\c0.n46_adj_3443 ));
    Odrv12 I__15041 (
            .O(N__63590),
            .I(\c0.n46_adj_3443 ));
    CascadeMux I__15040 (
            .O(N__63583),
            .I(N__63580));
    InMux I__15039 (
            .O(N__63580),
            .I(N__63577));
    LocalMux I__15038 (
            .O(N__63577),
            .I(N__63570));
    InMux I__15037 (
            .O(N__63576),
            .I(N__63567));
    CascadeMux I__15036 (
            .O(N__63575),
            .I(N__63564));
    InMux I__15035 (
            .O(N__63574),
            .I(N__63561));
    CascadeMux I__15034 (
            .O(N__63573),
            .I(N__63557));
    Span4Mux_v I__15033 (
            .O(N__63570),
            .I(N__63552));
    LocalMux I__15032 (
            .O(N__63567),
            .I(N__63552));
    InMux I__15031 (
            .O(N__63564),
            .I(N__63549));
    LocalMux I__15030 (
            .O(N__63561),
            .I(N__63546));
    InMux I__15029 (
            .O(N__63560),
            .I(N__63543));
    InMux I__15028 (
            .O(N__63557),
            .I(N__63540));
    Span4Mux_v I__15027 (
            .O(N__63552),
            .I(N__63535));
    LocalMux I__15026 (
            .O(N__63549),
            .I(N__63535));
    Span4Mux_v I__15025 (
            .O(N__63546),
            .I(N__63529));
    LocalMux I__15024 (
            .O(N__63543),
            .I(N__63529));
    LocalMux I__15023 (
            .O(N__63540),
            .I(N__63526));
    Span4Mux_h I__15022 (
            .O(N__63535),
            .I(N__63523));
    CascadeMux I__15021 (
            .O(N__63534),
            .I(N__63520));
    Sp12to4 I__15020 (
            .O(N__63529),
            .I(N__63517));
    Span4Mux_h I__15019 (
            .O(N__63526),
            .I(N__63512));
    Span4Mux_h I__15018 (
            .O(N__63523),
            .I(N__63512));
    InMux I__15017 (
            .O(N__63520),
            .I(N__63509));
    Span12Mux_h I__15016 (
            .O(N__63517),
            .I(N__63506));
    Span4Mux_v I__15015 (
            .O(N__63512),
            .I(N__63503));
    LocalMux I__15014 (
            .O(N__63509),
            .I(\c0.data_in_frame_15_0 ));
    Odrv12 I__15013 (
            .O(N__63506),
            .I(\c0.data_in_frame_15_0 ));
    Odrv4 I__15012 (
            .O(N__63503),
            .I(\c0.data_in_frame_15_0 ));
    InMux I__15011 (
            .O(N__63496),
            .I(N__63489));
    InMux I__15010 (
            .O(N__63495),
            .I(N__63489));
    InMux I__15009 (
            .O(N__63494),
            .I(N__63486));
    LocalMux I__15008 (
            .O(N__63489),
            .I(N__63482));
    LocalMux I__15007 (
            .O(N__63486),
            .I(N__63479));
    InMux I__15006 (
            .O(N__63485),
            .I(N__63476));
    Span4Mux_v I__15005 (
            .O(N__63482),
            .I(N__63473));
    Span4Mux_v I__15004 (
            .O(N__63479),
            .I(N__63468));
    LocalMux I__15003 (
            .O(N__63476),
            .I(N__63468));
    Sp12to4 I__15002 (
            .O(N__63473),
            .I(N__63465));
    Span4Mux_h I__15001 (
            .O(N__63468),
            .I(N__63462));
    Odrv12 I__15000 (
            .O(N__63465),
            .I(\c0.n40_adj_3413 ));
    Odrv4 I__14999 (
            .O(N__63462),
            .I(\c0.n40_adj_3413 ));
    CascadeMux I__14998 (
            .O(N__63457),
            .I(N__63452));
    CascadeMux I__14997 (
            .O(N__63456),
            .I(N__63449));
    InMux I__14996 (
            .O(N__63455),
            .I(N__63446));
    InMux I__14995 (
            .O(N__63452),
            .I(N__63441));
    InMux I__14994 (
            .O(N__63449),
            .I(N__63441));
    LocalMux I__14993 (
            .O(N__63446),
            .I(N__63438));
    LocalMux I__14992 (
            .O(N__63441),
            .I(N__63435));
    Sp12to4 I__14991 (
            .O(N__63438),
            .I(N__63432));
    Span4Mux_h I__14990 (
            .O(N__63435),
            .I(N__63429));
    Span12Mux_v I__14989 (
            .O(N__63432),
            .I(N__63426));
    Span4Mux_v I__14988 (
            .O(N__63429),
            .I(N__63423));
    Odrv12 I__14987 (
            .O(N__63426),
            .I(\c0.n45_adj_3138 ));
    Odrv4 I__14986 (
            .O(N__63423),
            .I(\c0.n45_adj_3138 ));
    InMux I__14985 (
            .O(N__63418),
            .I(N__63409));
    InMux I__14984 (
            .O(N__63417),
            .I(N__63404));
    InMux I__14983 (
            .O(N__63416),
            .I(N__63404));
    InMux I__14982 (
            .O(N__63415),
            .I(N__63399));
    InMux I__14981 (
            .O(N__63414),
            .I(N__63399));
    InMux I__14980 (
            .O(N__63413),
            .I(N__63396));
    InMux I__14979 (
            .O(N__63412),
            .I(N__63391));
    LocalMux I__14978 (
            .O(N__63409),
            .I(N__63386));
    LocalMux I__14977 (
            .O(N__63404),
            .I(N__63381));
    LocalMux I__14976 (
            .O(N__63399),
            .I(N__63381));
    LocalMux I__14975 (
            .O(N__63396),
            .I(N__63374));
    InMux I__14974 (
            .O(N__63395),
            .I(N__63371));
    InMux I__14973 (
            .O(N__63394),
            .I(N__63368));
    LocalMux I__14972 (
            .O(N__63391),
            .I(N__63365));
    CascadeMux I__14971 (
            .O(N__63390),
            .I(N__63362));
    CascadeMux I__14970 (
            .O(N__63389),
            .I(N__63359));
    Span4Mux_v I__14969 (
            .O(N__63386),
            .I(N__63348));
    Span4Mux_v I__14968 (
            .O(N__63381),
            .I(N__63348));
    InMux I__14967 (
            .O(N__63380),
            .I(N__63343));
    InMux I__14966 (
            .O(N__63379),
            .I(N__63343));
    InMux I__14965 (
            .O(N__63378),
            .I(N__63340));
    InMux I__14964 (
            .O(N__63377),
            .I(N__63337));
    Span4Mux_h I__14963 (
            .O(N__63374),
            .I(N__63334));
    LocalMux I__14962 (
            .O(N__63371),
            .I(N__63331));
    LocalMux I__14961 (
            .O(N__63368),
            .I(N__63328));
    Span4Mux_v I__14960 (
            .O(N__63365),
            .I(N__63325));
    InMux I__14959 (
            .O(N__63362),
            .I(N__63318));
    InMux I__14958 (
            .O(N__63359),
            .I(N__63318));
    InMux I__14957 (
            .O(N__63358),
            .I(N__63318));
    InMux I__14956 (
            .O(N__63357),
            .I(N__63315));
    InMux I__14955 (
            .O(N__63356),
            .I(N__63312));
    InMux I__14954 (
            .O(N__63355),
            .I(N__63305));
    InMux I__14953 (
            .O(N__63354),
            .I(N__63305));
    InMux I__14952 (
            .O(N__63353),
            .I(N__63305));
    Span4Mux_h I__14951 (
            .O(N__63348),
            .I(N__63300));
    LocalMux I__14950 (
            .O(N__63343),
            .I(N__63300));
    LocalMux I__14949 (
            .O(N__63340),
            .I(N__63295));
    LocalMux I__14948 (
            .O(N__63337),
            .I(N__63295));
    Span4Mux_h I__14947 (
            .O(N__63334),
            .I(N__63292));
    Span4Mux_h I__14946 (
            .O(N__63331),
            .I(N__63287));
    Span4Mux_h I__14945 (
            .O(N__63328),
            .I(N__63287));
    Sp12to4 I__14944 (
            .O(N__63325),
            .I(N__63282));
    LocalMux I__14943 (
            .O(N__63318),
            .I(N__63282));
    LocalMux I__14942 (
            .O(N__63315),
            .I(N__63273));
    LocalMux I__14941 (
            .O(N__63312),
            .I(N__63273));
    LocalMux I__14940 (
            .O(N__63305),
            .I(N__63273));
    Span4Mux_v I__14939 (
            .O(N__63300),
            .I(N__63270));
    Span12Mux_h I__14938 (
            .O(N__63295),
            .I(N__63265));
    Sp12to4 I__14937 (
            .O(N__63292),
            .I(N__63265));
    Sp12to4 I__14936 (
            .O(N__63287),
            .I(N__63260));
    Span12Mux_h I__14935 (
            .O(N__63282),
            .I(N__63260));
    InMux I__14934 (
            .O(N__63281),
            .I(N__63257));
    InMux I__14933 (
            .O(N__63280),
            .I(N__63254));
    Span4Mux_v I__14932 (
            .O(N__63273),
            .I(N__63251));
    Sp12to4 I__14931 (
            .O(N__63270),
            .I(N__63246));
    Span12Mux_v I__14930 (
            .O(N__63265),
            .I(N__63246));
    Span12Mux_v I__14929 (
            .O(N__63260),
            .I(N__63243));
    LocalMux I__14928 (
            .O(N__63257),
            .I(\c0.n19115 ));
    LocalMux I__14927 (
            .O(N__63254),
            .I(\c0.n19115 ));
    Odrv4 I__14926 (
            .O(N__63251),
            .I(\c0.n19115 ));
    Odrv12 I__14925 (
            .O(N__63246),
            .I(\c0.n19115 ));
    Odrv12 I__14924 (
            .O(N__63243),
            .I(\c0.n19115 ));
    InMux I__14923 (
            .O(N__63232),
            .I(N__63228));
    InMux I__14922 (
            .O(N__63231),
            .I(N__63225));
    LocalMux I__14921 (
            .O(N__63228),
            .I(N__63219));
    LocalMux I__14920 (
            .O(N__63225),
            .I(N__63219));
    InMux I__14919 (
            .O(N__63224),
            .I(N__63215));
    Span4Mux_h I__14918 (
            .O(N__63219),
            .I(N__63212));
    InMux I__14917 (
            .O(N__63218),
            .I(N__63209));
    LocalMux I__14916 (
            .O(N__63215),
            .I(\c0.data_in_frame_9_3 ));
    Odrv4 I__14915 (
            .O(N__63212),
            .I(\c0.data_in_frame_9_3 ));
    LocalMux I__14914 (
            .O(N__63209),
            .I(\c0.data_in_frame_9_3 ));
    InMux I__14913 (
            .O(N__63202),
            .I(N__63198));
    InMux I__14912 (
            .O(N__63201),
            .I(N__63194));
    LocalMux I__14911 (
            .O(N__63198),
            .I(N__63191));
    InMux I__14910 (
            .O(N__63197),
            .I(N__63188));
    LocalMux I__14909 (
            .O(N__63194),
            .I(\c0.data_in_frame_11_5 ));
    Odrv12 I__14908 (
            .O(N__63191),
            .I(\c0.data_in_frame_11_5 ));
    LocalMux I__14907 (
            .O(N__63188),
            .I(\c0.data_in_frame_11_5 ));
    InMux I__14906 (
            .O(N__63181),
            .I(N__63175));
    InMux I__14905 (
            .O(N__63180),
            .I(N__63175));
    LocalMux I__14904 (
            .O(N__63175),
            .I(N__63172));
    Span12Mux_h I__14903 (
            .O(N__63172),
            .I(N__63169));
    Odrv12 I__14902 (
            .O(N__63169),
            .I(\c0.n5_adj_3043 ));
    CascadeMux I__14901 (
            .O(N__63166),
            .I(N__63163));
    InMux I__14900 (
            .O(N__63163),
            .I(N__63159));
    InMux I__14899 (
            .O(N__63162),
            .I(N__63156));
    LocalMux I__14898 (
            .O(N__63159),
            .I(N__63150));
    LocalMux I__14897 (
            .O(N__63156),
            .I(N__63150));
    InMux I__14896 (
            .O(N__63155),
            .I(N__63145));
    Span4Mux_v I__14895 (
            .O(N__63150),
            .I(N__63142));
    CascadeMux I__14894 (
            .O(N__63149),
            .I(N__63139));
    CascadeMux I__14893 (
            .O(N__63148),
            .I(N__63136));
    LocalMux I__14892 (
            .O(N__63145),
            .I(N__63132));
    Span4Mux_h I__14891 (
            .O(N__63142),
            .I(N__63129));
    InMux I__14890 (
            .O(N__63139),
            .I(N__63124));
    InMux I__14889 (
            .O(N__63136),
            .I(N__63124));
    InMux I__14888 (
            .O(N__63135),
            .I(N__63121));
    Span12Mux_v I__14887 (
            .O(N__63132),
            .I(N__63118));
    Odrv4 I__14886 (
            .O(N__63129),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__14885 (
            .O(N__63124),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__14884 (
            .O(N__63121),
            .I(\c0.data_in_frame_7_1 ));
    Odrv12 I__14883 (
            .O(N__63118),
            .I(\c0.data_in_frame_7_1 ));
    InMux I__14882 (
            .O(N__63109),
            .I(N__63106));
    LocalMux I__14881 (
            .O(N__63106),
            .I(N__63101));
    InMux I__14880 (
            .O(N__63105),
            .I(N__63096));
    InMux I__14879 (
            .O(N__63104),
            .I(N__63093));
    Span4Mux_h I__14878 (
            .O(N__63101),
            .I(N__63090));
    InMux I__14877 (
            .O(N__63100),
            .I(N__63087));
    InMux I__14876 (
            .O(N__63099),
            .I(N__63084));
    LocalMux I__14875 (
            .O(N__63096),
            .I(N__63081));
    LocalMux I__14874 (
            .O(N__63093),
            .I(\c0.data_in_frame_9_0 ));
    Odrv4 I__14873 (
            .O(N__63090),
            .I(\c0.data_in_frame_9_0 ));
    LocalMux I__14872 (
            .O(N__63087),
            .I(\c0.data_in_frame_9_0 ));
    LocalMux I__14871 (
            .O(N__63084),
            .I(\c0.data_in_frame_9_0 ));
    Odrv12 I__14870 (
            .O(N__63081),
            .I(\c0.data_in_frame_9_0 ));
    CascadeMux I__14869 (
            .O(N__63070),
            .I(N__63067));
    InMux I__14868 (
            .O(N__63067),
            .I(N__63062));
    InMux I__14867 (
            .O(N__63066),
            .I(N__63057));
    InMux I__14866 (
            .O(N__63065),
            .I(N__63057));
    LocalMux I__14865 (
            .O(N__63062),
            .I(N__63054));
    LocalMux I__14864 (
            .O(N__63057),
            .I(\c0.data_in_frame_11_3 ));
    Odrv12 I__14863 (
            .O(N__63054),
            .I(\c0.data_in_frame_11_3 ));
    InMux I__14862 (
            .O(N__63049),
            .I(N__63045));
    CascadeMux I__14861 (
            .O(N__63048),
            .I(N__63041));
    LocalMux I__14860 (
            .O(N__63045),
            .I(N__63038));
    InMux I__14859 (
            .O(N__63044),
            .I(N__63035));
    InMux I__14858 (
            .O(N__63041),
            .I(N__63031));
    Span4Mux_v I__14857 (
            .O(N__63038),
            .I(N__63028));
    LocalMux I__14856 (
            .O(N__63035),
            .I(N__63025));
    InMux I__14855 (
            .O(N__63034),
            .I(N__63022));
    LocalMux I__14854 (
            .O(N__63031),
            .I(\c0.data_in_frame_13_4 ));
    Odrv4 I__14853 (
            .O(N__63028),
            .I(\c0.data_in_frame_13_4 ));
    Odrv4 I__14852 (
            .O(N__63025),
            .I(\c0.data_in_frame_13_4 ));
    LocalMux I__14851 (
            .O(N__63022),
            .I(\c0.data_in_frame_13_4 ));
    CascadeMux I__14850 (
            .O(N__63013),
            .I(N__63010));
    InMux I__14849 (
            .O(N__63010),
            .I(N__63007));
    LocalMux I__14848 (
            .O(N__63007),
            .I(N__63004));
    Span4Mux_v I__14847 (
            .O(N__63004),
            .I(N__63001));
    Span4Mux_h I__14846 (
            .O(N__63001),
            .I(N__62998));
    Odrv4 I__14845 (
            .O(N__62998),
            .I(\c0.n11_adj_3492 ));
    CascadeMux I__14844 (
            .O(N__62995),
            .I(\c0.n11_adj_3492_cascade_ ));
    InMux I__14843 (
            .O(N__62992),
            .I(N__62989));
    LocalMux I__14842 (
            .O(N__62989),
            .I(N__62985));
    InMux I__14841 (
            .O(N__62988),
            .I(N__62982));
    Span4Mux_v I__14840 (
            .O(N__62985),
            .I(N__62976));
    LocalMux I__14839 (
            .O(N__62982),
            .I(N__62976));
    InMux I__14838 (
            .O(N__62981),
            .I(N__62973));
    Span4Mux_h I__14837 (
            .O(N__62976),
            .I(N__62970));
    LocalMux I__14836 (
            .O(N__62973),
            .I(N__62965));
    Span4Mux_h I__14835 (
            .O(N__62970),
            .I(N__62962));
    InMux I__14834 (
            .O(N__62969),
            .I(N__62957));
    InMux I__14833 (
            .O(N__62968),
            .I(N__62957));
    Odrv4 I__14832 (
            .O(N__62965),
            .I(data_in_frame_16_0));
    Odrv4 I__14831 (
            .O(N__62962),
            .I(data_in_frame_16_0));
    LocalMux I__14830 (
            .O(N__62957),
            .I(data_in_frame_16_0));
    InMux I__14829 (
            .O(N__62950),
            .I(N__62947));
    LocalMux I__14828 (
            .O(N__62947),
            .I(N__62944));
    Span4Mux_h I__14827 (
            .O(N__62944),
            .I(N__62941));
    Span4Mux_v I__14826 (
            .O(N__62941),
            .I(N__62938));
    Odrv4 I__14825 (
            .O(N__62938),
            .I(\c0.n20_adj_3527 ));
    InMux I__14824 (
            .O(N__62935),
            .I(N__62931));
    CascadeMux I__14823 (
            .O(N__62934),
            .I(N__62928));
    LocalMux I__14822 (
            .O(N__62931),
            .I(N__62923));
    InMux I__14821 (
            .O(N__62928),
            .I(N__62916));
    InMux I__14820 (
            .O(N__62927),
            .I(N__62916));
    InMux I__14819 (
            .O(N__62926),
            .I(N__62916));
    Odrv4 I__14818 (
            .O(N__62923),
            .I(\c0.data_in_frame_11_1 ));
    LocalMux I__14817 (
            .O(N__62916),
            .I(\c0.data_in_frame_11_1 ));
    InMux I__14816 (
            .O(N__62911),
            .I(N__62908));
    LocalMux I__14815 (
            .O(N__62908),
            .I(N__62905));
    Span4Mux_h I__14814 (
            .O(N__62905),
            .I(N__62901));
    InMux I__14813 (
            .O(N__62904),
            .I(N__62898));
    Span4Mux_h I__14812 (
            .O(N__62901),
            .I(N__62895));
    LocalMux I__14811 (
            .O(N__62898),
            .I(\c0.n19229 ));
    Odrv4 I__14810 (
            .O(N__62895),
            .I(\c0.n19229 ));
    InMux I__14809 (
            .O(N__62890),
            .I(N__62886));
    InMux I__14808 (
            .O(N__62889),
            .I(N__62882));
    LocalMux I__14807 (
            .O(N__62886),
            .I(N__62879));
    CascadeMux I__14806 (
            .O(N__62885),
            .I(N__62875));
    LocalMux I__14805 (
            .O(N__62882),
            .I(N__62872));
    Span4Mux_v I__14804 (
            .O(N__62879),
            .I(N__62869));
    CascadeMux I__14803 (
            .O(N__62878),
            .I(N__62866));
    InMux I__14802 (
            .O(N__62875),
            .I(N__62863));
    Span4Mux_v I__14801 (
            .O(N__62872),
            .I(N__62858));
    Span4Mux_h I__14800 (
            .O(N__62869),
            .I(N__62858));
    InMux I__14799 (
            .O(N__62866),
            .I(N__62855));
    LocalMux I__14798 (
            .O(N__62863),
            .I(\c0.data_in_frame_11_2 ));
    Odrv4 I__14797 (
            .O(N__62858),
            .I(\c0.data_in_frame_11_2 ));
    LocalMux I__14796 (
            .O(N__62855),
            .I(\c0.data_in_frame_11_2 ));
    InMux I__14795 (
            .O(N__62848),
            .I(N__62839));
    InMux I__14794 (
            .O(N__62847),
            .I(N__62839));
    InMux I__14793 (
            .O(N__62846),
            .I(N__62834));
    InMux I__14792 (
            .O(N__62845),
            .I(N__62831));
    InMux I__14791 (
            .O(N__62844),
            .I(N__62827));
    LocalMux I__14790 (
            .O(N__62839),
            .I(N__62824));
    InMux I__14789 (
            .O(N__62838),
            .I(N__62819));
    InMux I__14788 (
            .O(N__62837),
            .I(N__62819));
    LocalMux I__14787 (
            .O(N__62834),
            .I(N__62816));
    LocalMux I__14786 (
            .O(N__62831),
            .I(N__62813));
    InMux I__14785 (
            .O(N__62830),
            .I(N__62807));
    LocalMux I__14784 (
            .O(N__62827),
            .I(N__62804));
    Span4Mux_v I__14783 (
            .O(N__62824),
            .I(N__62798));
    LocalMux I__14782 (
            .O(N__62819),
            .I(N__62795));
    Span4Mux_v I__14781 (
            .O(N__62816),
            .I(N__62788));
    Span4Mux_v I__14780 (
            .O(N__62813),
            .I(N__62788));
    InMux I__14779 (
            .O(N__62812),
            .I(N__62785));
    InMux I__14778 (
            .O(N__62811),
            .I(N__62782));
    InMux I__14777 (
            .O(N__62810),
            .I(N__62779));
    LocalMux I__14776 (
            .O(N__62807),
            .I(N__62774));
    Span4Mux_v I__14775 (
            .O(N__62804),
            .I(N__62774));
    InMux I__14774 (
            .O(N__62803),
            .I(N__62771));
    InMux I__14773 (
            .O(N__62802),
            .I(N__62766));
    InMux I__14772 (
            .O(N__62801),
            .I(N__62766));
    Sp12to4 I__14771 (
            .O(N__62798),
            .I(N__62763));
    Sp12to4 I__14770 (
            .O(N__62795),
            .I(N__62760));
    InMux I__14769 (
            .O(N__62794),
            .I(N__62755));
    InMux I__14768 (
            .O(N__62793),
            .I(N__62755));
    Sp12to4 I__14767 (
            .O(N__62788),
            .I(N__62752));
    LocalMux I__14766 (
            .O(N__62785),
            .I(N__62743));
    LocalMux I__14765 (
            .O(N__62782),
            .I(N__62743));
    LocalMux I__14764 (
            .O(N__62779),
            .I(N__62743));
    Sp12to4 I__14763 (
            .O(N__62774),
            .I(N__62743));
    LocalMux I__14762 (
            .O(N__62771),
            .I(N__62734));
    LocalMux I__14761 (
            .O(N__62766),
            .I(N__62734));
    Span12Mux_h I__14760 (
            .O(N__62763),
            .I(N__62734));
    Span12Mux_s11_v I__14759 (
            .O(N__62760),
            .I(N__62734));
    LocalMux I__14758 (
            .O(N__62755),
            .I(\c0.n19134 ));
    Odrv12 I__14757 (
            .O(N__62752),
            .I(\c0.n19134 ));
    Odrv12 I__14756 (
            .O(N__62743),
            .I(\c0.n19134 ));
    Odrv12 I__14755 (
            .O(N__62734),
            .I(\c0.n19134 ));
    CascadeMux I__14754 (
            .O(N__62725),
            .I(N__62721));
    CascadeMux I__14753 (
            .O(N__62724),
            .I(N__62717));
    InMux I__14752 (
            .O(N__62721),
            .I(N__62713));
    InMux I__14751 (
            .O(N__62720),
            .I(N__62710));
    InMux I__14750 (
            .O(N__62717),
            .I(N__62705));
    InMux I__14749 (
            .O(N__62716),
            .I(N__62705));
    LocalMux I__14748 (
            .O(N__62713),
            .I(\c0.data_in_frame_10_7 ));
    LocalMux I__14747 (
            .O(N__62710),
            .I(\c0.data_in_frame_10_7 ));
    LocalMux I__14746 (
            .O(N__62705),
            .I(\c0.data_in_frame_10_7 ));
    CascadeMux I__14745 (
            .O(N__62698),
            .I(N__62695));
    InMux I__14744 (
            .O(N__62695),
            .I(N__62692));
    LocalMux I__14743 (
            .O(N__62692),
            .I(N__62689));
    Span4Mux_h I__14742 (
            .O(N__62689),
            .I(N__62686));
    Odrv4 I__14741 (
            .O(N__62686),
            .I(\c0.n6_adj_3037 ));
    InMux I__14740 (
            .O(N__62683),
            .I(N__62676));
    InMux I__14739 (
            .O(N__62682),
            .I(N__62673));
    CascadeMux I__14738 (
            .O(N__62681),
            .I(N__62670));
    InMux I__14737 (
            .O(N__62680),
            .I(N__62667));
    InMux I__14736 (
            .O(N__62679),
            .I(N__62664));
    LocalMux I__14735 (
            .O(N__62676),
            .I(N__62659));
    LocalMux I__14734 (
            .O(N__62673),
            .I(N__62659));
    InMux I__14733 (
            .O(N__62670),
            .I(N__62655));
    LocalMux I__14732 (
            .O(N__62667),
            .I(N__62650));
    LocalMux I__14731 (
            .O(N__62664),
            .I(N__62650));
    Span12Mux_v I__14730 (
            .O(N__62659),
            .I(N__62647));
    InMux I__14729 (
            .O(N__62658),
            .I(N__62644));
    LocalMux I__14728 (
            .O(N__62655),
            .I(\c0.data_in_frame_5_7 ));
    Odrv12 I__14727 (
            .O(N__62650),
            .I(\c0.data_in_frame_5_7 ));
    Odrv12 I__14726 (
            .O(N__62647),
            .I(\c0.data_in_frame_5_7 ));
    LocalMux I__14725 (
            .O(N__62644),
            .I(\c0.data_in_frame_5_7 ));
    InMux I__14724 (
            .O(N__62635),
            .I(N__62632));
    LocalMux I__14723 (
            .O(N__62632),
            .I(\c0.n4_adj_3036 ));
    CascadeMux I__14722 (
            .O(N__62629),
            .I(\c0.n6_adj_3037_cascade_ ));
    CascadeMux I__14721 (
            .O(N__62626),
            .I(N__62621));
    InMux I__14720 (
            .O(N__62625),
            .I(N__62615));
    InMux I__14719 (
            .O(N__62624),
            .I(N__62612));
    InMux I__14718 (
            .O(N__62621),
            .I(N__62609));
    InMux I__14717 (
            .O(N__62620),
            .I(N__62606));
    InMux I__14716 (
            .O(N__62619),
            .I(N__62601));
    InMux I__14715 (
            .O(N__62618),
            .I(N__62601));
    LocalMux I__14714 (
            .O(N__62615),
            .I(N__62596));
    LocalMux I__14713 (
            .O(N__62612),
            .I(N__62596));
    LocalMux I__14712 (
            .O(N__62609),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__14711 (
            .O(N__62606),
            .I(\c0.data_in_frame_3_5 ));
    LocalMux I__14710 (
            .O(N__62601),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__14709 (
            .O(N__62596),
            .I(\c0.data_in_frame_3_5 ));
    InMux I__14708 (
            .O(N__62587),
            .I(N__62584));
    LocalMux I__14707 (
            .O(N__62584),
            .I(N__62579));
    InMux I__14706 (
            .O(N__62583),
            .I(N__62576));
    InMux I__14705 (
            .O(N__62582),
            .I(N__62573));
    Span4Mux_h I__14704 (
            .O(N__62579),
            .I(N__62570));
    LocalMux I__14703 (
            .O(N__62576),
            .I(N__62567));
    LocalMux I__14702 (
            .O(N__62573),
            .I(N__62564));
    Span4Mux_h I__14701 (
            .O(N__62570),
            .I(N__62561));
    Span4Mux_h I__14700 (
            .O(N__62567),
            .I(N__62556));
    Span4Mux_h I__14699 (
            .O(N__62564),
            .I(N__62556));
    Odrv4 I__14698 (
            .O(N__62561),
            .I(\c0.n19560 ));
    Odrv4 I__14697 (
            .O(N__62556),
            .I(\c0.n19560 ));
    CascadeMux I__14696 (
            .O(N__62551),
            .I(N__62548));
    InMux I__14695 (
            .O(N__62548),
            .I(N__62545));
    LocalMux I__14694 (
            .O(N__62545),
            .I(N__62541));
    CascadeMux I__14693 (
            .O(N__62544),
            .I(N__62538));
    Span4Mux_v I__14692 (
            .O(N__62541),
            .I(N__62535));
    InMux I__14691 (
            .O(N__62538),
            .I(N__62532));
    Odrv4 I__14690 (
            .O(N__62535),
            .I(\c0.data_out_frame_0__7__N_1540 ));
    LocalMux I__14689 (
            .O(N__62532),
            .I(\c0.data_out_frame_0__7__N_1540 ));
    InMux I__14688 (
            .O(N__62527),
            .I(N__62524));
    LocalMux I__14687 (
            .O(N__62524),
            .I(N__62519));
    InMux I__14686 (
            .O(N__62523),
            .I(N__62516));
    CascadeMux I__14685 (
            .O(N__62522),
            .I(N__62513));
    Span4Mux_v I__14684 (
            .O(N__62519),
            .I(N__62507));
    LocalMux I__14683 (
            .O(N__62516),
            .I(N__62507));
    InMux I__14682 (
            .O(N__62513),
            .I(N__62502));
    InMux I__14681 (
            .O(N__62512),
            .I(N__62502));
    Odrv4 I__14680 (
            .O(N__62507),
            .I(\c0.data_in_frame_6_6 ));
    LocalMux I__14679 (
            .O(N__62502),
            .I(\c0.data_in_frame_6_6 ));
    InMux I__14678 (
            .O(N__62497),
            .I(N__62492));
    CascadeMux I__14677 (
            .O(N__62496),
            .I(N__62489));
    InMux I__14676 (
            .O(N__62495),
            .I(N__62486));
    LocalMux I__14675 (
            .O(N__62492),
            .I(N__62483));
    InMux I__14674 (
            .O(N__62489),
            .I(N__62480));
    LocalMux I__14673 (
            .O(N__62486),
            .I(N__62477));
    Span4Mux_v I__14672 (
            .O(N__62483),
            .I(N__62474));
    LocalMux I__14671 (
            .O(N__62480),
            .I(\c0.n19258 ));
    Odrv4 I__14670 (
            .O(N__62477),
            .I(\c0.n19258 ));
    Odrv4 I__14669 (
            .O(N__62474),
            .I(\c0.n19258 ));
    InMux I__14668 (
            .O(N__62467),
            .I(N__62461));
    InMux I__14667 (
            .O(N__62466),
            .I(N__62456));
    InMux I__14666 (
            .O(N__62465),
            .I(N__62456));
    CascadeMux I__14665 (
            .O(N__62464),
            .I(N__62453));
    LocalMux I__14664 (
            .O(N__62461),
            .I(N__62448));
    LocalMux I__14663 (
            .O(N__62456),
            .I(N__62448));
    InMux I__14662 (
            .O(N__62453),
            .I(N__62444));
    Span4Mux_v I__14661 (
            .O(N__62448),
            .I(N__62441));
    InMux I__14660 (
            .O(N__62447),
            .I(N__62437));
    LocalMux I__14659 (
            .O(N__62444),
            .I(N__62434));
    Span4Mux_h I__14658 (
            .O(N__62441),
            .I(N__62431));
    InMux I__14657 (
            .O(N__62440),
            .I(N__62428));
    LocalMux I__14656 (
            .O(N__62437),
            .I(\c0.data_in_frame_8_0 ));
    Odrv4 I__14655 (
            .O(N__62434),
            .I(\c0.data_in_frame_8_0 ));
    Odrv4 I__14654 (
            .O(N__62431),
            .I(\c0.data_in_frame_8_0 ));
    LocalMux I__14653 (
            .O(N__62428),
            .I(\c0.data_in_frame_8_0 ));
    InMux I__14652 (
            .O(N__62419),
            .I(N__62415));
    InMux I__14651 (
            .O(N__62418),
            .I(N__62412));
    LocalMux I__14650 (
            .O(N__62415),
            .I(N__62406));
    LocalMux I__14649 (
            .O(N__62412),
            .I(N__62403));
    InMux I__14648 (
            .O(N__62411),
            .I(N__62400));
    CascadeMux I__14647 (
            .O(N__62410),
            .I(N__62396));
    InMux I__14646 (
            .O(N__62409),
            .I(N__62393));
    Span4Mux_v I__14645 (
            .O(N__62406),
            .I(N__62386));
    Span4Mux_v I__14644 (
            .O(N__62403),
            .I(N__62386));
    LocalMux I__14643 (
            .O(N__62400),
            .I(N__62386));
    InMux I__14642 (
            .O(N__62399),
            .I(N__62383));
    InMux I__14641 (
            .O(N__62396),
            .I(N__62379));
    LocalMux I__14640 (
            .O(N__62393),
            .I(N__62374));
    Span4Mux_h I__14639 (
            .O(N__62386),
            .I(N__62374));
    LocalMux I__14638 (
            .O(N__62383),
            .I(N__62371));
    InMux I__14637 (
            .O(N__62382),
            .I(N__62368));
    LocalMux I__14636 (
            .O(N__62379),
            .I(\c0.data_in_frame_7_7 ));
    Odrv4 I__14635 (
            .O(N__62374),
            .I(\c0.data_in_frame_7_7 ));
    Odrv4 I__14634 (
            .O(N__62371),
            .I(\c0.data_in_frame_7_7 ));
    LocalMux I__14633 (
            .O(N__62368),
            .I(\c0.data_in_frame_7_7 ));
    CascadeMux I__14632 (
            .O(N__62359),
            .I(N__62356));
    InMux I__14631 (
            .O(N__62356),
            .I(N__62350));
    InMux I__14630 (
            .O(N__62355),
            .I(N__62347));
    InMux I__14629 (
            .O(N__62354),
            .I(N__62344));
    InMux I__14628 (
            .O(N__62353),
            .I(N__62340));
    LocalMux I__14627 (
            .O(N__62350),
            .I(N__62335));
    LocalMux I__14626 (
            .O(N__62347),
            .I(N__62335));
    LocalMux I__14625 (
            .O(N__62344),
            .I(N__62332));
    InMux I__14624 (
            .O(N__62343),
            .I(N__62329));
    LocalMux I__14623 (
            .O(N__62340),
            .I(\c0.data_in_frame_5_6 ));
    Odrv4 I__14622 (
            .O(N__62335),
            .I(\c0.data_in_frame_5_6 ));
    Odrv4 I__14621 (
            .O(N__62332),
            .I(\c0.data_in_frame_5_6 ));
    LocalMux I__14620 (
            .O(N__62329),
            .I(\c0.data_in_frame_5_6 ));
    InMux I__14619 (
            .O(N__62320),
            .I(N__62317));
    LocalMux I__14618 (
            .O(N__62317),
            .I(\c0.n8_adj_3020 ));
    CascadeMux I__14617 (
            .O(N__62314),
            .I(N__62310));
    CascadeMux I__14616 (
            .O(N__62313),
            .I(N__62304));
    InMux I__14615 (
            .O(N__62310),
            .I(N__62301));
    CascadeMux I__14614 (
            .O(N__62309),
            .I(N__62298));
    InMux I__14613 (
            .O(N__62308),
            .I(N__62293));
    InMux I__14612 (
            .O(N__62307),
            .I(N__62293));
    InMux I__14611 (
            .O(N__62304),
            .I(N__62290));
    LocalMux I__14610 (
            .O(N__62301),
            .I(N__62287));
    InMux I__14609 (
            .O(N__62298),
            .I(N__62284));
    LocalMux I__14608 (
            .O(N__62293),
            .I(N__62281));
    LocalMux I__14607 (
            .O(N__62290),
            .I(N__62278));
    Span4Mux_v I__14606 (
            .O(N__62287),
            .I(N__62275));
    LocalMux I__14605 (
            .O(N__62284),
            .I(N__62270));
    Span4Mux_v I__14604 (
            .O(N__62281),
            .I(N__62270));
    Span4Mux_h I__14603 (
            .O(N__62278),
            .I(N__62267));
    Span4Mux_h I__14602 (
            .O(N__62275),
            .I(N__62264));
    Odrv4 I__14601 (
            .O(N__62270),
            .I(\c0.data_in_frame_13_3 ));
    Odrv4 I__14600 (
            .O(N__62267),
            .I(\c0.data_in_frame_13_3 ));
    Odrv4 I__14599 (
            .O(N__62264),
            .I(\c0.data_in_frame_13_3 ));
    InMux I__14598 (
            .O(N__62257),
            .I(N__62251));
    InMux I__14597 (
            .O(N__62256),
            .I(N__62247));
    InMux I__14596 (
            .O(N__62255),
            .I(N__62244));
    CascadeMux I__14595 (
            .O(N__62254),
            .I(N__62241));
    LocalMux I__14594 (
            .O(N__62251),
            .I(N__62238));
    InMux I__14593 (
            .O(N__62250),
            .I(N__62235));
    LocalMux I__14592 (
            .O(N__62247),
            .I(N__62232));
    LocalMux I__14591 (
            .O(N__62244),
            .I(N__62229));
    InMux I__14590 (
            .O(N__62241),
            .I(N__62226));
    Span4Mux_v I__14589 (
            .O(N__62238),
            .I(N__62223));
    LocalMux I__14588 (
            .O(N__62235),
            .I(N__62218));
    Span4Mux_h I__14587 (
            .O(N__62232),
            .I(N__62218));
    Span12Mux_v I__14586 (
            .O(N__62229),
            .I(N__62215));
    LocalMux I__14585 (
            .O(N__62226),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__14584 (
            .O(N__62223),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__14583 (
            .O(N__62218),
            .I(\c0.data_in_frame_9_2 ));
    Odrv12 I__14582 (
            .O(N__62215),
            .I(\c0.data_in_frame_9_2 ));
    InMux I__14581 (
            .O(N__62206),
            .I(N__62203));
    LocalMux I__14580 (
            .O(N__62203),
            .I(N__62200));
    Span4Mux_h I__14579 (
            .O(N__62200),
            .I(N__62194));
    InMux I__14578 (
            .O(N__62199),
            .I(N__62187));
    InMux I__14577 (
            .O(N__62198),
            .I(N__62187));
    InMux I__14576 (
            .O(N__62197),
            .I(N__62187));
    Odrv4 I__14575 (
            .O(N__62194),
            .I(\c0.n20095 ));
    LocalMux I__14574 (
            .O(N__62187),
            .I(\c0.n20095 ));
    InMux I__14573 (
            .O(N__62182),
            .I(N__62177));
    InMux I__14572 (
            .O(N__62181),
            .I(N__62173));
    InMux I__14571 (
            .O(N__62180),
            .I(N__62169));
    LocalMux I__14570 (
            .O(N__62177),
            .I(N__62166));
    InMux I__14569 (
            .O(N__62176),
            .I(N__62160));
    LocalMux I__14568 (
            .O(N__62173),
            .I(N__62157));
    InMux I__14567 (
            .O(N__62172),
            .I(N__62153));
    LocalMux I__14566 (
            .O(N__62169),
            .I(N__62148));
    Span4Mux_v I__14565 (
            .O(N__62166),
            .I(N__62148));
    InMux I__14564 (
            .O(N__62165),
            .I(N__62145));
    InMux I__14563 (
            .O(N__62164),
            .I(N__62140));
    InMux I__14562 (
            .O(N__62163),
            .I(N__62140));
    LocalMux I__14561 (
            .O(N__62160),
            .I(N__62135));
    Span4Mux_v I__14560 (
            .O(N__62157),
            .I(N__62135));
    InMux I__14559 (
            .O(N__62156),
            .I(N__62132));
    LocalMux I__14558 (
            .O(N__62153),
            .I(N__62123));
    Span4Mux_h I__14557 (
            .O(N__62148),
            .I(N__62118));
    LocalMux I__14556 (
            .O(N__62145),
            .I(N__62118));
    LocalMux I__14555 (
            .O(N__62140),
            .I(N__62111));
    Span4Mux_h I__14554 (
            .O(N__62135),
            .I(N__62111));
    LocalMux I__14553 (
            .O(N__62132),
            .I(N__62111));
    InMux I__14552 (
            .O(N__62131),
            .I(N__62108));
    InMux I__14551 (
            .O(N__62130),
            .I(N__62105));
    InMux I__14550 (
            .O(N__62129),
            .I(N__62100));
    InMux I__14549 (
            .O(N__62128),
            .I(N__62100));
    InMux I__14548 (
            .O(N__62127),
            .I(N__62095));
    InMux I__14547 (
            .O(N__62126),
            .I(N__62095));
    Odrv4 I__14546 (
            .O(N__62123),
            .I(data_in_frame_0_3));
    Odrv4 I__14545 (
            .O(N__62118),
            .I(data_in_frame_0_3));
    Odrv4 I__14544 (
            .O(N__62111),
            .I(data_in_frame_0_3));
    LocalMux I__14543 (
            .O(N__62108),
            .I(data_in_frame_0_3));
    LocalMux I__14542 (
            .O(N__62105),
            .I(data_in_frame_0_3));
    LocalMux I__14541 (
            .O(N__62100),
            .I(data_in_frame_0_3));
    LocalMux I__14540 (
            .O(N__62095),
            .I(data_in_frame_0_3));
    CascadeMux I__14539 (
            .O(N__62080),
            .I(N__62077));
    InMux I__14538 (
            .O(N__62077),
            .I(N__62073));
    InMux I__14537 (
            .O(N__62076),
            .I(N__62070));
    LocalMux I__14536 (
            .O(N__62073),
            .I(N__62067));
    LocalMux I__14535 (
            .O(N__62070),
            .I(\c0.n5240 ));
    Odrv12 I__14534 (
            .O(N__62067),
            .I(\c0.n5240 ));
    CascadeMux I__14533 (
            .O(N__62062),
            .I(\c0.n7_cascade_ ));
    InMux I__14532 (
            .O(N__62059),
            .I(N__62053));
    InMux I__14531 (
            .O(N__62058),
            .I(N__62053));
    LocalMux I__14530 (
            .O(N__62053),
            .I(N__62050));
    Span4Mux_v I__14529 (
            .O(N__62050),
            .I(N__62045));
    CascadeMux I__14528 (
            .O(N__62049),
            .I(N__62042));
    CascadeMux I__14527 (
            .O(N__62048),
            .I(N__62036));
    Span4Mux_h I__14526 (
            .O(N__62045),
            .I(N__62031));
    InMux I__14525 (
            .O(N__62042),
            .I(N__62027));
    InMux I__14524 (
            .O(N__62041),
            .I(N__62024));
    InMux I__14523 (
            .O(N__62040),
            .I(N__62019));
    InMux I__14522 (
            .O(N__62039),
            .I(N__62019));
    InMux I__14521 (
            .O(N__62036),
            .I(N__62013));
    InMux I__14520 (
            .O(N__62035),
            .I(N__62013));
    InMux I__14519 (
            .O(N__62034),
            .I(N__62010));
    Span4Mux_v I__14518 (
            .O(N__62031),
            .I(N__62006));
    InMux I__14517 (
            .O(N__62030),
            .I(N__62003));
    LocalMux I__14516 (
            .O(N__62027),
            .I(N__61997));
    LocalMux I__14515 (
            .O(N__62024),
            .I(N__61997));
    LocalMux I__14514 (
            .O(N__62019),
            .I(N__61994));
    InMux I__14513 (
            .O(N__62018),
            .I(N__61991));
    LocalMux I__14512 (
            .O(N__62013),
            .I(N__61988));
    LocalMux I__14511 (
            .O(N__62010),
            .I(N__61984));
    InMux I__14510 (
            .O(N__62009),
            .I(N__61981));
    Span4Mux_h I__14509 (
            .O(N__62006),
            .I(N__61976));
    LocalMux I__14508 (
            .O(N__62003),
            .I(N__61976));
    CascadeMux I__14507 (
            .O(N__62002),
            .I(N__61973));
    Span4Mux_v I__14506 (
            .O(N__61997),
            .I(N__61968));
    Span4Mux_v I__14505 (
            .O(N__61994),
            .I(N__61968));
    LocalMux I__14504 (
            .O(N__61991),
            .I(N__61965));
    Span4Mux_v I__14503 (
            .O(N__61988),
            .I(N__61962));
    CascadeMux I__14502 (
            .O(N__61987),
            .I(N__61959));
    Span4Mux_v I__14501 (
            .O(N__61984),
            .I(N__61956));
    LocalMux I__14500 (
            .O(N__61981),
            .I(N__61951));
    Span4Mux_v I__14499 (
            .O(N__61976),
            .I(N__61948));
    InMux I__14498 (
            .O(N__61973),
            .I(N__61945));
    Span4Mux_h I__14497 (
            .O(N__61968),
            .I(N__61942));
    Span4Mux_v I__14496 (
            .O(N__61965),
            .I(N__61937));
    Span4Mux_h I__14495 (
            .O(N__61962),
            .I(N__61937));
    InMux I__14494 (
            .O(N__61959),
            .I(N__61934));
    Sp12to4 I__14493 (
            .O(N__61956),
            .I(N__61931));
    InMux I__14492 (
            .O(N__61955),
            .I(N__61928));
    InMux I__14491 (
            .O(N__61954),
            .I(N__61924));
    Span4Mux_v I__14490 (
            .O(N__61951),
            .I(N__61921));
    Span4Mux_h I__14489 (
            .O(N__61948),
            .I(N__61916));
    LocalMux I__14488 (
            .O(N__61945),
            .I(N__61916));
    Span4Mux_h I__14487 (
            .O(N__61942),
            .I(N__61911));
    Span4Mux_v I__14486 (
            .O(N__61937),
            .I(N__61911));
    LocalMux I__14485 (
            .O(N__61934),
            .I(N__61904));
    Span12Mux_h I__14484 (
            .O(N__61931),
            .I(N__61904));
    LocalMux I__14483 (
            .O(N__61928),
            .I(N__61904));
    InMux I__14482 (
            .O(N__61927),
            .I(N__61901));
    LocalMux I__14481 (
            .O(N__61924),
            .I(N__61898));
    Span4Mux_h I__14480 (
            .O(N__61921),
            .I(N__61893));
    Span4Mux_h I__14479 (
            .O(N__61916),
            .I(N__61893));
    Sp12to4 I__14478 (
            .O(N__61911),
            .I(N__61888));
    Span12Mux_v I__14477 (
            .O(N__61904),
            .I(N__61888));
    LocalMux I__14476 (
            .O(N__61901),
            .I(\c0.n9_adj_3038 ));
    Odrv4 I__14475 (
            .O(N__61898),
            .I(\c0.n9_adj_3038 ));
    Odrv4 I__14474 (
            .O(N__61893),
            .I(\c0.n9_adj_3038 ));
    Odrv12 I__14473 (
            .O(N__61888),
            .I(\c0.n9_adj_3038 ));
    InMux I__14472 (
            .O(N__61879),
            .I(N__61875));
    InMux I__14471 (
            .O(N__61878),
            .I(N__61868));
    LocalMux I__14470 (
            .O(N__61875),
            .I(N__61865));
    InMux I__14469 (
            .O(N__61874),
            .I(N__61862));
    InMux I__14468 (
            .O(N__61873),
            .I(N__61857));
    InMux I__14467 (
            .O(N__61872),
            .I(N__61852));
    InMux I__14466 (
            .O(N__61871),
            .I(N__61852));
    LocalMux I__14465 (
            .O(N__61868),
            .I(N__61847));
    Span4Mux_h I__14464 (
            .O(N__61865),
            .I(N__61847));
    LocalMux I__14463 (
            .O(N__61862),
            .I(N__61844));
    CascadeMux I__14462 (
            .O(N__61861),
            .I(N__61841));
    InMux I__14461 (
            .O(N__61860),
            .I(N__61838));
    LocalMux I__14460 (
            .O(N__61857),
            .I(N__61833));
    LocalMux I__14459 (
            .O(N__61852),
            .I(N__61833));
    Span4Mux_v I__14458 (
            .O(N__61847),
            .I(N__61830));
    Span4Mux_h I__14457 (
            .O(N__61844),
            .I(N__61827));
    InMux I__14456 (
            .O(N__61841),
            .I(N__61823));
    LocalMux I__14455 (
            .O(N__61838),
            .I(N__61820));
    Span4Mux_v I__14454 (
            .O(N__61833),
            .I(N__61813));
    Span4Mux_h I__14453 (
            .O(N__61830),
            .I(N__61813));
    Span4Mux_h I__14452 (
            .O(N__61827),
            .I(N__61813));
    InMux I__14451 (
            .O(N__61826),
            .I(N__61810));
    LocalMux I__14450 (
            .O(N__61823),
            .I(\c0.data_in_frame_6_7 ));
    Odrv12 I__14449 (
            .O(N__61820),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__14448 (
            .O(N__61813),
            .I(\c0.data_in_frame_6_7 ));
    LocalMux I__14447 (
            .O(N__61810),
            .I(\c0.data_in_frame_6_7 ));
    InMux I__14446 (
            .O(N__61801),
            .I(N__61798));
    LocalMux I__14445 (
            .O(N__61798),
            .I(N__61791));
    InMux I__14444 (
            .O(N__61797),
            .I(N__61786));
    InMux I__14443 (
            .O(N__61796),
            .I(N__61786));
    InMux I__14442 (
            .O(N__61795),
            .I(N__61781));
    InMux I__14441 (
            .O(N__61794),
            .I(N__61781));
    Span4Mux_v I__14440 (
            .O(N__61791),
            .I(N__61774));
    LocalMux I__14439 (
            .O(N__61786),
            .I(N__61769));
    LocalMux I__14438 (
            .O(N__61781),
            .I(N__61769));
    InMux I__14437 (
            .O(N__61780),
            .I(N__61761));
    InMux I__14436 (
            .O(N__61779),
            .I(N__61761));
    CascadeMux I__14435 (
            .O(N__61778),
            .I(N__61749));
    CascadeMux I__14434 (
            .O(N__61777),
            .I(N__61746));
    Span4Mux_h I__14433 (
            .O(N__61774),
            .I(N__61739));
    Span4Mux_v I__14432 (
            .O(N__61769),
            .I(N__61739));
    InMux I__14431 (
            .O(N__61768),
            .I(N__61732));
    InMux I__14430 (
            .O(N__61767),
            .I(N__61732));
    InMux I__14429 (
            .O(N__61766),
            .I(N__61732));
    LocalMux I__14428 (
            .O(N__61761),
            .I(N__61727));
    InMux I__14427 (
            .O(N__61760),
            .I(N__61716));
    InMux I__14426 (
            .O(N__61759),
            .I(N__61716));
    InMux I__14425 (
            .O(N__61758),
            .I(N__61716));
    InMux I__14424 (
            .O(N__61757),
            .I(N__61713));
    InMux I__14423 (
            .O(N__61756),
            .I(N__61702));
    InMux I__14422 (
            .O(N__61755),
            .I(N__61702));
    InMux I__14421 (
            .O(N__61754),
            .I(N__61702));
    InMux I__14420 (
            .O(N__61753),
            .I(N__61702));
    InMux I__14419 (
            .O(N__61752),
            .I(N__61702));
    InMux I__14418 (
            .O(N__61749),
            .I(N__61693));
    InMux I__14417 (
            .O(N__61746),
            .I(N__61693));
    InMux I__14416 (
            .O(N__61745),
            .I(N__61693));
    InMux I__14415 (
            .O(N__61744),
            .I(N__61693));
    Span4Mux_h I__14414 (
            .O(N__61739),
            .I(N__61678));
    LocalMux I__14413 (
            .O(N__61732),
            .I(N__61678));
    InMux I__14412 (
            .O(N__61731),
            .I(N__61674));
    InMux I__14411 (
            .O(N__61730),
            .I(N__61667));
    Span4Mux_v I__14410 (
            .O(N__61727),
            .I(N__61664));
    InMux I__14409 (
            .O(N__61726),
            .I(N__61659));
    InMux I__14408 (
            .O(N__61725),
            .I(N__61659));
    InMux I__14407 (
            .O(N__61724),
            .I(N__61654));
    InMux I__14406 (
            .O(N__61723),
            .I(N__61654));
    LocalMux I__14405 (
            .O(N__61716),
            .I(N__61651));
    LocalMux I__14404 (
            .O(N__61713),
            .I(N__61644));
    LocalMux I__14403 (
            .O(N__61702),
            .I(N__61644));
    LocalMux I__14402 (
            .O(N__61693),
            .I(N__61644));
    InMux I__14401 (
            .O(N__61692),
            .I(N__61635));
    InMux I__14400 (
            .O(N__61691),
            .I(N__61635));
    InMux I__14399 (
            .O(N__61690),
            .I(N__61635));
    InMux I__14398 (
            .O(N__61689),
            .I(N__61635));
    InMux I__14397 (
            .O(N__61688),
            .I(N__61632));
    InMux I__14396 (
            .O(N__61687),
            .I(N__61627));
    InMux I__14395 (
            .O(N__61686),
            .I(N__61627));
    InMux I__14394 (
            .O(N__61685),
            .I(N__61624));
    InMux I__14393 (
            .O(N__61684),
            .I(N__61619));
    InMux I__14392 (
            .O(N__61683),
            .I(N__61619));
    Span4Mux_h I__14391 (
            .O(N__61678),
            .I(N__61616));
    InMux I__14390 (
            .O(N__61677),
            .I(N__61612));
    LocalMux I__14389 (
            .O(N__61674),
            .I(N__61609));
    InMux I__14388 (
            .O(N__61673),
            .I(N__61600));
    InMux I__14387 (
            .O(N__61672),
            .I(N__61600));
    InMux I__14386 (
            .O(N__61671),
            .I(N__61600));
    InMux I__14385 (
            .O(N__61670),
            .I(N__61600));
    LocalMux I__14384 (
            .O(N__61667),
            .I(N__61584));
    Span4Mux_h I__14383 (
            .O(N__61664),
            .I(N__61584));
    LocalMux I__14382 (
            .O(N__61659),
            .I(N__61584));
    LocalMux I__14381 (
            .O(N__61654),
            .I(N__61584));
    Span4Mux_v I__14380 (
            .O(N__61651),
            .I(N__61577));
    Span4Mux_v I__14379 (
            .O(N__61644),
            .I(N__61577));
    LocalMux I__14378 (
            .O(N__61635),
            .I(N__61577));
    LocalMux I__14377 (
            .O(N__61632),
            .I(N__61572));
    LocalMux I__14376 (
            .O(N__61627),
            .I(N__61572));
    LocalMux I__14375 (
            .O(N__61624),
            .I(N__61567));
    LocalMux I__14374 (
            .O(N__61619),
            .I(N__61567));
    Span4Mux_v I__14373 (
            .O(N__61616),
            .I(N__61564));
    InMux I__14372 (
            .O(N__61615),
            .I(N__61561));
    LocalMux I__14371 (
            .O(N__61612),
            .I(N__61553));
    Span4Mux_v I__14370 (
            .O(N__61609),
            .I(N__61553));
    LocalMux I__14369 (
            .O(N__61600),
            .I(N__61553));
    CascadeMux I__14368 (
            .O(N__61599),
            .I(N__61546));
    InMux I__14367 (
            .O(N__61598),
            .I(N__61543));
    InMux I__14366 (
            .O(N__61597),
            .I(N__61538));
    InMux I__14365 (
            .O(N__61596),
            .I(N__61538));
    InMux I__14364 (
            .O(N__61595),
            .I(N__61531));
    InMux I__14363 (
            .O(N__61594),
            .I(N__61531));
    InMux I__14362 (
            .O(N__61593),
            .I(N__61531));
    Span4Mux_v I__14361 (
            .O(N__61584),
            .I(N__61522));
    Span4Mux_h I__14360 (
            .O(N__61577),
            .I(N__61522));
    Span4Mux_v I__14359 (
            .O(N__61572),
            .I(N__61522));
    Span4Mux_v I__14358 (
            .O(N__61567),
            .I(N__61522));
    Sp12to4 I__14357 (
            .O(N__61564),
            .I(N__61519));
    LocalMux I__14356 (
            .O(N__61561),
            .I(N__61516));
    InMux I__14355 (
            .O(N__61560),
            .I(N__61513));
    Span4Mux_h I__14354 (
            .O(N__61553),
            .I(N__61510));
    InMux I__14353 (
            .O(N__61552),
            .I(N__61501));
    InMux I__14352 (
            .O(N__61551),
            .I(N__61501));
    InMux I__14351 (
            .O(N__61550),
            .I(N__61501));
    InMux I__14350 (
            .O(N__61549),
            .I(N__61501));
    InMux I__14349 (
            .O(N__61546),
            .I(N__61498));
    LocalMux I__14348 (
            .O(N__61543),
            .I(N__61485));
    LocalMux I__14347 (
            .O(N__61538),
            .I(N__61485));
    LocalMux I__14346 (
            .O(N__61531),
            .I(N__61485));
    Sp12to4 I__14345 (
            .O(N__61522),
            .I(N__61485));
    Span12Mux_s7_h I__14344 (
            .O(N__61519),
            .I(N__61485));
    Sp12to4 I__14343 (
            .O(N__61516),
            .I(N__61485));
    LocalMux I__14342 (
            .O(N__61513),
            .I(N__61478));
    Span4Mux_h I__14341 (
            .O(N__61510),
            .I(N__61478));
    LocalMux I__14340 (
            .O(N__61501),
            .I(N__61478));
    LocalMux I__14339 (
            .O(N__61498),
            .I(N__61475));
    Span12Mux_h I__14338 (
            .O(N__61485),
            .I(N__61472));
    Sp12to4 I__14337 (
            .O(N__61478),
            .I(N__61469));
    Span12Mux_h I__14336 (
            .O(N__61475),
            .I(N__61466));
    Span12Mux_v I__14335 (
            .O(N__61472),
            .I(N__61461));
    Span12Mux_v I__14334 (
            .O(N__61469),
            .I(N__61461));
    Odrv12 I__14333 (
            .O(N__61466),
            .I(\c0.n19098 ));
    Odrv12 I__14332 (
            .O(N__61461),
            .I(\c0.n19098 ));
    InMux I__14331 (
            .O(N__61456),
            .I(N__61450));
    InMux I__14330 (
            .O(N__61455),
            .I(N__61443));
    InMux I__14329 (
            .O(N__61454),
            .I(N__61443));
    InMux I__14328 (
            .O(N__61453),
            .I(N__61440));
    LocalMux I__14327 (
            .O(N__61450),
            .I(N__61437));
    CascadeMux I__14326 (
            .O(N__61449),
            .I(N__61434));
    InMux I__14325 (
            .O(N__61448),
            .I(N__61431));
    LocalMux I__14324 (
            .O(N__61443),
            .I(N__61425));
    LocalMux I__14323 (
            .O(N__61440),
            .I(N__61425));
    Span4Mux_h I__14322 (
            .O(N__61437),
            .I(N__61421));
    InMux I__14321 (
            .O(N__61434),
            .I(N__61418));
    LocalMux I__14320 (
            .O(N__61431),
            .I(N__61415));
    InMux I__14319 (
            .O(N__61430),
            .I(N__61412));
    Span4Mux_v I__14318 (
            .O(N__61425),
            .I(N__61409));
    CascadeMux I__14317 (
            .O(N__61424),
            .I(N__61404));
    Span4Mux_v I__14316 (
            .O(N__61421),
            .I(N__61401));
    LocalMux I__14315 (
            .O(N__61418),
            .I(N__61398));
    Span4Mux_v I__14314 (
            .O(N__61415),
            .I(N__61395));
    LocalMux I__14313 (
            .O(N__61412),
            .I(N__61392));
    Span4Mux_v I__14312 (
            .O(N__61409),
            .I(N__61389));
    InMux I__14311 (
            .O(N__61408),
            .I(N__61384));
    InMux I__14310 (
            .O(N__61407),
            .I(N__61384));
    InMux I__14309 (
            .O(N__61404),
            .I(N__61381));
    Sp12to4 I__14308 (
            .O(N__61401),
            .I(N__61378));
    Span4Mux_v I__14307 (
            .O(N__61398),
            .I(N__61373));
    Span4Mux_v I__14306 (
            .O(N__61395),
            .I(N__61373));
    Span4Mux_v I__14305 (
            .O(N__61392),
            .I(N__61368));
    Span4Mux_h I__14304 (
            .O(N__61389),
            .I(N__61368));
    LocalMux I__14303 (
            .O(N__61384),
            .I(N__61361));
    LocalMux I__14302 (
            .O(N__61381),
            .I(N__61361));
    Span12Mux_v I__14301 (
            .O(N__61378),
            .I(N__61361));
    Sp12to4 I__14300 (
            .O(N__61373),
            .I(N__61354));
    Sp12to4 I__14299 (
            .O(N__61368),
            .I(N__61354));
    Span12Mux_v I__14298 (
            .O(N__61361),
            .I(N__61354));
    Odrv12 I__14297 (
            .O(N__61354),
            .I(\c0.n9_adj_3251 ));
    InMux I__14296 (
            .O(N__61351),
            .I(N__61348));
    LocalMux I__14295 (
            .O(N__61348),
            .I(N__61342));
    InMux I__14294 (
            .O(N__61347),
            .I(N__61337));
    InMux I__14293 (
            .O(N__61346),
            .I(N__61337));
    CascadeMux I__14292 (
            .O(N__61345),
            .I(N__61334));
    Span4Mux_h I__14291 (
            .O(N__61342),
            .I(N__61331));
    LocalMux I__14290 (
            .O(N__61337),
            .I(N__61328));
    InMux I__14289 (
            .O(N__61334),
            .I(N__61323));
    Span4Mux_h I__14288 (
            .O(N__61331),
            .I(N__61318));
    Span4Mux_v I__14287 (
            .O(N__61328),
            .I(N__61318));
    InMux I__14286 (
            .O(N__61327),
            .I(N__61313));
    InMux I__14285 (
            .O(N__61326),
            .I(N__61313));
    LocalMux I__14284 (
            .O(N__61323),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__14283 (
            .O(N__61318),
            .I(\c0.data_in_frame_3_4 ));
    LocalMux I__14282 (
            .O(N__61313),
            .I(\c0.data_in_frame_3_4 ));
    InMux I__14281 (
            .O(N__61306),
            .I(N__61303));
    LocalMux I__14280 (
            .O(N__61303),
            .I(\c0.n12_adj_2998 ));
    InMux I__14279 (
            .O(N__61300),
            .I(N__61297));
    LocalMux I__14278 (
            .O(N__61297),
            .I(N__61294));
    Span4Mux_h I__14277 (
            .O(N__61294),
            .I(N__61291));
    Span4Mux_h I__14276 (
            .O(N__61291),
            .I(N__61288));
    Odrv4 I__14275 (
            .O(N__61288),
            .I(\c0.n19176 ));
    InMux I__14274 (
            .O(N__61285),
            .I(N__61281));
    InMux I__14273 (
            .O(N__61284),
            .I(N__61278));
    LocalMux I__14272 (
            .O(N__61281),
            .I(N__61275));
    LocalMux I__14271 (
            .O(N__61278),
            .I(N__61272));
    Span4Mux_h I__14270 (
            .O(N__61275),
            .I(N__61269));
    Span12Mux_v I__14269 (
            .O(N__61272),
            .I(N__61266));
    Odrv4 I__14268 (
            .O(N__61269),
            .I(\c0.n11953 ));
    Odrv12 I__14267 (
            .O(N__61266),
            .I(\c0.n11953 ));
    InMux I__14266 (
            .O(N__61261),
            .I(N__61258));
    LocalMux I__14265 (
            .O(N__61258),
            .I(N__61255));
    Span4Mux_v I__14264 (
            .O(N__61255),
            .I(N__61251));
    InMux I__14263 (
            .O(N__61254),
            .I(N__61248));
    Sp12to4 I__14262 (
            .O(N__61251),
            .I(N__61241));
    LocalMux I__14261 (
            .O(N__61248),
            .I(N__61241));
    InMux I__14260 (
            .O(N__61247),
            .I(N__61236));
    InMux I__14259 (
            .O(N__61246),
            .I(N__61236));
    Odrv12 I__14258 (
            .O(N__61241),
            .I(\c0.data_in_frame_5_2 ));
    LocalMux I__14257 (
            .O(N__61236),
            .I(\c0.data_in_frame_5_2 ));
    InMux I__14256 (
            .O(N__61231),
            .I(N__61228));
    LocalMux I__14255 (
            .O(N__61228),
            .I(N__61222));
    InMux I__14254 (
            .O(N__61227),
            .I(N__61219));
    InMux I__14253 (
            .O(N__61226),
            .I(N__61216));
    InMux I__14252 (
            .O(N__61225),
            .I(N__61213));
    Span4Mux_v I__14251 (
            .O(N__61222),
            .I(N__61209));
    LocalMux I__14250 (
            .O(N__61219),
            .I(N__61206));
    LocalMux I__14249 (
            .O(N__61216),
            .I(N__61202));
    LocalMux I__14248 (
            .O(N__61213),
            .I(N__61199));
    InMux I__14247 (
            .O(N__61212),
            .I(N__61190));
    Span4Mux_h I__14246 (
            .O(N__61209),
            .I(N__61187));
    Span4Mux_h I__14245 (
            .O(N__61206),
            .I(N__61184));
    InMux I__14244 (
            .O(N__61205),
            .I(N__61181));
    Span4Mux_h I__14243 (
            .O(N__61202),
            .I(N__61176));
    Span4Mux_h I__14242 (
            .O(N__61199),
            .I(N__61176));
    InMux I__14241 (
            .O(N__61198),
            .I(N__61173));
    InMux I__14240 (
            .O(N__61197),
            .I(N__61170));
    InMux I__14239 (
            .O(N__61196),
            .I(N__61163));
    InMux I__14238 (
            .O(N__61195),
            .I(N__61163));
    InMux I__14237 (
            .O(N__61194),
            .I(N__61163));
    InMux I__14236 (
            .O(N__61193),
            .I(N__61160));
    LocalMux I__14235 (
            .O(N__61190),
            .I(data_in_frame_1_3));
    Odrv4 I__14234 (
            .O(N__61187),
            .I(data_in_frame_1_3));
    Odrv4 I__14233 (
            .O(N__61184),
            .I(data_in_frame_1_3));
    LocalMux I__14232 (
            .O(N__61181),
            .I(data_in_frame_1_3));
    Odrv4 I__14231 (
            .O(N__61176),
            .I(data_in_frame_1_3));
    LocalMux I__14230 (
            .O(N__61173),
            .I(data_in_frame_1_3));
    LocalMux I__14229 (
            .O(N__61170),
            .I(data_in_frame_1_3));
    LocalMux I__14228 (
            .O(N__61163),
            .I(data_in_frame_1_3));
    LocalMux I__14227 (
            .O(N__61160),
            .I(data_in_frame_1_3));
    CascadeMux I__14226 (
            .O(N__61141),
            .I(N__61138));
    InMux I__14225 (
            .O(N__61138),
            .I(N__61135));
    LocalMux I__14224 (
            .O(N__61135),
            .I(\c0.n55_adj_3500 ));
    CascadeMux I__14223 (
            .O(N__61132),
            .I(N__61128));
    InMux I__14222 (
            .O(N__61131),
            .I(N__61123));
    InMux I__14221 (
            .O(N__61128),
            .I(N__61119));
    InMux I__14220 (
            .O(N__61127),
            .I(N__61112));
    InMux I__14219 (
            .O(N__61126),
            .I(N__61112));
    LocalMux I__14218 (
            .O(N__61123),
            .I(N__61109));
    InMux I__14217 (
            .O(N__61122),
            .I(N__61106));
    LocalMux I__14216 (
            .O(N__61119),
            .I(N__61103));
    InMux I__14215 (
            .O(N__61118),
            .I(N__61100));
    InMux I__14214 (
            .O(N__61117),
            .I(N__61096));
    LocalMux I__14213 (
            .O(N__61112),
            .I(N__61093));
    Span4Mux_h I__14212 (
            .O(N__61109),
            .I(N__61087));
    LocalMux I__14211 (
            .O(N__61106),
            .I(N__61087));
    Span4Mux_h I__14210 (
            .O(N__61103),
            .I(N__61082));
    LocalMux I__14209 (
            .O(N__61100),
            .I(N__61082));
    CascadeMux I__14208 (
            .O(N__61099),
            .I(N__61074));
    LocalMux I__14207 (
            .O(N__61096),
            .I(N__61070));
    Span4Mux_v I__14206 (
            .O(N__61093),
            .I(N__61067));
    InMux I__14205 (
            .O(N__61092),
            .I(N__61064));
    Span4Mux_v I__14204 (
            .O(N__61087),
            .I(N__61061));
    Span4Mux_h I__14203 (
            .O(N__61082),
            .I(N__61058));
    InMux I__14202 (
            .O(N__61081),
            .I(N__61055));
    InMux I__14201 (
            .O(N__61080),
            .I(N__61048));
    InMux I__14200 (
            .O(N__61079),
            .I(N__61048));
    InMux I__14199 (
            .O(N__61078),
            .I(N__61048));
    InMux I__14198 (
            .O(N__61077),
            .I(N__61045));
    InMux I__14197 (
            .O(N__61074),
            .I(N__61040));
    InMux I__14196 (
            .O(N__61073),
            .I(N__61040));
    Span4Mux_h I__14195 (
            .O(N__61070),
            .I(N__61033));
    Span4Mux_h I__14194 (
            .O(N__61067),
            .I(N__61033));
    LocalMux I__14193 (
            .O(N__61064),
            .I(N__61033));
    Odrv4 I__14192 (
            .O(N__61061),
            .I(data_in_frame_0_2));
    Odrv4 I__14191 (
            .O(N__61058),
            .I(data_in_frame_0_2));
    LocalMux I__14190 (
            .O(N__61055),
            .I(data_in_frame_0_2));
    LocalMux I__14189 (
            .O(N__61048),
            .I(data_in_frame_0_2));
    LocalMux I__14188 (
            .O(N__61045),
            .I(data_in_frame_0_2));
    LocalMux I__14187 (
            .O(N__61040),
            .I(data_in_frame_0_2));
    Odrv4 I__14186 (
            .O(N__61033),
            .I(data_in_frame_0_2));
    InMux I__14185 (
            .O(N__61018),
            .I(N__61015));
    LocalMux I__14184 (
            .O(N__61015),
            .I(\c0.n7 ));
    CascadeMux I__14183 (
            .O(N__61012),
            .I(N__61008));
    CascadeMux I__14182 (
            .O(N__61011),
            .I(N__61005));
    InMux I__14181 (
            .O(N__61008),
            .I(N__61002));
    InMux I__14180 (
            .O(N__61005),
            .I(N__60999));
    LocalMux I__14179 (
            .O(N__61002),
            .I(N__60994));
    LocalMux I__14178 (
            .O(N__60999),
            .I(N__60994));
    Span4Mux_h I__14177 (
            .O(N__60994),
            .I(N__60991));
    Odrv4 I__14176 (
            .O(N__60991),
            .I(\c0.n19241 ));
    CascadeMux I__14175 (
            .O(N__60988),
            .I(N__60984));
    InMux I__14174 (
            .O(N__60987),
            .I(N__60980));
    InMux I__14173 (
            .O(N__60984),
            .I(N__60977));
    CascadeMux I__14172 (
            .O(N__60983),
            .I(N__60973));
    LocalMux I__14171 (
            .O(N__60980),
            .I(N__60970));
    LocalMux I__14170 (
            .O(N__60977),
            .I(N__60967));
    InMux I__14169 (
            .O(N__60976),
            .I(N__60964));
    InMux I__14168 (
            .O(N__60973),
            .I(N__60961));
    Span4Mux_h I__14167 (
            .O(N__60970),
            .I(N__60958));
    Span4Mux_h I__14166 (
            .O(N__60967),
            .I(N__60953));
    LocalMux I__14165 (
            .O(N__60964),
            .I(N__60950));
    LocalMux I__14164 (
            .O(N__60961),
            .I(N__60945));
    Span4Mux_h I__14163 (
            .O(N__60958),
            .I(N__60945));
    InMux I__14162 (
            .O(N__60957),
            .I(N__60940));
    InMux I__14161 (
            .O(N__60956),
            .I(N__60940));
    Odrv4 I__14160 (
            .O(N__60953),
            .I(\c0.data_in_frame_2_4 ));
    Odrv12 I__14159 (
            .O(N__60950),
            .I(\c0.data_in_frame_2_4 ));
    Odrv4 I__14158 (
            .O(N__60945),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__14157 (
            .O(N__60940),
            .I(\c0.data_in_frame_2_4 ));
    InMux I__14156 (
            .O(N__60931),
            .I(N__60928));
    LocalMux I__14155 (
            .O(N__60928),
            .I(N__60923));
    InMux I__14154 (
            .O(N__60927),
            .I(N__60917));
    InMux I__14153 (
            .O(N__60926),
            .I(N__60917));
    Span4Mux_v I__14152 (
            .O(N__60923),
            .I(N__60913));
    InMux I__14151 (
            .O(N__60922),
            .I(N__60910));
    LocalMux I__14150 (
            .O(N__60917),
            .I(N__60902));
    InMux I__14149 (
            .O(N__60916),
            .I(N__60896));
    Span4Mux_h I__14148 (
            .O(N__60913),
            .I(N__60893));
    LocalMux I__14147 (
            .O(N__60910),
            .I(N__60890));
    InMux I__14146 (
            .O(N__60909),
            .I(N__60887));
    InMux I__14145 (
            .O(N__60908),
            .I(N__60884));
    InMux I__14144 (
            .O(N__60907),
            .I(N__60881));
    InMux I__14143 (
            .O(N__60906),
            .I(N__60876));
    InMux I__14142 (
            .O(N__60905),
            .I(N__60876));
    Span4Mux_h I__14141 (
            .O(N__60902),
            .I(N__60873));
    InMux I__14140 (
            .O(N__60901),
            .I(N__60868));
    InMux I__14139 (
            .O(N__60900),
            .I(N__60868));
    InMux I__14138 (
            .O(N__60899),
            .I(N__60865));
    LocalMux I__14137 (
            .O(N__60896),
            .I(data_in_frame_1_4));
    Odrv4 I__14136 (
            .O(N__60893),
            .I(data_in_frame_1_4));
    Odrv4 I__14135 (
            .O(N__60890),
            .I(data_in_frame_1_4));
    LocalMux I__14134 (
            .O(N__60887),
            .I(data_in_frame_1_4));
    LocalMux I__14133 (
            .O(N__60884),
            .I(data_in_frame_1_4));
    LocalMux I__14132 (
            .O(N__60881),
            .I(data_in_frame_1_4));
    LocalMux I__14131 (
            .O(N__60876),
            .I(data_in_frame_1_4));
    Odrv4 I__14130 (
            .O(N__60873),
            .I(data_in_frame_1_4));
    LocalMux I__14129 (
            .O(N__60868),
            .I(data_in_frame_1_4));
    LocalMux I__14128 (
            .O(N__60865),
            .I(data_in_frame_1_4));
    InMux I__14127 (
            .O(N__60844),
            .I(N__60839));
    InMux I__14126 (
            .O(N__60843),
            .I(N__60836));
    InMux I__14125 (
            .O(N__60842),
            .I(N__60833));
    LocalMux I__14124 (
            .O(N__60839),
            .I(N__60830));
    LocalMux I__14123 (
            .O(N__60836),
            .I(N__60826));
    LocalMux I__14122 (
            .O(N__60833),
            .I(N__60823));
    Span12Mux_h I__14121 (
            .O(N__60830),
            .I(N__60820));
    InMux I__14120 (
            .O(N__60829),
            .I(N__60817));
    Span4Mux_v I__14119 (
            .O(N__60826),
            .I(N__60814));
    Span4Mux_h I__14118 (
            .O(N__60823),
            .I(N__60811));
    Span12Mux_v I__14117 (
            .O(N__60820),
            .I(N__60808));
    LocalMux I__14116 (
            .O(N__60817),
            .I(N__60805));
    Span4Mux_v I__14115 (
            .O(N__60814),
            .I(N__60802));
    Odrv4 I__14114 (
            .O(N__60811),
            .I(\c0.n11833 ));
    Odrv12 I__14113 (
            .O(N__60808),
            .I(\c0.n11833 ));
    Odrv4 I__14112 (
            .O(N__60805),
            .I(\c0.n11833 ));
    Odrv4 I__14111 (
            .O(N__60802),
            .I(\c0.n11833 ));
    InMux I__14110 (
            .O(N__60793),
            .I(N__60788));
    InMux I__14109 (
            .O(N__60792),
            .I(N__60785));
    InMux I__14108 (
            .O(N__60791),
            .I(N__60782));
    LocalMux I__14107 (
            .O(N__60788),
            .I(N__60779));
    LocalMux I__14106 (
            .O(N__60785),
            .I(N__60775));
    LocalMux I__14105 (
            .O(N__60782),
            .I(N__60772));
    Span4Mux_v I__14104 (
            .O(N__60779),
            .I(N__60768));
    InMux I__14103 (
            .O(N__60778),
            .I(N__60765));
    Span4Mux_h I__14102 (
            .O(N__60775),
            .I(N__60762));
    Span4Mux_v I__14101 (
            .O(N__60772),
            .I(N__60759));
    InMux I__14100 (
            .O(N__60771),
            .I(N__60756));
    Odrv4 I__14099 (
            .O(N__60768),
            .I(\c0.n19456 ));
    LocalMux I__14098 (
            .O(N__60765),
            .I(\c0.n19456 ));
    Odrv4 I__14097 (
            .O(N__60762),
            .I(\c0.n19456 ));
    Odrv4 I__14096 (
            .O(N__60759),
            .I(\c0.n19456 ));
    LocalMux I__14095 (
            .O(N__60756),
            .I(\c0.n19456 ));
    InMux I__14094 (
            .O(N__60745),
            .I(N__60742));
    LocalMux I__14093 (
            .O(N__60742),
            .I(N__60739));
    Span4Mux_v I__14092 (
            .O(N__60739),
            .I(N__60736));
    Odrv4 I__14091 (
            .O(N__60736),
            .I(\c0.n5595 ));
    InMux I__14090 (
            .O(N__60733),
            .I(N__60730));
    LocalMux I__14089 (
            .O(N__60730),
            .I(N__60726));
    InMux I__14088 (
            .O(N__60729),
            .I(N__60723));
    Span4Mux_v I__14087 (
            .O(N__60726),
            .I(N__60718));
    LocalMux I__14086 (
            .O(N__60723),
            .I(N__60718));
    Span4Mux_h I__14085 (
            .O(N__60718),
            .I(N__60714));
    InMux I__14084 (
            .O(N__60717),
            .I(N__60711));
    Span4Mux_v I__14083 (
            .O(N__60714),
            .I(N__60704));
    LocalMux I__14082 (
            .O(N__60711),
            .I(N__60704));
    InMux I__14081 (
            .O(N__60710),
            .I(N__60699));
    InMux I__14080 (
            .O(N__60709),
            .I(N__60699));
    Span4Mux_h I__14079 (
            .O(N__60704),
            .I(N__60696));
    LocalMux I__14078 (
            .O(N__60699),
            .I(N__60683));
    Span4Mux_v I__14077 (
            .O(N__60696),
            .I(N__60680));
    InMux I__14076 (
            .O(N__60695),
            .I(N__60677));
    InMux I__14075 (
            .O(N__60694),
            .I(N__60668));
    InMux I__14074 (
            .O(N__60693),
            .I(N__60668));
    InMux I__14073 (
            .O(N__60692),
            .I(N__60668));
    InMux I__14072 (
            .O(N__60691),
            .I(N__60668));
    InMux I__14071 (
            .O(N__60690),
            .I(N__60663));
    InMux I__14070 (
            .O(N__60689),
            .I(N__60663));
    InMux I__14069 (
            .O(N__60688),
            .I(N__60660));
    InMux I__14068 (
            .O(N__60687),
            .I(N__60655));
    InMux I__14067 (
            .O(N__60686),
            .I(N__60655));
    Span4Mux_v I__14066 (
            .O(N__60683),
            .I(N__60647));
    Span4Mux_v I__14065 (
            .O(N__60680),
            .I(N__60644));
    LocalMux I__14064 (
            .O(N__60677),
            .I(N__60641));
    LocalMux I__14063 (
            .O(N__60668),
            .I(N__60636));
    LocalMux I__14062 (
            .O(N__60663),
            .I(N__60636));
    LocalMux I__14061 (
            .O(N__60660),
            .I(N__60629));
    LocalMux I__14060 (
            .O(N__60655),
            .I(N__60626));
    InMux I__14059 (
            .O(N__60654),
            .I(N__60621));
    InMux I__14058 (
            .O(N__60653),
            .I(N__60621));
    InMux I__14057 (
            .O(N__60652),
            .I(N__60612));
    InMux I__14056 (
            .O(N__60651),
            .I(N__60612));
    InMux I__14055 (
            .O(N__60650),
            .I(N__60609));
    Sp12to4 I__14054 (
            .O(N__60647),
            .I(N__60606));
    Span4Mux_v I__14053 (
            .O(N__60644),
            .I(N__60603));
    Span4Mux_v I__14052 (
            .O(N__60641),
            .I(N__60600));
    Span4Mux_v I__14051 (
            .O(N__60636),
            .I(N__60597));
    InMux I__14050 (
            .O(N__60635),
            .I(N__60592));
    InMux I__14049 (
            .O(N__60634),
            .I(N__60592));
    InMux I__14048 (
            .O(N__60633),
            .I(N__60589));
    InMux I__14047 (
            .O(N__60632),
            .I(N__60586));
    Span4Mux_v I__14046 (
            .O(N__60629),
            .I(N__60576));
    Span4Mux_h I__14045 (
            .O(N__60626),
            .I(N__60576));
    LocalMux I__14044 (
            .O(N__60621),
            .I(N__60576));
    InMux I__14043 (
            .O(N__60620),
            .I(N__60567));
    InMux I__14042 (
            .O(N__60619),
            .I(N__60567));
    InMux I__14041 (
            .O(N__60618),
            .I(N__60567));
    InMux I__14040 (
            .O(N__60617),
            .I(N__60567));
    LocalMux I__14039 (
            .O(N__60612),
            .I(N__60560));
    LocalMux I__14038 (
            .O(N__60609),
            .I(N__60560));
    Span12Mux_h I__14037 (
            .O(N__60606),
            .I(N__60560));
    Span4Mux_v I__14036 (
            .O(N__60603),
            .I(N__60555));
    Span4Mux_h I__14035 (
            .O(N__60600),
            .I(N__60555));
    Span4Mux_v I__14034 (
            .O(N__60597),
            .I(N__60552));
    LocalMux I__14033 (
            .O(N__60592),
            .I(N__60549));
    LocalMux I__14032 (
            .O(N__60589),
            .I(N__60546));
    LocalMux I__14031 (
            .O(N__60586),
            .I(N__60543));
    InMux I__14030 (
            .O(N__60585),
            .I(N__60538));
    InMux I__14029 (
            .O(N__60584),
            .I(N__60538));
    InMux I__14028 (
            .O(N__60583),
            .I(N__60535));
    Sp12to4 I__14027 (
            .O(N__60576),
            .I(N__60528));
    LocalMux I__14026 (
            .O(N__60567),
            .I(N__60528));
    Span12Mux_v I__14025 (
            .O(N__60560),
            .I(N__60528));
    Odrv4 I__14024 (
            .O(N__60555),
            .I(n2108));
    Odrv4 I__14023 (
            .O(N__60552),
            .I(n2108));
    Odrv12 I__14022 (
            .O(N__60549),
            .I(n2108));
    Odrv4 I__14021 (
            .O(N__60546),
            .I(n2108));
    Odrv4 I__14020 (
            .O(N__60543),
            .I(n2108));
    LocalMux I__14019 (
            .O(N__60538),
            .I(n2108));
    LocalMux I__14018 (
            .O(N__60535),
            .I(n2108));
    Odrv12 I__14017 (
            .O(N__60528),
            .I(n2108));
    SRMux I__14016 (
            .O(N__60511),
            .I(N__60508));
    LocalMux I__14015 (
            .O(N__60508),
            .I(N__60505));
    Span4Mux_h I__14014 (
            .O(N__60505),
            .I(N__60502));
    Span4Mux_h I__14013 (
            .O(N__60502),
            .I(N__60499));
    Span4Mux_h I__14012 (
            .O(N__60499),
            .I(N__60496));
    Odrv4 I__14011 (
            .O(N__60496),
            .I(\c0.n6_adj_3140 ));
    CascadeMux I__14010 (
            .O(N__60493),
            .I(N__60489));
    InMux I__14009 (
            .O(N__60492),
            .I(N__60482));
    InMux I__14008 (
            .O(N__60489),
            .I(N__60482));
    InMux I__14007 (
            .O(N__60488),
            .I(N__60479));
    InMux I__14006 (
            .O(N__60487),
            .I(N__60475));
    LocalMux I__14005 (
            .O(N__60482),
            .I(N__60472));
    LocalMux I__14004 (
            .O(N__60479),
            .I(N__60469));
    InMux I__14003 (
            .O(N__60478),
            .I(N__60466));
    LocalMux I__14002 (
            .O(N__60475),
            .I(N__60461));
    Span4Mux_h I__14001 (
            .O(N__60472),
            .I(N__60461));
    Span4Mux_h I__14000 (
            .O(N__60469),
            .I(N__60458));
    LocalMux I__13999 (
            .O(N__60466),
            .I(\c0.data_in_frame_6_0 ));
    Odrv4 I__13998 (
            .O(N__60461),
            .I(\c0.data_in_frame_6_0 ));
    Odrv4 I__13997 (
            .O(N__60458),
            .I(\c0.data_in_frame_6_0 ));
    InMux I__13996 (
            .O(N__60451),
            .I(N__60445));
    InMux I__13995 (
            .O(N__60450),
            .I(N__60442));
    CascadeMux I__13994 (
            .O(N__60449),
            .I(N__60439));
    InMux I__13993 (
            .O(N__60448),
            .I(N__60436));
    LocalMux I__13992 (
            .O(N__60445),
            .I(N__60433));
    LocalMux I__13991 (
            .O(N__60442),
            .I(N__60430));
    InMux I__13990 (
            .O(N__60439),
            .I(N__60427));
    LocalMux I__13989 (
            .O(N__60436),
            .I(N__60422));
    Span4Mux_h I__13988 (
            .O(N__60433),
            .I(N__60422));
    Span4Mux_h I__13987 (
            .O(N__60430),
            .I(N__60419));
    LocalMux I__13986 (
            .O(N__60427),
            .I(\c0.data_in_frame_6_2 ));
    Odrv4 I__13985 (
            .O(N__60422),
            .I(\c0.data_in_frame_6_2 ));
    Odrv4 I__13984 (
            .O(N__60419),
            .I(\c0.data_in_frame_6_2 ));
    InMux I__13983 (
            .O(N__60412),
            .I(N__60408));
    InMux I__13982 (
            .O(N__60411),
            .I(N__60405));
    LocalMux I__13981 (
            .O(N__60408),
            .I(N__60402));
    LocalMux I__13980 (
            .O(N__60405),
            .I(N__60399));
    Span4Mux_v I__13979 (
            .O(N__60402),
            .I(N__60395));
    Span4Mux_h I__13978 (
            .O(N__60399),
            .I(N__60392));
    InMux I__13977 (
            .O(N__60398),
            .I(N__60385));
    Span4Mux_h I__13976 (
            .O(N__60395),
            .I(N__60382));
    Span4Mux_h I__13975 (
            .O(N__60392),
            .I(N__60379));
    InMux I__13974 (
            .O(N__60391),
            .I(N__60372));
    InMux I__13973 (
            .O(N__60390),
            .I(N__60372));
    InMux I__13972 (
            .O(N__60389),
            .I(N__60372));
    InMux I__13971 (
            .O(N__60388),
            .I(N__60369));
    LocalMux I__13970 (
            .O(N__60385),
            .I(data_in_frame_1_2));
    Odrv4 I__13969 (
            .O(N__60382),
            .I(data_in_frame_1_2));
    Odrv4 I__13968 (
            .O(N__60379),
            .I(data_in_frame_1_2));
    LocalMux I__13967 (
            .O(N__60372),
            .I(data_in_frame_1_2));
    LocalMux I__13966 (
            .O(N__60369),
            .I(data_in_frame_1_2));
    CascadeMux I__13965 (
            .O(N__60358),
            .I(N__60355));
    InMux I__13964 (
            .O(N__60355),
            .I(N__60347));
    InMux I__13963 (
            .O(N__60354),
            .I(N__60347));
    InMux I__13962 (
            .O(N__60353),
            .I(N__60343));
    InMux I__13961 (
            .O(N__60352),
            .I(N__60340));
    LocalMux I__13960 (
            .O(N__60347),
            .I(N__60337));
    InMux I__13959 (
            .O(N__60346),
            .I(N__60333));
    LocalMux I__13958 (
            .O(N__60343),
            .I(N__60330));
    LocalMux I__13957 (
            .O(N__60340),
            .I(N__60326));
    Span4Mux_v I__13956 (
            .O(N__60337),
            .I(N__60323));
    InMux I__13955 (
            .O(N__60336),
            .I(N__60320));
    LocalMux I__13954 (
            .O(N__60333),
            .I(N__60316));
    Sp12to4 I__13953 (
            .O(N__60330),
            .I(N__60313));
    CascadeMux I__13952 (
            .O(N__60329),
            .I(N__60310));
    Span4Mux_v I__13951 (
            .O(N__60326),
            .I(N__60302));
    Span4Mux_h I__13950 (
            .O(N__60323),
            .I(N__60302));
    LocalMux I__13949 (
            .O(N__60320),
            .I(N__60302));
    InMux I__13948 (
            .O(N__60319),
            .I(N__60299));
    Span4Mux_v I__13947 (
            .O(N__60316),
            .I(N__60296));
    Span12Mux_s10_v I__13946 (
            .O(N__60313),
            .I(N__60293));
    InMux I__13945 (
            .O(N__60310),
            .I(N__60288));
    InMux I__13944 (
            .O(N__60309),
            .I(N__60288));
    Span4Mux_h I__13943 (
            .O(N__60302),
            .I(N__60281));
    LocalMux I__13942 (
            .O(N__60299),
            .I(N__60281));
    Span4Mux_v I__13941 (
            .O(N__60296),
            .I(N__60281));
    Odrv12 I__13940 (
            .O(N__60293),
            .I(\c0.n9_adj_3101 ));
    LocalMux I__13939 (
            .O(N__60288),
            .I(\c0.n9_adj_3101 ));
    Odrv4 I__13938 (
            .O(N__60281),
            .I(\c0.n9_adj_3101 ));
    InMux I__13937 (
            .O(N__60274),
            .I(N__60269));
    InMux I__13936 (
            .O(N__60273),
            .I(N__60265));
    InMux I__13935 (
            .O(N__60272),
            .I(N__60260));
    LocalMux I__13934 (
            .O(N__60269),
            .I(N__60257));
    InMux I__13933 (
            .O(N__60268),
            .I(N__60253));
    LocalMux I__13932 (
            .O(N__60265),
            .I(N__60249));
    CascadeMux I__13931 (
            .O(N__60264),
            .I(N__60246));
    CascadeMux I__13930 (
            .O(N__60263),
            .I(N__60243));
    LocalMux I__13929 (
            .O(N__60260),
            .I(N__60239));
    Span4Mux_v I__13928 (
            .O(N__60257),
            .I(N__60236));
    InMux I__13927 (
            .O(N__60256),
            .I(N__60232));
    LocalMux I__13926 (
            .O(N__60253),
            .I(N__60229));
    InMux I__13925 (
            .O(N__60252),
            .I(N__60226));
    Span4Mux_v I__13924 (
            .O(N__60249),
            .I(N__60223));
    InMux I__13923 (
            .O(N__60246),
            .I(N__60220));
    InMux I__13922 (
            .O(N__60243),
            .I(N__60215));
    InMux I__13921 (
            .O(N__60242),
            .I(N__60215));
    Span4Mux_v I__13920 (
            .O(N__60239),
            .I(N__60212));
    Span4Mux_v I__13919 (
            .O(N__60236),
            .I(N__60209));
    CascadeMux I__13918 (
            .O(N__60235),
            .I(N__60205));
    LocalMux I__13917 (
            .O(N__60232),
            .I(N__60201));
    Span4Mux_v I__13916 (
            .O(N__60229),
            .I(N__60198));
    LocalMux I__13915 (
            .O(N__60226),
            .I(N__60195));
    Span4Mux_h I__13914 (
            .O(N__60223),
            .I(N__60192));
    LocalMux I__13913 (
            .O(N__60220),
            .I(N__60189));
    LocalMux I__13912 (
            .O(N__60215),
            .I(N__60186));
    Span4Mux_v I__13911 (
            .O(N__60212),
            .I(N__60183));
    Span4Mux_h I__13910 (
            .O(N__60209),
            .I(N__60180));
    InMux I__13909 (
            .O(N__60208),
            .I(N__60177));
    InMux I__13908 (
            .O(N__60205),
            .I(N__60174));
    InMux I__13907 (
            .O(N__60204),
            .I(N__60171));
    Span4Mux_v I__13906 (
            .O(N__60201),
            .I(N__60168));
    Span4Mux_h I__13905 (
            .O(N__60198),
            .I(N__60163));
    Span4Mux_v I__13904 (
            .O(N__60195),
            .I(N__60163));
    Span4Mux_h I__13903 (
            .O(N__60192),
            .I(N__60154));
    Span4Mux_v I__13902 (
            .O(N__60189),
            .I(N__60154));
    Span4Mux_v I__13901 (
            .O(N__60186),
            .I(N__60154));
    Span4Mux_v I__13900 (
            .O(N__60183),
            .I(N__60154));
    Span4Mux_v I__13899 (
            .O(N__60180),
            .I(N__60151));
    LocalMux I__13898 (
            .O(N__60177),
            .I(N__60148));
    LocalMux I__13897 (
            .O(N__60174),
            .I(FRAME_MATCHER_i_0));
    LocalMux I__13896 (
            .O(N__60171),
            .I(FRAME_MATCHER_i_0));
    Odrv4 I__13895 (
            .O(N__60168),
            .I(FRAME_MATCHER_i_0));
    Odrv4 I__13894 (
            .O(N__60163),
            .I(FRAME_MATCHER_i_0));
    Odrv4 I__13893 (
            .O(N__60154),
            .I(FRAME_MATCHER_i_0));
    Odrv4 I__13892 (
            .O(N__60151),
            .I(FRAME_MATCHER_i_0));
    Odrv4 I__13891 (
            .O(N__60148),
            .I(FRAME_MATCHER_i_0));
    CascadeMux I__13890 (
            .O(N__60133),
            .I(N__60129));
    InMux I__13889 (
            .O(N__60132),
            .I(N__60125));
    InMux I__13888 (
            .O(N__60129),
            .I(N__60122));
    InMux I__13887 (
            .O(N__60128),
            .I(N__60118));
    LocalMux I__13886 (
            .O(N__60125),
            .I(N__60112));
    LocalMux I__13885 (
            .O(N__60122),
            .I(N__60109));
    InMux I__13884 (
            .O(N__60121),
            .I(N__60105));
    LocalMux I__13883 (
            .O(N__60118),
            .I(N__60101));
    InMux I__13882 (
            .O(N__60117),
            .I(N__60098));
    InMux I__13881 (
            .O(N__60116),
            .I(N__60095));
    InMux I__13880 (
            .O(N__60115),
            .I(N__60092));
    Span4Mux_h I__13879 (
            .O(N__60112),
            .I(N__60089));
    Span4Mux_v I__13878 (
            .O(N__60109),
            .I(N__60086));
    InMux I__13877 (
            .O(N__60108),
            .I(N__60083));
    LocalMux I__13876 (
            .O(N__60105),
            .I(N__60080));
    InMux I__13875 (
            .O(N__60104),
            .I(N__60077));
    Span4Mux_h I__13874 (
            .O(N__60101),
            .I(N__60072));
    LocalMux I__13873 (
            .O(N__60098),
            .I(N__60072));
    LocalMux I__13872 (
            .O(N__60095),
            .I(N__60069));
    LocalMux I__13871 (
            .O(N__60092),
            .I(N__60064));
    Span4Mux_h I__13870 (
            .O(N__60089),
            .I(N__60064));
    Sp12to4 I__13869 (
            .O(N__60086),
            .I(N__60061));
    LocalMux I__13868 (
            .O(N__60083),
            .I(N__60058));
    Span4Mux_v I__13867 (
            .O(N__60080),
            .I(N__60053));
    LocalMux I__13866 (
            .O(N__60077),
            .I(N__60053));
    Span4Mux_v I__13865 (
            .O(N__60072),
            .I(N__60050));
    Span4Mux_h I__13864 (
            .O(N__60069),
            .I(N__60042));
    Span4Mux_v I__13863 (
            .O(N__60064),
            .I(N__60042));
    Span12Mux_h I__13862 (
            .O(N__60061),
            .I(N__60038));
    Span4Mux_h I__13861 (
            .O(N__60058),
            .I(N__60035));
    Span4Mux_v I__13860 (
            .O(N__60053),
            .I(N__60032));
    Sp12to4 I__13859 (
            .O(N__60050),
            .I(N__60029));
    InMux I__13858 (
            .O(N__60049),
            .I(N__60022));
    InMux I__13857 (
            .O(N__60048),
            .I(N__60022));
    InMux I__13856 (
            .O(N__60047),
            .I(N__60022));
    Sp12to4 I__13855 (
            .O(N__60042),
            .I(N__60019));
    InMux I__13854 (
            .O(N__60041),
            .I(N__60016));
    Odrv12 I__13853 (
            .O(N__60038),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__13852 (
            .O(N__60035),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__13851 (
            .O(N__60032),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv12 I__13850 (
            .O(N__60029),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__13849 (
            .O(N__60022),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv12 I__13848 (
            .O(N__60019),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__13847 (
            .O(N__60016),
            .I(\c0.FRAME_MATCHER_i_1 ));
    InMux I__13846 (
            .O(N__60001),
            .I(N__59997));
    InMux I__13845 (
            .O(N__60000),
            .I(N__59993));
    LocalMux I__13844 (
            .O(N__59997),
            .I(N__59989));
    InMux I__13843 (
            .O(N__59996),
            .I(N__59986));
    LocalMux I__13842 (
            .O(N__59993),
            .I(N__59982));
    InMux I__13841 (
            .O(N__59992),
            .I(N__59979));
    Span4Mux_v I__13840 (
            .O(N__59989),
            .I(N__59972));
    LocalMux I__13839 (
            .O(N__59986),
            .I(N__59972));
    InMux I__13838 (
            .O(N__59985),
            .I(N__59969));
    Span4Mux_h I__13837 (
            .O(N__59982),
            .I(N__59966));
    LocalMux I__13836 (
            .O(N__59979),
            .I(N__59962));
    InMux I__13835 (
            .O(N__59978),
            .I(N__59959));
    InMux I__13834 (
            .O(N__59977),
            .I(N__59956));
    Span4Mux_h I__13833 (
            .O(N__59972),
            .I(N__59951));
    LocalMux I__13832 (
            .O(N__59969),
            .I(N__59951));
    Span4Mux_h I__13831 (
            .O(N__59966),
            .I(N__59948));
    CascadeMux I__13830 (
            .O(N__59965),
            .I(N__59945));
    Span4Mux_v I__13829 (
            .O(N__59962),
            .I(N__59939));
    LocalMux I__13828 (
            .O(N__59959),
            .I(N__59939));
    LocalMux I__13827 (
            .O(N__59956),
            .I(N__59934));
    Span4Mux_h I__13826 (
            .O(N__59951),
            .I(N__59934));
    Span4Mux_v I__13825 (
            .O(N__59948),
            .I(N__59931));
    InMux I__13824 (
            .O(N__59945),
            .I(N__59928));
    CascadeMux I__13823 (
            .O(N__59944),
            .I(N__59924));
    Span4Mux_h I__13822 (
            .O(N__59939),
            .I(N__59914));
    Span4Mux_h I__13821 (
            .O(N__59934),
            .I(N__59914));
    Span4Mux_v I__13820 (
            .O(N__59931),
            .I(N__59914));
    LocalMux I__13819 (
            .O(N__59928),
            .I(N__59911));
    InMux I__13818 (
            .O(N__59927),
            .I(N__59908));
    InMux I__13817 (
            .O(N__59924),
            .I(N__59899));
    InMux I__13816 (
            .O(N__59923),
            .I(N__59899));
    InMux I__13815 (
            .O(N__59922),
            .I(N__59899));
    InMux I__13814 (
            .O(N__59921),
            .I(N__59899));
    Span4Mux_v I__13813 (
            .O(N__59914),
            .I(N__59896));
    Span12Mux_v I__13812 (
            .O(N__59911),
            .I(N__59893));
    LocalMux I__13811 (
            .O(N__59908),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__13810 (
            .O(N__59899),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__13809 (
            .O(N__59896),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv12 I__13808 (
            .O(N__59893),
            .I(\c0.FRAME_MATCHER_i_2 ));
    InMux I__13807 (
            .O(N__59884),
            .I(N__59880));
    InMux I__13806 (
            .O(N__59883),
            .I(N__59877));
    LocalMux I__13805 (
            .O(N__59880),
            .I(N__59870));
    LocalMux I__13804 (
            .O(N__59877),
            .I(N__59870));
    InMux I__13803 (
            .O(N__59876),
            .I(N__59861));
    InMux I__13802 (
            .O(N__59875),
            .I(N__59861));
    Span4Mux_h I__13801 (
            .O(N__59870),
            .I(N__59858));
    InMux I__13800 (
            .O(N__59869),
            .I(N__59855));
    InMux I__13799 (
            .O(N__59868),
            .I(N__59848));
    InMux I__13798 (
            .O(N__59867),
            .I(N__59848));
    InMux I__13797 (
            .O(N__59866),
            .I(N__59848));
    LocalMux I__13796 (
            .O(N__59861),
            .I(N__59845));
    Span4Mux_h I__13795 (
            .O(N__59858),
            .I(N__59842));
    LocalMux I__13794 (
            .O(N__59855),
            .I(n19100));
    LocalMux I__13793 (
            .O(N__59848),
            .I(n19100));
    Odrv12 I__13792 (
            .O(N__59845),
            .I(n19100));
    Odrv4 I__13791 (
            .O(N__59842),
            .I(n19100));
    InMux I__13790 (
            .O(N__59833),
            .I(N__59829));
    InMux I__13789 (
            .O(N__59832),
            .I(N__59825));
    LocalMux I__13788 (
            .O(N__59829),
            .I(N__59822));
    InMux I__13787 (
            .O(N__59828),
            .I(N__59819));
    LocalMux I__13786 (
            .O(N__59825),
            .I(\c0.n17942 ));
    Odrv12 I__13785 (
            .O(N__59822),
            .I(\c0.n17942 ));
    LocalMux I__13784 (
            .O(N__59819),
            .I(\c0.n17942 ));
    CascadeMux I__13783 (
            .O(N__59812),
            .I(\c0.n77_adj_3396_cascade_ ));
    InMux I__13782 (
            .O(N__59809),
            .I(N__59806));
    LocalMux I__13781 (
            .O(N__59806),
            .I(N__59803));
    Span4Mux_h I__13780 (
            .O(N__59803),
            .I(N__59800));
    Span4Mux_v I__13779 (
            .O(N__59800),
            .I(N__59797));
    Odrv4 I__13778 (
            .O(N__59797),
            .I(\c0.n90_adj_3400 ));
    CascadeMux I__13777 (
            .O(N__59794),
            .I(N__59791));
    InMux I__13776 (
            .O(N__59791),
            .I(N__59788));
    LocalMux I__13775 (
            .O(N__59788),
            .I(N__59785));
    Span4Mux_v I__13774 (
            .O(N__59785),
            .I(N__59780));
    CascadeMux I__13773 (
            .O(N__59784),
            .I(N__59776));
    CascadeMux I__13772 (
            .O(N__59783),
            .I(N__59772));
    Span4Mux_h I__13771 (
            .O(N__59780),
            .I(N__59769));
    InMux I__13770 (
            .O(N__59779),
            .I(N__59766));
    InMux I__13769 (
            .O(N__59776),
            .I(N__59763));
    InMux I__13768 (
            .O(N__59775),
            .I(N__59760));
    InMux I__13767 (
            .O(N__59772),
            .I(N__59757));
    Sp12to4 I__13766 (
            .O(N__59769),
            .I(N__59748));
    LocalMux I__13765 (
            .O(N__59766),
            .I(N__59748));
    LocalMux I__13764 (
            .O(N__59763),
            .I(N__59748));
    LocalMux I__13763 (
            .O(N__59760),
            .I(N__59748));
    LocalMux I__13762 (
            .O(N__59757),
            .I(\c0.data_in_frame_25_7 ));
    Odrv12 I__13761 (
            .O(N__59748),
            .I(\c0.data_in_frame_25_7 ));
    InMux I__13760 (
            .O(N__59743),
            .I(N__59739));
    InMux I__13759 (
            .O(N__59742),
            .I(N__59735));
    LocalMux I__13758 (
            .O(N__59739),
            .I(N__59732));
    InMux I__13757 (
            .O(N__59738),
            .I(N__59729));
    LocalMux I__13756 (
            .O(N__59735),
            .I(N__59726));
    Span4Mux_v I__13755 (
            .O(N__59732),
            .I(N__59723));
    LocalMux I__13754 (
            .O(N__59729),
            .I(N__59720));
    Span4Mux_v I__13753 (
            .O(N__59726),
            .I(N__59712));
    Span4Mux_h I__13752 (
            .O(N__59723),
            .I(N__59712));
    Span4Mux_v I__13751 (
            .O(N__59720),
            .I(N__59712));
    InMux I__13750 (
            .O(N__59719),
            .I(N__59709));
    Span4Mux_v I__13749 (
            .O(N__59712),
            .I(N__59706));
    LocalMux I__13748 (
            .O(N__59709),
            .I(\c0.data_in_frame_25_5 ));
    Odrv4 I__13747 (
            .O(N__59706),
            .I(\c0.data_in_frame_25_5 ));
    CascadeMux I__13746 (
            .O(N__59701),
            .I(N__59696));
    InMux I__13745 (
            .O(N__59700),
            .I(N__59693));
    InMux I__13744 (
            .O(N__59699),
            .I(N__59689));
    InMux I__13743 (
            .O(N__59696),
            .I(N__59685));
    LocalMux I__13742 (
            .O(N__59693),
            .I(N__59682));
    CascadeMux I__13741 (
            .O(N__59692),
            .I(N__59679));
    LocalMux I__13740 (
            .O(N__59689),
            .I(N__59676));
    InMux I__13739 (
            .O(N__59688),
            .I(N__59673));
    LocalMux I__13738 (
            .O(N__59685),
            .I(N__59670));
    Span4Mux_v I__13737 (
            .O(N__59682),
            .I(N__59666));
    InMux I__13736 (
            .O(N__59679),
            .I(N__59663));
    Span4Mux_v I__13735 (
            .O(N__59676),
            .I(N__59660));
    LocalMux I__13734 (
            .O(N__59673),
            .I(N__59657));
    Span4Mux_v I__13733 (
            .O(N__59670),
            .I(N__59654));
    CascadeMux I__13732 (
            .O(N__59669),
            .I(N__59651));
    Sp12to4 I__13731 (
            .O(N__59666),
            .I(N__59644));
    LocalMux I__13730 (
            .O(N__59663),
            .I(N__59644));
    Sp12to4 I__13729 (
            .O(N__59660),
            .I(N__59644));
    Span4Mux_v I__13728 (
            .O(N__59657),
            .I(N__59639));
    Span4Mux_h I__13727 (
            .O(N__59654),
            .I(N__59639));
    InMux I__13726 (
            .O(N__59651),
            .I(N__59636));
    Span12Mux_h I__13725 (
            .O(N__59644),
            .I(N__59633));
    Span4Mux_v I__13724 (
            .O(N__59639),
            .I(N__59630));
    LocalMux I__13723 (
            .O(N__59636),
            .I(\c0.data_in_frame_25_4 ));
    Odrv12 I__13722 (
            .O(N__59633),
            .I(\c0.data_in_frame_25_4 ));
    Odrv4 I__13721 (
            .O(N__59630),
            .I(\c0.data_in_frame_25_4 ));
    CascadeMux I__13720 (
            .O(N__59623),
            .I(\c0.n19214_cascade_ ));
    InMux I__13719 (
            .O(N__59620),
            .I(N__59617));
    LocalMux I__13718 (
            .O(N__59617),
            .I(N__59613));
    InMux I__13717 (
            .O(N__59616),
            .I(N__59609));
    Span4Mux_h I__13716 (
            .O(N__59613),
            .I(N__59606));
    InMux I__13715 (
            .O(N__59612),
            .I(N__59603));
    LocalMux I__13714 (
            .O(N__59609),
            .I(data_in_frame_24_5));
    Odrv4 I__13713 (
            .O(N__59606),
            .I(data_in_frame_24_5));
    LocalMux I__13712 (
            .O(N__59603),
            .I(data_in_frame_24_5));
    InMux I__13711 (
            .O(N__59596),
            .I(N__59592));
    InMux I__13710 (
            .O(N__59595),
            .I(N__59589));
    LocalMux I__13709 (
            .O(N__59592),
            .I(N__59585));
    LocalMux I__13708 (
            .O(N__59589),
            .I(N__59582));
    InMux I__13707 (
            .O(N__59588),
            .I(N__59579));
    Span4Mux_v I__13706 (
            .O(N__59585),
            .I(N__59576));
    Span4Mux_v I__13705 (
            .O(N__59582),
            .I(N__59571));
    LocalMux I__13704 (
            .O(N__59579),
            .I(N__59571));
    Span4Mux_h I__13703 (
            .O(N__59576),
            .I(N__59568));
    Span4Mux_h I__13702 (
            .O(N__59571),
            .I(N__59565));
    Odrv4 I__13701 (
            .O(N__59568),
            .I(\c0.n12_adj_3214 ));
    Odrv4 I__13700 (
            .O(N__59565),
            .I(\c0.n12_adj_3214 ));
    InMux I__13699 (
            .O(N__59560),
            .I(N__59557));
    LocalMux I__13698 (
            .O(N__59557),
            .I(N__59553));
    CascadeMux I__13697 (
            .O(N__59556),
            .I(N__59550));
    Span4Mux_h I__13696 (
            .O(N__59553),
            .I(N__59545));
    InMux I__13695 (
            .O(N__59550),
            .I(N__59540));
    InMux I__13694 (
            .O(N__59549),
            .I(N__59540));
    InMux I__13693 (
            .O(N__59548),
            .I(N__59537));
    Odrv4 I__13692 (
            .O(N__59545),
            .I(\c0.data_in_frame_25_6 ));
    LocalMux I__13691 (
            .O(N__59540),
            .I(\c0.data_in_frame_25_6 ));
    LocalMux I__13690 (
            .O(N__59537),
            .I(\c0.data_in_frame_25_6 ));
    InMux I__13689 (
            .O(N__59530),
            .I(N__59527));
    LocalMux I__13688 (
            .O(N__59527),
            .I(N__59524));
    Span4Mux_h I__13687 (
            .O(N__59524),
            .I(N__59521));
    Span4Mux_v I__13686 (
            .O(N__59521),
            .I(N__59518));
    Span4Mux_v I__13685 (
            .O(N__59518),
            .I(N__59515));
    Odrv4 I__13684 (
            .O(N__59515),
            .I(\c0.n5784 ));
    InMux I__13683 (
            .O(N__59512),
            .I(N__59508));
    InMux I__13682 (
            .O(N__59511),
            .I(N__59505));
    LocalMux I__13681 (
            .O(N__59508),
            .I(N__59501));
    LocalMux I__13680 (
            .O(N__59505),
            .I(N__59498));
    InMux I__13679 (
            .O(N__59504),
            .I(N__59495));
    Span4Mux_v I__13678 (
            .O(N__59501),
            .I(N__59488));
    Span4Mux_v I__13677 (
            .O(N__59498),
            .I(N__59488));
    LocalMux I__13676 (
            .O(N__59495),
            .I(N__59488));
    Odrv4 I__13675 (
            .O(N__59488),
            .I(\c0.n18431 ));
    InMux I__13674 (
            .O(N__59485),
            .I(N__59482));
    LocalMux I__13673 (
            .O(N__59482),
            .I(N__59475));
    InMux I__13672 (
            .O(N__59481),
            .I(N__59472));
    InMux I__13671 (
            .O(N__59480),
            .I(N__59469));
    InMux I__13670 (
            .O(N__59479),
            .I(N__59466));
    InMux I__13669 (
            .O(N__59478),
            .I(N__59463));
    Span4Mux_v I__13668 (
            .O(N__59475),
            .I(N__59460));
    LocalMux I__13667 (
            .O(N__59472),
            .I(N__59456));
    LocalMux I__13666 (
            .O(N__59469),
            .I(N__59452));
    LocalMux I__13665 (
            .O(N__59466),
            .I(N__59449));
    LocalMux I__13664 (
            .O(N__59463),
            .I(N__59443));
    Span4Mux_v I__13663 (
            .O(N__59460),
            .I(N__59443));
    InMux I__13662 (
            .O(N__59459),
            .I(N__59440));
    Span4Mux_v I__13661 (
            .O(N__59456),
            .I(N__59436));
    InMux I__13660 (
            .O(N__59455),
            .I(N__59433));
    Span4Mux_h I__13659 (
            .O(N__59452),
            .I(N__59429));
    Span4Mux_v I__13658 (
            .O(N__59449),
            .I(N__59426));
    InMux I__13657 (
            .O(N__59448),
            .I(N__59423));
    Span4Mux_h I__13656 (
            .O(N__59443),
            .I(N__59418));
    LocalMux I__13655 (
            .O(N__59440),
            .I(N__59418));
    InMux I__13654 (
            .O(N__59439),
            .I(N__59415));
    Span4Mux_v I__13653 (
            .O(N__59436),
            .I(N__59412));
    LocalMux I__13652 (
            .O(N__59433),
            .I(N__59409));
    InMux I__13651 (
            .O(N__59432),
            .I(N__59406));
    Span4Mux_v I__13650 (
            .O(N__59429),
            .I(N__59403));
    Span4Mux_h I__13649 (
            .O(N__59426),
            .I(N__59396));
    LocalMux I__13648 (
            .O(N__59423),
            .I(N__59396));
    Span4Mux_v I__13647 (
            .O(N__59418),
            .I(N__59396));
    LocalMux I__13646 (
            .O(N__59415),
            .I(N__59393));
    Odrv4 I__13645 (
            .O(N__59412),
            .I(\c0.n15701 ));
    Odrv4 I__13644 (
            .O(N__59409),
            .I(\c0.n15701 ));
    LocalMux I__13643 (
            .O(N__59406),
            .I(\c0.n15701 ));
    Odrv4 I__13642 (
            .O(N__59403),
            .I(\c0.n15701 ));
    Odrv4 I__13641 (
            .O(N__59396),
            .I(\c0.n15701 ));
    Odrv4 I__13640 (
            .O(N__59393),
            .I(\c0.n15701 ));
    InMux I__13639 (
            .O(N__59380),
            .I(N__59377));
    LocalMux I__13638 (
            .O(N__59377),
            .I(N__59374));
    Span4Mux_v I__13637 (
            .O(N__59374),
            .I(N__59371));
    Span4Mux_h I__13636 (
            .O(N__59371),
            .I(N__59368));
    Span4Mux_v I__13635 (
            .O(N__59368),
            .I(N__59365));
    Span4Mux_h I__13634 (
            .O(N__59365),
            .I(N__59362));
    Odrv4 I__13633 (
            .O(N__59362),
            .I(\c0.n7_adj_3047 ));
    InMux I__13632 (
            .O(N__59359),
            .I(N__59355));
    InMux I__13631 (
            .O(N__59358),
            .I(N__59352));
    LocalMux I__13630 (
            .O(N__59355),
            .I(N__59349));
    LocalMux I__13629 (
            .O(N__59352),
            .I(N__59346));
    Span4Mux_h I__13628 (
            .O(N__59349),
            .I(N__59340));
    Span4Mux_v I__13627 (
            .O(N__59346),
            .I(N__59340));
    InMux I__13626 (
            .O(N__59345),
            .I(N__59337));
    Odrv4 I__13625 (
            .O(N__59340),
            .I(\c0.n20965 ));
    LocalMux I__13624 (
            .O(N__59337),
            .I(\c0.n20965 ));
    InMux I__13623 (
            .O(N__59332),
            .I(N__59329));
    LocalMux I__13622 (
            .O(N__59329),
            .I(N__59326));
    Span4Mux_h I__13621 (
            .O(N__59326),
            .I(N__59321));
    CascadeMux I__13620 (
            .O(N__59325),
            .I(N__59318));
    CascadeMux I__13619 (
            .O(N__59324),
            .I(N__59315));
    Span4Mux_h I__13618 (
            .O(N__59321),
            .I(N__59312));
    InMux I__13617 (
            .O(N__59318),
            .I(N__59307));
    InMux I__13616 (
            .O(N__59315),
            .I(N__59307));
    Odrv4 I__13615 (
            .O(N__59312),
            .I(\c0.data_in_frame_26_0 ));
    LocalMux I__13614 (
            .O(N__59307),
            .I(\c0.data_in_frame_26_0 ));
    InMux I__13613 (
            .O(N__59302),
            .I(N__59297));
    InMux I__13612 (
            .O(N__59301),
            .I(N__59294));
    CascadeMux I__13611 (
            .O(N__59300),
            .I(N__59291));
    LocalMux I__13610 (
            .O(N__59297),
            .I(N__59288));
    LocalMux I__13609 (
            .O(N__59294),
            .I(N__59285));
    InMux I__13608 (
            .O(N__59291),
            .I(N__59282));
    Span4Mux_h I__13607 (
            .O(N__59288),
            .I(N__59279));
    Span4Mux_h I__13606 (
            .O(N__59285),
            .I(N__59276));
    LocalMux I__13605 (
            .O(N__59282),
            .I(N__59269));
    Span4Mux_h I__13604 (
            .O(N__59279),
            .I(N__59269));
    Span4Mux_h I__13603 (
            .O(N__59276),
            .I(N__59266));
    InMux I__13602 (
            .O(N__59275),
            .I(N__59261));
    InMux I__13601 (
            .O(N__59274),
            .I(N__59261));
    Odrv4 I__13600 (
            .O(N__59269),
            .I(\c0.data_in_frame_27_1 ));
    Odrv4 I__13599 (
            .O(N__59266),
            .I(\c0.data_in_frame_27_1 ));
    LocalMux I__13598 (
            .O(N__59261),
            .I(\c0.data_in_frame_27_1 ));
    CascadeMux I__13597 (
            .O(N__59254),
            .I(N__59251));
    InMux I__13596 (
            .O(N__59251),
            .I(N__59247));
    InMux I__13595 (
            .O(N__59250),
            .I(N__59244));
    LocalMux I__13594 (
            .O(N__59247),
            .I(N__59241));
    LocalMux I__13593 (
            .O(N__59244),
            .I(N__59238));
    Span4Mux_h I__13592 (
            .O(N__59241),
            .I(N__59232));
    Span4Mux_h I__13591 (
            .O(N__59238),
            .I(N__59232));
    InMux I__13590 (
            .O(N__59237),
            .I(N__59227));
    Span4Mux_h I__13589 (
            .O(N__59232),
            .I(N__59224));
    InMux I__13588 (
            .O(N__59231),
            .I(N__59219));
    InMux I__13587 (
            .O(N__59230),
            .I(N__59219));
    LocalMux I__13586 (
            .O(N__59227),
            .I(\c0.data_in_frame_27_2 ));
    Odrv4 I__13585 (
            .O(N__59224),
            .I(\c0.data_in_frame_27_2 ));
    LocalMux I__13584 (
            .O(N__59219),
            .I(\c0.data_in_frame_27_2 ));
    InMux I__13583 (
            .O(N__59212),
            .I(N__59208));
    CascadeMux I__13582 (
            .O(N__59211),
            .I(N__59205));
    LocalMux I__13581 (
            .O(N__59208),
            .I(N__59202));
    InMux I__13580 (
            .O(N__59205),
            .I(N__59199));
    Span12Mux_s9_v I__13579 (
            .O(N__59202),
            .I(N__59196));
    LocalMux I__13578 (
            .O(N__59199),
            .I(\c0.data_in_frame_28_2 ));
    Odrv12 I__13577 (
            .O(N__59196),
            .I(\c0.data_in_frame_28_2 ));
    InMux I__13576 (
            .O(N__59191),
            .I(N__59187));
    InMux I__13575 (
            .O(N__59190),
            .I(N__59184));
    LocalMux I__13574 (
            .O(N__59187),
            .I(\c0.n20709 ));
    LocalMux I__13573 (
            .O(N__59184),
            .I(\c0.n20709 ));
    CascadeMux I__13572 (
            .O(N__59179),
            .I(N__59175));
    InMux I__13571 (
            .O(N__59178),
            .I(N__59172));
    InMux I__13570 (
            .O(N__59175),
            .I(N__59169));
    LocalMux I__13569 (
            .O(N__59172),
            .I(N__59166));
    LocalMux I__13568 (
            .O(N__59169),
            .I(N__59162));
    Span4Mux_h I__13567 (
            .O(N__59166),
            .I(N__59159));
    InMux I__13566 (
            .O(N__59165),
            .I(N__59156));
    Odrv4 I__13565 (
            .O(N__59162),
            .I(\c0.n38_adj_3062 ));
    Odrv4 I__13564 (
            .O(N__59159),
            .I(\c0.n38_adj_3062 ));
    LocalMux I__13563 (
            .O(N__59156),
            .I(\c0.n38_adj_3062 ));
    CascadeMux I__13562 (
            .O(N__59149),
            .I(N__59146));
    InMux I__13561 (
            .O(N__59146),
            .I(N__59143));
    LocalMux I__13560 (
            .O(N__59143),
            .I(N__59140));
    Odrv12 I__13559 (
            .O(N__59140),
            .I(\c0.n83_adj_3442 ));
    CascadeMux I__13558 (
            .O(N__59137),
            .I(N__59134));
    InMux I__13557 (
            .O(N__59134),
            .I(N__59130));
    InMux I__13556 (
            .O(N__59133),
            .I(N__59127));
    LocalMux I__13555 (
            .O(N__59130),
            .I(N__59123));
    LocalMux I__13554 (
            .O(N__59127),
            .I(N__59120));
    InMux I__13553 (
            .O(N__59126),
            .I(N__59117));
    Span4Mux_v I__13552 (
            .O(N__59123),
            .I(N__59112));
    Span4Mux_v I__13551 (
            .O(N__59120),
            .I(N__59107));
    LocalMux I__13550 (
            .O(N__59117),
            .I(N__59107));
    InMux I__13549 (
            .O(N__59116),
            .I(N__59104));
    InMux I__13548 (
            .O(N__59115),
            .I(N__59101));
    Span4Mux_h I__13547 (
            .O(N__59112),
            .I(N__59098));
    Span4Mux_v I__13546 (
            .O(N__59107),
            .I(N__59095));
    LocalMux I__13545 (
            .O(N__59104),
            .I(data_in_frame_18_7));
    LocalMux I__13544 (
            .O(N__59101),
            .I(data_in_frame_18_7));
    Odrv4 I__13543 (
            .O(N__59098),
            .I(data_in_frame_18_7));
    Odrv4 I__13542 (
            .O(N__59095),
            .I(data_in_frame_18_7));
    InMux I__13541 (
            .O(N__59086),
            .I(N__59082));
    InMux I__13540 (
            .O(N__59085),
            .I(N__59079));
    LocalMux I__13539 (
            .O(N__59082),
            .I(N__59076));
    LocalMux I__13538 (
            .O(N__59079),
            .I(N__59069));
    Span4Mux_v I__13537 (
            .O(N__59076),
            .I(N__59066));
    InMux I__13536 (
            .O(N__59075),
            .I(N__59061));
    InMux I__13535 (
            .O(N__59074),
            .I(N__59061));
    InMux I__13534 (
            .O(N__59073),
            .I(N__59056));
    InMux I__13533 (
            .O(N__59072),
            .I(N__59056));
    Odrv12 I__13532 (
            .O(N__59069),
            .I(\c0.n12052 ));
    Odrv4 I__13531 (
            .O(N__59066),
            .I(\c0.n12052 ));
    LocalMux I__13530 (
            .O(N__59061),
            .I(\c0.n12052 ));
    LocalMux I__13529 (
            .O(N__59056),
            .I(\c0.n12052 ));
    InMux I__13528 (
            .O(N__59047),
            .I(N__59043));
    InMux I__13527 (
            .O(N__59046),
            .I(N__59040));
    LocalMux I__13526 (
            .O(N__59043),
            .I(N__59036));
    LocalMux I__13525 (
            .O(N__59040),
            .I(N__59033));
    InMux I__13524 (
            .O(N__59039),
            .I(N__59029));
    Span4Mux_v I__13523 (
            .O(N__59036),
            .I(N__59024));
    Span4Mux_h I__13522 (
            .O(N__59033),
            .I(N__59024));
    InMux I__13521 (
            .O(N__59032),
            .I(N__59021));
    LocalMux I__13520 (
            .O(N__59029),
            .I(\c0.n19_adj_3056 ));
    Odrv4 I__13519 (
            .O(N__59024),
            .I(\c0.n19_adj_3056 ));
    LocalMux I__13518 (
            .O(N__59021),
            .I(\c0.n19_adj_3056 ));
    CascadeMux I__13517 (
            .O(N__59014),
            .I(\c0.n19_adj_3056_cascade_ ));
    InMux I__13516 (
            .O(N__59011),
            .I(N__59006));
    InMux I__13515 (
            .O(N__59010),
            .I(N__58999));
    InMux I__13514 (
            .O(N__59009),
            .I(N__58995));
    LocalMux I__13513 (
            .O(N__59006),
            .I(N__58992));
    InMux I__13512 (
            .O(N__59005),
            .I(N__58985));
    InMux I__13511 (
            .O(N__59004),
            .I(N__58985));
    InMux I__13510 (
            .O(N__59003),
            .I(N__58985));
    InMux I__13509 (
            .O(N__59002),
            .I(N__58982));
    LocalMux I__13508 (
            .O(N__58999),
            .I(N__58979));
    InMux I__13507 (
            .O(N__58998),
            .I(N__58976));
    LocalMux I__13506 (
            .O(N__58995),
            .I(N__58967));
    Sp12to4 I__13505 (
            .O(N__58992),
            .I(N__58967));
    LocalMux I__13504 (
            .O(N__58985),
            .I(N__58967));
    LocalMux I__13503 (
            .O(N__58982),
            .I(N__58967));
    Span4Mux_h I__13502 (
            .O(N__58979),
            .I(N__58962));
    LocalMux I__13501 (
            .O(N__58976),
            .I(N__58962));
    Span12Mux_v I__13500 (
            .O(N__58967),
            .I(N__58959));
    Odrv4 I__13499 (
            .O(N__58962),
            .I(\c0.n21045 ));
    Odrv12 I__13498 (
            .O(N__58959),
            .I(\c0.n21045 ));
    InMux I__13497 (
            .O(N__58954),
            .I(N__58951));
    LocalMux I__13496 (
            .O(N__58951),
            .I(N__58948));
    Span4Mux_h I__13495 (
            .O(N__58948),
            .I(N__58945));
    Odrv4 I__13494 (
            .O(N__58945),
            .I(\c0.n29_adj_3454 ));
    InMux I__13493 (
            .O(N__58942),
            .I(N__58937));
    InMux I__13492 (
            .O(N__58941),
            .I(N__58932));
    InMux I__13491 (
            .O(N__58940),
            .I(N__58932));
    LocalMux I__13490 (
            .O(N__58937),
            .I(N__58926));
    LocalMux I__13489 (
            .O(N__58932),
            .I(N__58926));
    InMux I__13488 (
            .O(N__58931),
            .I(N__58923));
    Span4Mux_v I__13487 (
            .O(N__58926),
            .I(N__58920));
    LocalMux I__13486 (
            .O(N__58923),
            .I(N__58917));
    Odrv4 I__13485 (
            .O(N__58920),
            .I(\c0.n18398 ));
    Odrv4 I__13484 (
            .O(N__58917),
            .I(\c0.n18398 ));
    InMux I__13483 (
            .O(N__58912),
            .I(N__58909));
    LocalMux I__13482 (
            .O(N__58909),
            .I(N__58906));
    Span4Mux_h I__13481 (
            .O(N__58906),
            .I(N__58903));
    Odrv4 I__13480 (
            .O(N__58903),
            .I(\c0.n6_adj_3239 ));
    InMux I__13479 (
            .O(N__58900),
            .I(N__58896));
    CascadeMux I__13478 (
            .O(N__58899),
            .I(N__58892));
    LocalMux I__13477 (
            .O(N__58896),
            .I(N__58889));
    InMux I__13476 (
            .O(N__58895),
            .I(N__58886));
    InMux I__13475 (
            .O(N__58892),
            .I(N__58883));
    Span4Mux_v I__13474 (
            .O(N__58889),
            .I(N__58878));
    LocalMux I__13473 (
            .O(N__58886),
            .I(N__58878));
    LocalMux I__13472 (
            .O(N__58883),
            .I(N__58875));
    Span4Mux_h I__13471 (
            .O(N__58878),
            .I(N__58872));
    Span4Mux_v I__13470 (
            .O(N__58875),
            .I(N__58868));
    Span4Mux_h I__13469 (
            .O(N__58872),
            .I(N__58865));
    InMux I__13468 (
            .O(N__58871),
            .I(N__58862));
    Span4Mux_h I__13467 (
            .O(N__58868),
            .I(N__58859));
    Span4Mux_v I__13466 (
            .O(N__58865),
            .I(N__58856));
    LocalMux I__13465 (
            .O(N__58862),
            .I(data_in_frame_22_2));
    Odrv4 I__13464 (
            .O(N__58859),
            .I(data_in_frame_22_2));
    Odrv4 I__13463 (
            .O(N__58856),
            .I(data_in_frame_22_2));
    CascadeMux I__13462 (
            .O(N__58849),
            .I(N__58846));
    InMux I__13461 (
            .O(N__58846),
            .I(N__58843));
    LocalMux I__13460 (
            .O(N__58843),
            .I(\c0.n19354 ));
    InMux I__13459 (
            .O(N__58840),
            .I(N__58836));
    InMux I__13458 (
            .O(N__58839),
            .I(N__58833));
    LocalMux I__13457 (
            .O(N__58836),
            .I(N__58829));
    LocalMux I__13456 (
            .O(N__58833),
            .I(N__58826));
    InMux I__13455 (
            .O(N__58832),
            .I(N__58823));
    Span4Mux_v I__13454 (
            .O(N__58829),
            .I(N__58819));
    Span4Mux_v I__13453 (
            .O(N__58826),
            .I(N__58814));
    LocalMux I__13452 (
            .O(N__58823),
            .I(N__58814));
    InMux I__13451 (
            .O(N__58822),
            .I(N__58811));
    Sp12to4 I__13450 (
            .O(N__58819),
            .I(N__58808));
    Span4Mux_h I__13449 (
            .O(N__58814),
            .I(N__58805));
    LocalMux I__13448 (
            .O(N__58811),
            .I(data_in_frame_22_7));
    Odrv12 I__13447 (
            .O(N__58808),
            .I(data_in_frame_22_7));
    Odrv4 I__13446 (
            .O(N__58805),
            .I(data_in_frame_22_7));
    InMux I__13445 (
            .O(N__58798),
            .I(N__58795));
    LocalMux I__13444 (
            .O(N__58795),
            .I(N__58791));
    InMux I__13443 (
            .O(N__58794),
            .I(N__58787));
    Span4Mux_h I__13442 (
            .O(N__58791),
            .I(N__58784));
    InMux I__13441 (
            .O(N__58790),
            .I(N__58781));
    LocalMux I__13440 (
            .O(N__58787),
            .I(N__58778));
    Span4Mux_v I__13439 (
            .O(N__58784),
            .I(N__58775));
    LocalMux I__13438 (
            .O(N__58781),
            .I(data_in_frame_22_3));
    Odrv4 I__13437 (
            .O(N__58778),
            .I(data_in_frame_22_3));
    Odrv4 I__13436 (
            .O(N__58775),
            .I(data_in_frame_22_3));
    InMux I__13435 (
            .O(N__58768),
            .I(N__58765));
    LocalMux I__13434 (
            .O(N__58765),
            .I(N__58762));
    Span4Mux_v I__13433 (
            .O(N__58762),
            .I(N__58757));
    InMux I__13432 (
            .O(N__58761),
            .I(N__58753));
    CascadeMux I__13431 (
            .O(N__58760),
            .I(N__58750));
    Sp12to4 I__13430 (
            .O(N__58757),
            .I(N__58747));
    InMux I__13429 (
            .O(N__58756),
            .I(N__58744));
    LocalMux I__13428 (
            .O(N__58753),
            .I(N__58741));
    InMux I__13427 (
            .O(N__58750),
            .I(N__58738));
    Span12Mux_h I__13426 (
            .O(N__58747),
            .I(N__58735));
    LocalMux I__13425 (
            .O(N__58744),
            .I(data_in_frame_24_0));
    Odrv4 I__13424 (
            .O(N__58741),
            .I(data_in_frame_24_0));
    LocalMux I__13423 (
            .O(N__58738),
            .I(data_in_frame_24_0));
    Odrv12 I__13422 (
            .O(N__58735),
            .I(data_in_frame_24_0));
    InMux I__13421 (
            .O(N__58726),
            .I(N__58719));
    InMux I__13420 (
            .O(N__58725),
            .I(N__58719));
    CascadeMux I__13419 (
            .O(N__58724),
            .I(N__58716));
    LocalMux I__13418 (
            .O(N__58719),
            .I(N__58712));
    InMux I__13417 (
            .O(N__58716),
            .I(N__58709));
    InMux I__13416 (
            .O(N__58715),
            .I(N__58705));
    Span4Mux_h I__13415 (
            .O(N__58712),
            .I(N__58700));
    LocalMux I__13414 (
            .O(N__58709),
            .I(N__58700));
    CascadeMux I__13413 (
            .O(N__58708),
            .I(N__58697));
    LocalMux I__13412 (
            .O(N__58705),
            .I(N__58694));
    Span4Mux_v I__13411 (
            .O(N__58700),
            .I(N__58691));
    InMux I__13410 (
            .O(N__58697),
            .I(N__58688));
    Span12Mux_v I__13409 (
            .O(N__58694),
            .I(N__58685));
    Sp12to4 I__13408 (
            .O(N__58691),
            .I(N__58682));
    LocalMux I__13407 (
            .O(N__58688),
            .I(\c0.data_in_frame_26_2 ));
    Odrv12 I__13406 (
            .O(N__58685),
            .I(\c0.data_in_frame_26_2 ));
    Odrv12 I__13405 (
            .O(N__58682),
            .I(\c0.data_in_frame_26_2 ));
    InMux I__13404 (
            .O(N__58675),
            .I(N__58672));
    LocalMux I__13403 (
            .O(N__58672),
            .I(\c0.n93_adj_3385 ));
    InMux I__13402 (
            .O(N__58669),
            .I(N__58664));
    InMux I__13401 (
            .O(N__58668),
            .I(N__58661));
    InMux I__13400 (
            .O(N__58667),
            .I(N__58658));
    LocalMux I__13399 (
            .O(N__58664),
            .I(N__58655));
    LocalMux I__13398 (
            .O(N__58661),
            .I(N__58650));
    LocalMux I__13397 (
            .O(N__58658),
            .I(N__58650));
    Span4Mux_h I__13396 (
            .O(N__58655),
            .I(N__58646));
    Span4Mux_h I__13395 (
            .O(N__58650),
            .I(N__58643));
    InMux I__13394 (
            .O(N__58649),
            .I(N__58640));
    Odrv4 I__13393 (
            .O(N__58646),
            .I(\c0.n32_adj_3057 ));
    Odrv4 I__13392 (
            .O(N__58643),
            .I(\c0.n32_adj_3057 ));
    LocalMux I__13391 (
            .O(N__58640),
            .I(\c0.n32_adj_3057 ));
    InMux I__13390 (
            .O(N__58633),
            .I(N__58630));
    LocalMux I__13389 (
            .O(N__58630),
            .I(N__58626));
    InMux I__13388 (
            .O(N__58629),
            .I(N__58623));
    Span4Mux_h I__13387 (
            .O(N__58626),
            .I(N__58620));
    LocalMux I__13386 (
            .O(N__58623),
            .I(N__58617));
    Odrv4 I__13385 (
            .O(N__58620),
            .I(\c0.n62 ));
    Odrv4 I__13384 (
            .O(N__58617),
            .I(\c0.n62 ));
    InMux I__13383 (
            .O(N__58612),
            .I(N__58609));
    LocalMux I__13382 (
            .O(N__58609),
            .I(\c0.n68 ));
    InMux I__13381 (
            .O(N__58606),
            .I(N__58603));
    LocalMux I__13380 (
            .O(N__58603),
            .I(N__58600));
    Span4Mux_v I__13379 (
            .O(N__58600),
            .I(N__58595));
    InMux I__13378 (
            .O(N__58599),
            .I(N__58592));
    InMux I__13377 (
            .O(N__58598),
            .I(N__58589));
    Odrv4 I__13376 (
            .O(N__58595),
            .I(\c0.n19502 ));
    LocalMux I__13375 (
            .O(N__58592),
            .I(\c0.n19502 ));
    LocalMux I__13374 (
            .O(N__58589),
            .I(\c0.n19502 ));
    InMux I__13373 (
            .O(N__58582),
            .I(N__58579));
    LocalMux I__13372 (
            .O(N__58579),
            .I(N__58576));
    Odrv12 I__13371 (
            .O(N__58576),
            .I(\c0.n20_adj_3536 ));
    CascadeMux I__13370 (
            .O(N__58573),
            .I(N__58570));
    InMux I__13369 (
            .O(N__58570),
            .I(N__58567));
    LocalMux I__13368 (
            .O(N__58567),
            .I(N__58564));
    Span4Mux_v I__13367 (
            .O(N__58564),
            .I(N__58561));
    Span4Mux_h I__13366 (
            .O(N__58561),
            .I(N__58558));
    Span4Mux_v I__13365 (
            .O(N__58558),
            .I(N__58555));
    Odrv4 I__13364 (
            .O(N__58555),
            .I(\c0.n23_adj_3534 ));
    CascadeMux I__13363 (
            .O(N__58552),
            .I(N__58547));
    InMux I__13362 (
            .O(N__58551),
            .I(N__58544));
    CascadeMux I__13361 (
            .O(N__58550),
            .I(N__58541));
    InMux I__13360 (
            .O(N__58547),
            .I(N__58538));
    LocalMux I__13359 (
            .O(N__58544),
            .I(N__58535));
    InMux I__13358 (
            .O(N__58541),
            .I(N__58532));
    LocalMux I__13357 (
            .O(N__58538),
            .I(N__58529));
    Span4Mux_h I__13356 (
            .O(N__58535),
            .I(N__58526));
    LocalMux I__13355 (
            .O(N__58532),
            .I(N__58523));
    Span4Mux_v I__13354 (
            .O(N__58529),
            .I(N__58518));
    Span4Mux_h I__13353 (
            .O(N__58526),
            .I(N__58518));
    Span4Mux_h I__13352 (
            .O(N__58523),
            .I(N__58515));
    Odrv4 I__13351 (
            .O(N__58518),
            .I(\c0.n40_adj_3374 ));
    Odrv4 I__13350 (
            .O(N__58515),
            .I(\c0.n40_adj_3374 ));
    CascadeMux I__13349 (
            .O(N__58510),
            .I(\c0.n38_adj_3062_cascade_ ));
    InMux I__13348 (
            .O(N__58507),
            .I(N__58503));
    InMux I__13347 (
            .O(N__58506),
            .I(N__58500));
    LocalMux I__13346 (
            .O(N__58503),
            .I(\c0.n39_adj_3384 ));
    LocalMux I__13345 (
            .O(N__58500),
            .I(\c0.n39_adj_3384 ));
    InMux I__13344 (
            .O(N__58495),
            .I(N__58492));
    LocalMux I__13343 (
            .O(N__58492),
            .I(N__58488));
    InMux I__13342 (
            .O(N__58491),
            .I(N__58485));
    Span4Mux_h I__13341 (
            .O(N__58488),
            .I(N__58482));
    LocalMux I__13340 (
            .O(N__58485),
            .I(N__58479));
    Span4Mux_h I__13339 (
            .O(N__58482),
            .I(N__58476));
    Span4Mux_h I__13338 (
            .O(N__58479),
            .I(N__58473));
    Odrv4 I__13337 (
            .O(N__58476),
            .I(\c0.n93_adj_3329 ));
    Odrv4 I__13336 (
            .O(N__58473),
            .I(\c0.n93_adj_3329 ));
    InMux I__13335 (
            .O(N__58468),
            .I(N__58463));
    CascadeMux I__13334 (
            .O(N__58467),
            .I(N__58458));
    InMux I__13333 (
            .O(N__58466),
            .I(N__58455));
    LocalMux I__13332 (
            .O(N__58463),
            .I(N__58452));
    InMux I__13331 (
            .O(N__58462),
            .I(N__58449));
    InMux I__13330 (
            .O(N__58461),
            .I(N__58446));
    InMux I__13329 (
            .O(N__58458),
            .I(N__58443));
    LocalMux I__13328 (
            .O(N__58455),
            .I(N__58440));
    Span4Mux_v I__13327 (
            .O(N__58452),
            .I(N__58433));
    LocalMux I__13326 (
            .O(N__58449),
            .I(N__58433));
    LocalMux I__13325 (
            .O(N__58446),
            .I(N__58433));
    LocalMux I__13324 (
            .O(N__58443),
            .I(N__58428));
    Span4Mux_v I__13323 (
            .O(N__58440),
            .I(N__58423));
    Span4Mux_v I__13322 (
            .O(N__58433),
            .I(N__58423));
    InMux I__13321 (
            .O(N__58432),
            .I(N__58420));
    InMux I__13320 (
            .O(N__58431),
            .I(N__58417));
    Odrv12 I__13319 (
            .O(N__58428),
            .I(\c0.data_in_frame_8_3 ));
    Odrv4 I__13318 (
            .O(N__58423),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__13317 (
            .O(N__58420),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__13316 (
            .O(N__58417),
            .I(\c0.data_in_frame_8_3 ));
    CascadeMux I__13315 (
            .O(N__58408),
            .I(N__58405));
    InMux I__13314 (
            .O(N__58405),
            .I(N__58401));
    InMux I__13313 (
            .O(N__58404),
            .I(N__58398));
    LocalMux I__13312 (
            .O(N__58401),
            .I(N__58395));
    LocalMux I__13311 (
            .O(N__58398),
            .I(N__58392));
    Span4Mux_v I__13310 (
            .O(N__58395),
            .I(N__58387));
    Span4Mux_v I__13309 (
            .O(N__58392),
            .I(N__58387));
    Span4Mux_h I__13308 (
            .O(N__58387),
            .I(N__58384));
    Odrv4 I__13307 (
            .O(N__58384),
            .I(\c0.n19505 ));
    InMux I__13306 (
            .O(N__58381),
            .I(N__58378));
    LocalMux I__13305 (
            .O(N__58378),
            .I(\c0.n26_adj_3537 ));
    CascadeMux I__13304 (
            .O(N__58375),
            .I(\c0.n20917_cascade_ ));
    InMux I__13303 (
            .O(N__58372),
            .I(N__58369));
    LocalMux I__13302 (
            .O(N__58369),
            .I(N__58365));
    InMux I__13301 (
            .O(N__58368),
            .I(N__58362));
    Span4Mux_v I__13300 (
            .O(N__58365),
            .I(N__58359));
    LocalMux I__13299 (
            .O(N__58362),
            .I(N__58354));
    Span4Mux_h I__13298 (
            .O(N__58359),
            .I(N__58354));
    Span4Mux_v I__13297 (
            .O(N__58354),
            .I(N__58350));
    InMux I__13296 (
            .O(N__58353),
            .I(N__58347));
    Odrv4 I__13295 (
            .O(N__58350),
            .I(\c0.n19524 ));
    LocalMux I__13294 (
            .O(N__58347),
            .I(\c0.n19524 ));
    CascadeMux I__13293 (
            .O(N__58342),
            .I(\c0.n6_adj_3433_cascade_ ));
    CascadeMux I__13292 (
            .O(N__58339),
            .I(\c0.n18375_cascade_ ));
    InMux I__13291 (
            .O(N__58336),
            .I(N__58330));
    InMux I__13290 (
            .O(N__58335),
            .I(N__58330));
    LocalMux I__13289 (
            .O(N__58330),
            .I(\c0.n58 ));
    CascadeMux I__13288 (
            .O(N__58327),
            .I(N__58324));
    InMux I__13287 (
            .O(N__58324),
            .I(N__58321));
    LocalMux I__13286 (
            .O(N__58321),
            .I(N__58318));
    Span4Mux_h I__13285 (
            .O(N__58318),
            .I(N__58315));
    Span4Mux_h I__13284 (
            .O(N__58315),
            .I(N__58312));
    Span4Mux_v I__13283 (
            .O(N__58312),
            .I(N__58309));
    Odrv4 I__13282 (
            .O(N__58309),
            .I(\c0.n16_adj_3489 ));
    InMux I__13281 (
            .O(N__58306),
            .I(N__58300));
    InMux I__13280 (
            .O(N__58305),
            .I(N__58300));
    LocalMux I__13279 (
            .O(N__58300),
            .I(N__58297));
    Span4Mux_h I__13278 (
            .O(N__58297),
            .I(N__58294));
    Odrv4 I__13277 (
            .O(N__58294),
            .I(\c0.n31_adj_3126 ));
    CascadeMux I__13276 (
            .O(N__58291),
            .I(\c0.n10_adj_3425_cascade_ ));
    InMux I__13275 (
            .O(N__58288),
            .I(N__58284));
    InMux I__13274 (
            .O(N__58287),
            .I(N__58281));
    LocalMux I__13273 (
            .O(N__58284),
            .I(\c0.n42_adj_3130 ));
    LocalMux I__13272 (
            .O(N__58281),
            .I(\c0.n42_adj_3130 ));
    InMux I__13271 (
            .O(N__58276),
            .I(N__58273));
    LocalMux I__13270 (
            .O(N__58273),
            .I(N__58270));
    Span4Mux_h I__13269 (
            .O(N__58270),
            .I(N__58267));
    Odrv4 I__13268 (
            .O(N__58267),
            .I(\c0.n92_adj_3272 ));
    InMux I__13267 (
            .O(N__58264),
            .I(N__58261));
    LocalMux I__13266 (
            .O(N__58261),
            .I(\c0.n39_adj_3269 ));
    InMux I__13265 (
            .O(N__58258),
            .I(N__58255));
    LocalMux I__13264 (
            .O(N__58255),
            .I(N__58252));
    Span4Mux_h I__13263 (
            .O(N__58252),
            .I(N__58249));
    Span4Mux_v I__13262 (
            .O(N__58249),
            .I(N__58244));
    InMux I__13261 (
            .O(N__58248),
            .I(N__58239));
    InMux I__13260 (
            .O(N__58247),
            .I(N__58239));
    Span4Mux_h I__13259 (
            .O(N__58244),
            .I(N__58236));
    LocalMux I__13258 (
            .O(N__58239),
            .I(N__58233));
    Odrv4 I__13257 (
            .O(N__58236),
            .I(\c0.n36_adj_3275 ));
    Odrv12 I__13256 (
            .O(N__58233),
            .I(\c0.n36_adj_3275 ));
    CascadeMux I__13255 (
            .O(N__58228),
            .I(N__58224));
    InMux I__13254 (
            .O(N__58227),
            .I(N__58221));
    InMux I__13253 (
            .O(N__58224),
            .I(N__58218));
    LocalMux I__13252 (
            .O(N__58221),
            .I(N__58212));
    LocalMux I__13251 (
            .O(N__58218),
            .I(N__58212));
    InMux I__13250 (
            .O(N__58217),
            .I(N__58209));
    Odrv4 I__13249 (
            .O(N__58212),
            .I(\c0.n38_adj_3270 ));
    LocalMux I__13248 (
            .O(N__58209),
            .I(\c0.n38_adj_3270 ));
    CascadeMux I__13247 (
            .O(N__58204),
            .I(\c0.n39_adj_3269_cascade_ ));
    InMux I__13246 (
            .O(N__58201),
            .I(N__58194));
    InMux I__13245 (
            .O(N__58200),
            .I(N__58194));
    InMux I__13244 (
            .O(N__58199),
            .I(N__58191));
    LocalMux I__13243 (
            .O(N__58194),
            .I(\c0.n37_adj_3268 ));
    LocalMux I__13242 (
            .O(N__58191),
            .I(\c0.n37_adj_3268 ));
    InMux I__13241 (
            .O(N__58186),
            .I(N__58183));
    LocalMux I__13240 (
            .O(N__58183),
            .I(N__58180));
    Span4Mux_v I__13239 (
            .O(N__58180),
            .I(N__58177));
    Span4Mux_h I__13238 (
            .O(N__58177),
            .I(N__58174));
    Odrv4 I__13237 (
            .O(N__58174),
            .I(\c0.n94_adj_3375 ));
    CascadeMux I__13236 (
            .O(N__58171),
            .I(\c0.n92_adj_3377_cascade_ ));
    InMux I__13235 (
            .O(N__58168),
            .I(N__58165));
    LocalMux I__13234 (
            .O(N__58165),
            .I(N__58162));
    Odrv4 I__13233 (
            .O(N__58162),
            .I(\c0.n91_adj_3389 ));
    InMux I__13232 (
            .O(N__58159),
            .I(N__58156));
    LocalMux I__13231 (
            .O(N__58156),
            .I(N__58153));
    Odrv12 I__13230 (
            .O(N__58153),
            .I(\c0.n100_adj_3420 ));
    CascadeMux I__13229 (
            .O(N__58150),
            .I(N__58147));
    InMux I__13228 (
            .O(N__58147),
            .I(N__58144));
    LocalMux I__13227 (
            .O(N__58144),
            .I(N__58141));
    Span4Mux_h I__13226 (
            .O(N__58141),
            .I(N__58138));
    Span4Mux_v I__13225 (
            .O(N__58138),
            .I(N__58135));
    Span4Mux_h I__13224 (
            .O(N__58135),
            .I(N__58132));
    Span4Mux_h I__13223 (
            .O(N__58132),
            .I(N__58127));
    InMux I__13222 (
            .O(N__58131),
            .I(N__58124));
    InMux I__13221 (
            .O(N__58130),
            .I(N__58121));
    Odrv4 I__13220 (
            .O(N__58127),
            .I(\c0.n11942 ));
    LocalMux I__13219 (
            .O(N__58124),
            .I(\c0.n11942 ));
    LocalMux I__13218 (
            .O(N__58121),
            .I(\c0.n11942 ));
    CascadeMux I__13217 (
            .O(N__58114),
            .I(N__58111));
    InMux I__13216 (
            .O(N__58111),
            .I(N__58108));
    LocalMux I__13215 (
            .O(N__58108),
            .I(N__58105));
    Span4Mux_h I__13214 (
            .O(N__58105),
            .I(N__58102));
    Odrv4 I__13213 (
            .O(N__58102),
            .I(\c0.n12_adj_3208 ));
    InMux I__13212 (
            .O(N__58099),
            .I(N__58094));
    InMux I__13211 (
            .O(N__58098),
            .I(N__58089));
    InMux I__13210 (
            .O(N__58097),
            .I(N__58089));
    LocalMux I__13209 (
            .O(N__58094),
            .I(\c0.n10_adj_3425 ));
    LocalMux I__13208 (
            .O(N__58089),
            .I(\c0.n10_adj_3425 ));
    InMux I__13207 (
            .O(N__58084),
            .I(N__58081));
    LocalMux I__13206 (
            .O(N__58081),
            .I(N__58078));
    Span4Mux_v I__13205 (
            .O(N__58078),
            .I(N__58075));
    Odrv4 I__13204 (
            .O(N__58075),
            .I(\c0.n82 ));
    InMux I__13203 (
            .O(N__58072),
            .I(N__58069));
    LocalMux I__13202 (
            .O(N__58069),
            .I(N__58064));
    InMux I__13201 (
            .O(N__58068),
            .I(N__58059));
    InMux I__13200 (
            .O(N__58067),
            .I(N__58059));
    Span4Mux_v I__13199 (
            .O(N__58064),
            .I(N__58054));
    LocalMux I__13198 (
            .O(N__58059),
            .I(N__58054));
    Span4Mux_h I__13197 (
            .O(N__58054),
            .I(N__58050));
    InMux I__13196 (
            .O(N__58053),
            .I(N__58047));
    Odrv4 I__13195 (
            .O(N__58050),
            .I(\c0.n20085 ));
    LocalMux I__13194 (
            .O(N__58047),
            .I(\c0.n20085 ));
    InMux I__13193 (
            .O(N__58042),
            .I(N__58038));
    InMux I__13192 (
            .O(N__58041),
            .I(N__58034));
    LocalMux I__13191 (
            .O(N__58038),
            .I(N__58031));
    InMux I__13190 (
            .O(N__58037),
            .I(N__58028));
    LocalMux I__13189 (
            .O(N__58034),
            .I(N__58025));
    Span4Mux_h I__13188 (
            .O(N__58031),
            .I(N__58017));
    LocalMux I__13187 (
            .O(N__58028),
            .I(N__58017));
    Span4Mux_v I__13186 (
            .O(N__58025),
            .I(N__58017));
    InMux I__13185 (
            .O(N__58024),
            .I(N__58014));
    Odrv4 I__13184 (
            .O(N__58017),
            .I(\c0.n19244 ));
    LocalMux I__13183 (
            .O(N__58014),
            .I(\c0.n19244 ));
    InMux I__13182 (
            .O(N__58009),
            .I(N__58006));
    LocalMux I__13181 (
            .O(N__58006),
            .I(N__58003));
    Span4Mux_h I__13180 (
            .O(N__58003),
            .I(N__58000));
    Span4Mux_h I__13179 (
            .O(N__58000),
            .I(N__57997));
    Odrv4 I__13178 (
            .O(N__57997),
            .I(\c0.n88_adj_3422 ));
    InMux I__13177 (
            .O(N__57994),
            .I(N__57991));
    LocalMux I__13176 (
            .O(N__57991),
            .I(\c0.n25_adj_3510 ));
    InMux I__13175 (
            .O(N__57988),
            .I(N__57982));
    InMux I__13174 (
            .O(N__57987),
            .I(N__57982));
    LocalMux I__13173 (
            .O(N__57982),
            .I(N__57979));
    Span4Mux_h I__13172 (
            .O(N__57979),
            .I(N__57976));
    Odrv4 I__13171 (
            .O(N__57976),
            .I(\c0.n56 ));
    InMux I__13170 (
            .O(N__57973),
            .I(N__57970));
    LocalMux I__13169 (
            .O(N__57970),
            .I(N__57966));
    InMux I__13168 (
            .O(N__57969),
            .I(N__57963));
    Span4Mux_v I__13167 (
            .O(N__57966),
            .I(N__57960));
    LocalMux I__13166 (
            .O(N__57963),
            .I(N__57957));
    Odrv4 I__13165 (
            .O(N__57960),
            .I(\c0.n44_adj_3125 ));
    Odrv4 I__13164 (
            .O(N__57957),
            .I(\c0.n44_adj_3125 ));
    InMux I__13163 (
            .O(N__57952),
            .I(N__57948));
    InMux I__13162 (
            .O(N__57951),
            .I(N__57945));
    LocalMux I__13161 (
            .O(N__57948),
            .I(\c0.n11_adj_3124 ));
    LocalMux I__13160 (
            .O(N__57945),
            .I(\c0.n11_adj_3124 ));
    CascadeMux I__13159 (
            .O(N__57940),
            .I(N__57937));
    InMux I__13158 (
            .O(N__57937),
            .I(N__57934));
    LocalMux I__13157 (
            .O(N__57934),
            .I(\c0.n48_adj_3313 ));
    CascadeMux I__13156 (
            .O(N__57931),
            .I(\c0.n35_cascade_ ));
    InMux I__13155 (
            .O(N__57928),
            .I(N__57925));
    LocalMux I__13154 (
            .O(N__57925),
            .I(\c0.n67_adj_3092 ));
    InMux I__13153 (
            .O(N__57922),
            .I(N__57916));
    InMux I__13152 (
            .O(N__57921),
            .I(N__57916));
    LocalMux I__13151 (
            .O(N__57916),
            .I(N__57913));
    Odrv4 I__13150 (
            .O(N__57913),
            .I(\c0.n43_adj_3089 ));
    CascadeMux I__13149 (
            .O(N__57910),
            .I(N__57906));
    CascadeMux I__13148 (
            .O(N__57909),
            .I(N__57903));
    InMux I__13147 (
            .O(N__57906),
            .I(N__57900));
    InMux I__13146 (
            .O(N__57903),
            .I(N__57897));
    LocalMux I__13145 (
            .O(N__57900),
            .I(N__57894));
    LocalMux I__13144 (
            .O(N__57897),
            .I(N__57889));
    Span4Mux_h I__13143 (
            .O(N__57894),
            .I(N__57889));
    Span4Mux_v I__13142 (
            .O(N__57889),
            .I(N__57886));
    Odrv4 I__13141 (
            .O(N__57886),
            .I(\c0.n41_adj_3085 ));
    InMux I__13140 (
            .O(N__57883),
            .I(N__57879));
    InMux I__13139 (
            .O(N__57882),
            .I(N__57876));
    LocalMux I__13138 (
            .O(N__57879),
            .I(\c0.n42_adj_3086 ));
    LocalMux I__13137 (
            .O(N__57876),
            .I(\c0.n42_adj_3086 ));
    InMux I__13136 (
            .O(N__57871),
            .I(N__57868));
    LocalMux I__13135 (
            .O(N__57868),
            .I(\c0.n60_adj_3127 ));
    CascadeMux I__13134 (
            .O(N__57865),
            .I(\c0.n55_adj_3128_cascade_ ));
    InMux I__13133 (
            .O(N__57862),
            .I(N__57859));
    LocalMux I__13132 (
            .O(N__57859),
            .I(N__57854));
    InMux I__13131 (
            .O(N__57858),
            .I(N__57849));
    InMux I__13130 (
            .O(N__57857),
            .I(N__57849));
    Span4Mux_h I__13129 (
            .O(N__57854),
            .I(N__57846));
    LocalMux I__13128 (
            .O(N__57849),
            .I(N__57841));
    Span4Mux_h I__13127 (
            .O(N__57846),
            .I(N__57841));
    Odrv4 I__13126 (
            .O(N__57841),
            .I(\c0.n19749 ));
    InMux I__13125 (
            .O(N__57838),
            .I(N__57834));
    InMux I__13124 (
            .O(N__57837),
            .I(N__57831));
    LocalMux I__13123 (
            .O(N__57834),
            .I(N__57828));
    LocalMux I__13122 (
            .O(N__57831),
            .I(N__57825));
    Odrv4 I__13121 (
            .O(N__57828),
            .I(\c0.n69 ));
    Odrv4 I__13120 (
            .O(N__57825),
            .I(\c0.n69 ));
    CascadeMux I__13119 (
            .O(N__57820),
            .I(N__57816));
    InMux I__13118 (
            .O(N__57819),
            .I(N__57813));
    InMux I__13117 (
            .O(N__57816),
            .I(N__57810));
    LocalMux I__13116 (
            .O(N__57813),
            .I(N__57807));
    LocalMux I__13115 (
            .O(N__57810),
            .I(\c0.n28_adj_3059 ));
    Odrv4 I__13114 (
            .O(N__57807),
            .I(\c0.n28_adj_3059 ));
    CascadeMux I__13113 (
            .O(N__57802),
            .I(\c0.n38_adj_3058_cascade_ ));
    InMux I__13112 (
            .O(N__57799),
            .I(N__57796));
    LocalMux I__13111 (
            .O(N__57796),
            .I(\c0.n32_adj_3060 ));
    CascadeMux I__13110 (
            .O(N__57793),
            .I(\c0.n8_adj_3061_cascade_ ));
    InMux I__13109 (
            .O(N__57790),
            .I(N__57786));
    InMux I__13108 (
            .O(N__57789),
            .I(N__57783));
    LocalMux I__13107 (
            .O(N__57786),
            .I(N__57778));
    LocalMux I__13106 (
            .O(N__57783),
            .I(N__57778));
    Span4Mux_v I__13105 (
            .O(N__57778),
            .I(N__57775));
    Span4Mux_h I__13104 (
            .O(N__57775),
            .I(N__57772));
    Odrv4 I__13103 (
            .O(N__57772),
            .I(\c0.n52 ));
    InMux I__13102 (
            .O(N__57769),
            .I(N__57766));
    LocalMux I__13101 (
            .O(N__57766),
            .I(\c0.n8_adj_3061 ));
    CascadeMux I__13100 (
            .O(N__57763),
            .I(\c0.n43_adj_3285_cascade_ ));
    InMux I__13099 (
            .O(N__57760),
            .I(N__57757));
    LocalMux I__13098 (
            .O(N__57757),
            .I(\c0.n53 ));
    InMux I__13097 (
            .O(N__57754),
            .I(N__57751));
    LocalMux I__13096 (
            .O(N__57751),
            .I(N__57748));
    Span4Mux_h I__13095 (
            .O(N__57748),
            .I(N__57744));
    InMux I__13094 (
            .O(N__57747),
            .I(N__57741));
    Odrv4 I__13093 (
            .O(N__57744),
            .I(\c0.n4_adj_3123 ));
    LocalMux I__13092 (
            .O(N__57741),
            .I(\c0.n4_adj_3123 ));
    InMux I__13091 (
            .O(N__57736),
            .I(N__57733));
    LocalMux I__13090 (
            .O(N__57733),
            .I(N__57729));
    CascadeMux I__13089 (
            .O(N__57732),
            .I(N__57726));
    Span4Mux_v I__13088 (
            .O(N__57729),
            .I(N__57720));
    InMux I__13087 (
            .O(N__57726),
            .I(N__57717));
    InMux I__13086 (
            .O(N__57725),
            .I(N__57714));
    CascadeMux I__13085 (
            .O(N__57724),
            .I(N__57710));
    InMux I__13084 (
            .O(N__57723),
            .I(N__57706));
    Span4Mux_h I__13083 (
            .O(N__57720),
            .I(N__57701));
    LocalMux I__13082 (
            .O(N__57717),
            .I(N__57701));
    LocalMux I__13081 (
            .O(N__57714),
            .I(N__57698));
    InMux I__13080 (
            .O(N__57713),
            .I(N__57693));
    InMux I__13079 (
            .O(N__57710),
            .I(N__57693));
    InMux I__13078 (
            .O(N__57709),
            .I(N__57689));
    LocalMux I__13077 (
            .O(N__57706),
            .I(N__57682));
    Span4Mux_h I__13076 (
            .O(N__57701),
            .I(N__57682));
    Span4Mux_h I__13075 (
            .O(N__57698),
            .I(N__57682));
    LocalMux I__13074 (
            .O(N__57693),
            .I(N__57679));
    InMux I__13073 (
            .O(N__57692),
            .I(N__57676));
    LocalMux I__13072 (
            .O(N__57689),
            .I(N__57673));
    Span4Mux_v I__13071 (
            .O(N__57682),
            .I(N__57670));
    Span4Mux_v I__13070 (
            .O(N__57679),
            .I(N__57667));
    LocalMux I__13069 (
            .O(N__57676),
            .I(data_in_frame_16_7));
    Odrv12 I__13068 (
            .O(N__57673),
            .I(data_in_frame_16_7));
    Odrv4 I__13067 (
            .O(N__57670),
            .I(data_in_frame_16_7));
    Odrv4 I__13066 (
            .O(N__57667),
            .I(data_in_frame_16_7));
    InMux I__13065 (
            .O(N__57658),
            .I(N__57652));
    InMux I__13064 (
            .O(N__57657),
            .I(N__57647));
    InMux I__13063 (
            .O(N__57656),
            .I(N__57647));
    InMux I__13062 (
            .O(N__57655),
            .I(N__57642));
    LocalMux I__13061 (
            .O(N__57652),
            .I(N__57637));
    LocalMux I__13060 (
            .O(N__57647),
            .I(N__57637));
    InMux I__13059 (
            .O(N__57646),
            .I(N__57634));
    InMux I__13058 (
            .O(N__57645),
            .I(N__57629));
    LocalMux I__13057 (
            .O(N__57642),
            .I(N__57626));
    Span4Mux_v I__13056 (
            .O(N__57637),
            .I(N__57623));
    LocalMux I__13055 (
            .O(N__57634),
            .I(N__57620));
    CascadeMux I__13054 (
            .O(N__57633),
            .I(N__57617));
    InMux I__13053 (
            .O(N__57632),
            .I(N__57614));
    LocalMux I__13052 (
            .O(N__57629),
            .I(N__57611));
    Span4Mux_v I__13051 (
            .O(N__57626),
            .I(N__57606));
    Span4Mux_v I__13050 (
            .O(N__57623),
            .I(N__57606));
    Span4Mux_h I__13049 (
            .O(N__57620),
            .I(N__57603));
    InMux I__13048 (
            .O(N__57617),
            .I(N__57600));
    LocalMux I__13047 (
            .O(N__57614),
            .I(\c0.data_in_frame_12_5 ));
    Odrv12 I__13046 (
            .O(N__57611),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__13045 (
            .O(N__57606),
            .I(\c0.data_in_frame_12_5 ));
    Odrv4 I__13044 (
            .O(N__57603),
            .I(\c0.data_in_frame_12_5 ));
    LocalMux I__13043 (
            .O(N__57600),
            .I(\c0.data_in_frame_12_5 ));
    CascadeMux I__13042 (
            .O(N__57589),
            .I(\c0.n12_adj_3554_cascade_ ));
    InMux I__13041 (
            .O(N__57586),
            .I(N__57583));
    LocalMux I__13040 (
            .O(N__57583),
            .I(N__57578));
    InMux I__13039 (
            .O(N__57582),
            .I(N__57573));
    InMux I__13038 (
            .O(N__57581),
            .I(N__57573));
    Span4Mux_v I__13037 (
            .O(N__57578),
            .I(N__57568));
    LocalMux I__13036 (
            .O(N__57573),
            .I(N__57565));
    InMux I__13035 (
            .O(N__57572),
            .I(N__57562));
    InMux I__13034 (
            .O(N__57571),
            .I(N__57559));
    Span4Mux_h I__13033 (
            .O(N__57568),
            .I(N__57552));
    Span4Mux_v I__13032 (
            .O(N__57565),
            .I(N__57552));
    LocalMux I__13031 (
            .O(N__57562),
            .I(N__57552));
    LocalMux I__13030 (
            .O(N__57559),
            .I(\c0.n20151 ));
    Odrv4 I__13029 (
            .O(N__57552),
            .I(\c0.n20151 ));
    InMux I__13028 (
            .O(N__57547),
            .I(N__57544));
    LocalMux I__13027 (
            .O(N__57544),
            .I(N__57541));
    Span4Mux_h I__13026 (
            .O(N__57541),
            .I(N__57538));
    Odrv4 I__13025 (
            .O(N__57538),
            .I(\c0.n20542 ));
    CascadeMux I__13024 (
            .O(N__57535),
            .I(\c0.n20542_cascade_ ));
    InMux I__13023 (
            .O(N__57532),
            .I(N__57529));
    LocalMux I__13022 (
            .O(N__57529),
            .I(N__57526));
    Span4Mux_h I__13021 (
            .O(N__57526),
            .I(N__57522));
    InMux I__13020 (
            .O(N__57525),
            .I(N__57519));
    Odrv4 I__13019 (
            .O(N__57522),
            .I(\c0.n45_adj_3423 ));
    LocalMux I__13018 (
            .O(N__57519),
            .I(\c0.n45_adj_3423 ));
    CascadeMux I__13017 (
            .O(N__57514),
            .I(\c0.n25_adj_3510_cascade_ ));
    InMux I__13016 (
            .O(N__57511),
            .I(N__57508));
    LocalMux I__13015 (
            .O(N__57508),
            .I(N__57505));
    Odrv4 I__13014 (
            .O(N__57505),
            .I(\c0.n58_adj_3511 ));
    InMux I__13013 (
            .O(N__57502),
            .I(N__57496));
    InMux I__13012 (
            .O(N__57501),
            .I(N__57493));
    CascadeMux I__13011 (
            .O(N__57500),
            .I(N__57490));
    CascadeMux I__13010 (
            .O(N__57499),
            .I(N__57487));
    LocalMux I__13009 (
            .O(N__57496),
            .I(N__57484));
    LocalMux I__13008 (
            .O(N__57493),
            .I(N__57481));
    InMux I__13007 (
            .O(N__57490),
            .I(N__57478));
    InMux I__13006 (
            .O(N__57487),
            .I(N__57475));
    Span4Mux_h I__13005 (
            .O(N__57484),
            .I(N__57472));
    Span4Mux_v I__13004 (
            .O(N__57481),
            .I(N__57467));
    LocalMux I__13003 (
            .O(N__57478),
            .I(N__57467));
    LocalMux I__13002 (
            .O(N__57475),
            .I(\c0.data_in_frame_14_1 ));
    Odrv4 I__13001 (
            .O(N__57472),
            .I(\c0.data_in_frame_14_1 ));
    Odrv4 I__13000 (
            .O(N__57467),
            .I(\c0.data_in_frame_14_1 ));
    CascadeMux I__12999 (
            .O(N__57460),
            .I(N__57457));
    InMux I__12998 (
            .O(N__57457),
            .I(N__57447));
    InMux I__12997 (
            .O(N__57456),
            .I(N__57447));
    InMux I__12996 (
            .O(N__57455),
            .I(N__57447));
    InMux I__12995 (
            .O(N__57454),
            .I(N__57444));
    LocalMux I__12994 (
            .O(N__57447),
            .I(N__57438));
    LocalMux I__12993 (
            .O(N__57444),
            .I(N__57438));
    InMux I__12992 (
            .O(N__57443),
            .I(N__57435));
    Span4Mux_v I__12991 (
            .O(N__57438),
            .I(N__57429));
    LocalMux I__12990 (
            .O(N__57435),
            .I(N__57429));
    CascadeMux I__12989 (
            .O(N__57434),
            .I(N__57426));
    Span4Mux_h I__12988 (
            .O(N__57429),
            .I(N__57423));
    InMux I__12987 (
            .O(N__57426),
            .I(N__57420));
    Span4Mux_h I__12986 (
            .O(N__57423),
            .I(N__57417));
    LocalMux I__12985 (
            .O(N__57420),
            .I(\c0.data_in_frame_15_7 ));
    Odrv4 I__12984 (
            .O(N__57417),
            .I(\c0.data_in_frame_15_7 ));
    InMux I__12983 (
            .O(N__57412),
            .I(N__57409));
    LocalMux I__12982 (
            .O(N__57409),
            .I(N__57405));
    CascadeMux I__12981 (
            .O(N__57408),
            .I(N__57402));
    Span4Mux_h I__12980 (
            .O(N__57405),
            .I(N__57398));
    InMux I__12979 (
            .O(N__57402),
            .I(N__57395));
    InMux I__12978 (
            .O(N__57401),
            .I(N__57392));
    Span4Mux_h I__12977 (
            .O(N__57398),
            .I(N__57389));
    LocalMux I__12976 (
            .O(N__57395),
            .I(N__57384));
    LocalMux I__12975 (
            .O(N__57392),
            .I(N__57384));
    Odrv4 I__12974 (
            .O(N__57389),
            .I(\c0.data_in_frame_14_2 ));
    Odrv4 I__12973 (
            .O(N__57384),
            .I(\c0.data_in_frame_14_2 ));
    CascadeMux I__12972 (
            .O(N__57379),
            .I(N__57376));
    InMux I__12971 (
            .O(N__57376),
            .I(N__57373));
    LocalMux I__12970 (
            .O(N__57373),
            .I(N__57368));
    InMux I__12969 (
            .O(N__57372),
            .I(N__57365));
    InMux I__12968 (
            .O(N__57371),
            .I(N__57362));
    Span4Mux_h I__12967 (
            .O(N__57368),
            .I(N__57358));
    LocalMux I__12966 (
            .O(N__57365),
            .I(N__57355));
    LocalMux I__12965 (
            .O(N__57362),
            .I(N__57352));
    InMux I__12964 (
            .O(N__57361),
            .I(N__57349));
    Span4Mux_v I__12963 (
            .O(N__57358),
            .I(N__57346));
    Span4Mux_h I__12962 (
            .O(N__57355),
            .I(N__57343));
    Span4Mux_h I__12961 (
            .O(N__57352),
            .I(N__57340));
    LocalMux I__12960 (
            .O(N__57349),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__12959 (
            .O(N__57346),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__12958 (
            .O(N__57343),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__12957 (
            .O(N__57340),
            .I(\c0.data_in_frame_7_2 ));
    InMux I__12956 (
            .O(N__57331),
            .I(N__57325));
    InMux I__12955 (
            .O(N__57330),
            .I(N__57322));
    InMux I__12954 (
            .O(N__57329),
            .I(N__57317));
    InMux I__12953 (
            .O(N__57328),
            .I(N__57317));
    LocalMux I__12952 (
            .O(N__57325),
            .I(N__57314));
    LocalMux I__12951 (
            .O(N__57322),
            .I(N__57309));
    LocalMux I__12950 (
            .O(N__57317),
            .I(N__57309));
    Span4Mux_v I__12949 (
            .O(N__57314),
            .I(N__57302));
    Span4Mux_v I__12948 (
            .O(N__57309),
            .I(N__57302));
    InMux I__12947 (
            .O(N__57308),
            .I(N__57299));
    InMux I__12946 (
            .O(N__57307),
            .I(N__57296));
    Odrv4 I__12945 (
            .O(N__57302),
            .I(\c0.n20981 ));
    LocalMux I__12944 (
            .O(N__57299),
            .I(\c0.n20981 ));
    LocalMux I__12943 (
            .O(N__57296),
            .I(\c0.n20981 ));
    InMux I__12942 (
            .O(N__57289),
            .I(N__57286));
    LocalMux I__12941 (
            .O(N__57286),
            .I(N__57283));
    Span4Mux_h I__12940 (
            .O(N__57283),
            .I(N__57280));
    Span4Mux_v I__12939 (
            .O(N__57280),
            .I(N__57277));
    Span4Mux_h I__12938 (
            .O(N__57277),
            .I(N__57274));
    Odrv4 I__12937 (
            .O(N__57274),
            .I(\c0.n25_adj_3157 ));
    InMux I__12936 (
            .O(N__57271),
            .I(N__57268));
    LocalMux I__12935 (
            .O(N__57268),
            .I(N__57264));
    InMux I__12934 (
            .O(N__57267),
            .I(N__57261));
    Odrv4 I__12933 (
            .O(N__57264),
            .I(\c0.n5753 ));
    LocalMux I__12932 (
            .O(N__57261),
            .I(\c0.n5753 ));
    CascadeMux I__12931 (
            .O(N__57256),
            .I(N__57252));
    InMux I__12930 (
            .O(N__57255),
            .I(N__57248));
    InMux I__12929 (
            .O(N__57252),
            .I(N__57245));
    CascadeMux I__12928 (
            .O(N__57251),
            .I(N__57242));
    LocalMux I__12927 (
            .O(N__57248),
            .I(N__57239));
    LocalMux I__12926 (
            .O(N__57245),
            .I(N__57236));
    InMux I__12925 (
            .O(N__57242),
            .I(N__57232));
    Sp12to4 I__12924 (
            .O(N__57239),
            .I(N__57229));
    Span4Mux_h I__12923 (
            .O(N__57236),
            .I(N__57226));
    CascadeMux I__12922 (
            .O(N__57235),
            .I(N__57222));
    LocalMux I__12921 (
            .O(N__57232),
            .I(N__57219));
    Span12Mux_v I__12920 (
            .O(N__57229),
            .I(N__57216));
    Span4Mux_v I__12919 (
            .O(N__57226),
            .I(N__57213));
    InMux I__12918 (
            .O(N__57225),
            .I(N__57208));
    InMux I__12917 (
            .O(N__57222),
            .I(N__57208));
    Span4Mux_h I__12916 (
            .O(N__57219),
            .I(N__57205));
    Odrv12 I__12915 (
            .O(N__57216),
            .I(\c0.data_in_frame_14_0 ));
    Odrv4 I__12914 (
            .O(N__57213),
            .I(\c0.data_in_frame_14_0 ));
    LocalMux I__12913 (
            .O(N__57208),
            .I(\c0.data_in_frame_14_0 ));
    Odrv4 I__12912 (
            .O(N__57205),
            .I(\c0.data_in_frame_14_0 ));
    InMux I__12911 (
            .O(N__57196),
            .I(N__57192));
    CascadeMux I__12910 (
            .O(N__57195),
            .I(N__57188));
    LocalMux I__12909 (
            .O(N__57192),
            .I(N__57184));
    InMux I__12908 (
            .O(N__57191),
            .I(N__57181));
    InMux I__12907 (
            .O(N__57188),
            .I(N__57178));
    InMux I__12906 (
            .O(N__57187),
            .I(N__57175));
    Span4Mux_v I__12905 (
            .O(N__57184),
            .I(N__57170));
    LocalMux I__12904 (
            .O(N__57181),
            .I(N__57170));
    LocalMux I__12903 (
            .O(N__57178),
            .I(N__57165));
    LocalMux I__12902 (
            .O(N__57175),
            .I(N__57165));
    Span4Mux_v I__12901 (
            .O(N__57170),
            .I(N__57162));
    Odrv4 I__12900 (
            .O(N__57165),
            .I(\c0.data_in_frame_12_0 ));
    Odrv4 I__12899 (
            .O(N__57162),
            .I(\c0.data_in_frame_12_0 ));
    InMux I__12898 (
            .O(N__57157),
            .I(N__57154));
    LocalMux I__12897 (
            .O(N__57154),
            .I(N__57149));
    InMux I__12896 (
            .O(N__57153),
            .I(N__57144));
    InMux I__12895 (
            .O(N__57152),
            .I(N__57144));
    Span4Mux_v I__12894 (
            .O(N__57149),
            .I(N__57139));
    LocalMux I__12893 (
            .O(N__57144),
            .I(N__57136));
    InMux I__12892 (
            .O(N__57143),
            .I(N__57133));
    InMux I__12891 (
            .O(N__57142),
            .I(N__57130));
    Odrv4 I__12890 (
            .O(N__57139),
            .I(\c0.n20055 ));
    Odrv4 I__12889 (
            .O(N__57136),
            .I(\c0.n20055 ));
    LocalMux I__12888 (
            .O(N__57133),
            .I(\c0.n20055 ));
    LocalMux I__12887 (
            .O(N__57130),
            .I(\c0.n20055 ));
    CascadeMux I__12886 (
            .O(N__57121),
            .I(\c0.n20_adj_3536_cascade_ ));
    CascadeMux I__12885 (
            .O(N__57118),
            .I(\c0.n12_adj_3558_cascade_ ));
    InMux I__12884 (
            .O(N__57115),
            .I(N__57111));
    CascadeMux I__12883 (
            .O(N__57114),
            .I(N__57108));
    LocalMux I__12882 (
            .O(N__57111),
            .I(N__57104));
    InMux I__12881 (
            .O(N__57108),
            .I(N__57098));
    InMux I__12880 (
            .O(N__57107),
            .I(N__57098));
    Span4Mux_v I__12879 (
            .O(N__57104),
            .I(N__57095));
    InMux I__12878 (
            .O(N__57103),
            .I(N__57092));
    LocalMux I__12877 (
            .O(N__57098),
            .I(N__57084));
    Span4Mux_h I__12876 (
            .O(N__57095),
            .I(N__57084));
    LocalMux I__12875 (
            .O(N__57092),
            .I(N__57084));
    InMux I__12874 (
            .O(N__57091),
            .I(N__57081));
    Odrv4 I__12873 (
            .O(N__57084),
            .I(\c0.data_in_frame_8_5 ));
    LocalMux I__12872 (
            .O(N__57081),
            .I(\c0.data_in_frame_8_5 ));
    CascadeMux I__12871 (
            .O(N__57076),
            .I(N__57072));
    InMux I__12870 (
            .O(N__57075),
            .I(N__57068));
    InMux I__12869 (
            .O(N__57072),
            .I(N__57065));
    InMux I__12868 (
            .O(N__57071),
            .I(N__57062));
    LocalMux I__12867 (
            .O(N__57068),
            .I(N__57059));
    LocalMux I__12866 (
            .O(N__57065),
            .I(N__57056));
    LocalMux I__12865 (
            .O(N__57062),
            .I(N__57051));
    Span4Mux_h I__12864 (
            .O(N__57059),
            .I(N__57051));
    Odrv12 I__12863 (
            .O(N__57056),
            .I(\c0.data_in_frame_12_7 ));
    Odrv4 I__12862 (
            .O(N__57051),
            .I(\c0.data_in_frame_12_7 ));
    InMux I__12861 (
            .O(N__57046),
            .I(N__57040));
    InMux I__12860 (
            .O(N__57045),
            .I(N__57037));
    InMux I__12859 (
            .O(N__57044),
            .I(N__57034));
    InMux I__12858 (
            .O(N__57043),
            .I(N__57031));
    LocalMux I__12857 (
            .O(N__57040),
            .I(N__57028));
    LocalMux I__12856 (
            .O(N__57037),
            .I(N__57025));
    LocalMux I__12855 (
            .O(N__57034),
            .I(N__57021));
    LocalMux I__12854 (
            .O(N__57031),
            .I(N__57018));
    Span4Mux_h I__12853 (
            .O(N__57028),
            .I(N__57013));
    Span4Mux_h I__12852 (
            .O(N__57025),
            .I(N__57013));
    InMux I__12851 (
            .O(N__57024),
            .I(N__57010));
    Span4Mux_h I__12850 (
            .O(N__57021),
            .I(N__57007));
    Span4Mux_h I__12849 (
            .O(N__57018),
            .I(N__57001));
    Span4Mux_v I__12848 (
            .O(N__57013),
            .I(N__56998));
    LocalMux I__12847 (
            .O(N__57010),
            .I(N__56993));
    Sp12to4 I__12846 (
            .O(N__57007),
            .I(N__56993));
    InMux I__12845 (
            .O(N__57006),
            .I(N__56988));
    InMux I__12844 (
            .O(N__57005),
            .I(N__56988));
    InMux I__12843 (
            .O(N__57004),
            .I(N__56985));
    Odrv4 I__12842 (
            .O(N__57001),
            .I(\c0.n5_adj_3031 ));
    Odrv4 I__12841 (
            .O(N__56998),
            .I(\c0.n5_adj_3031 ));
    Odrv12 I__12840 (
            .O(N__56993),
            .I(\c0.n5_adj_3031 ));
    LocalMux I__12839 (
            .O(N__56988),
            .I(\c0.n5_adj_3031 ));
    LocalMux I__12838 (
            .O(N__56985),
            .I(\c0.n5_adj_3031 ));
    CascadeMux I__12837 (
            .O(N__56974),
            .I(\c0.n19359_cascade_ ));
    CascadeMux I__12836 (
            .O(N__56971),
            .I(N__56967));
    InMux I__12835 (
            .O(N__56970),
            .I(N__56964));
    InMux I__12834 (
            .O(N__56967),
            .I(N__56961));
    LocalMux I__12833 (
            .O(N__56964),
            .I(N__56958));
    LocalMux I__12832 (
            .O(N__56961),
            .I(N__56954));
    Span4Mux_h I__12831 (
            .O(N__56958),
            .I(N__56951));
    InMux I__12830 (
            .O(N__56957),
            .I(N__56948));
    Odrv4 I__12829 (
            .O(N__56954),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__12828 (
            .O(N__56951),
            .I(\c0.data_in_frame_8_4 ));
    LocalMux I__12827 (
            .O(N__56948),
            .I(\c0.data_in_frame_8_4 ));
    InMux I__12826 (
            .O(N__56941),
            .I(N__56933));
    InMux I__12825 (
            .O(N__56940),
            .I(N__56933));
    InMux I__12824 (
            .O(N__56939),
            .I(N__56930));
    InMux I__12823 (
            .O(N__56938),
            .I(N__56927));
    LocalMux I__12822 (
            .O(N__56933),
            .I(N__56922));
    LocalMux I__12821 (
            .O(N__56930),
            .I(N__56922));
    LocalMux I__12820 (
            .O(N__56927),
            .I(\c0.n11478 ));
    Odrv12 I__12819 (
            .O(N__56922),
            .I(\c0.n11478 ));
    InMux I__12818 (
            .O(N__56917),
            .I(N__56914));
    LocalMux I__12817 (
            .O(N__56914),
            .I(\c0.n19199 ));
    InMux I__12816 (
            .O(N__56911),
            .I(N__56908));
    LocalMux I__12815 (
            .O(N__56908),
            .I(N__56905));
    Span4Mux_h I__12814 (
            .O(N__56905),
            .I(N__56899));
    InMux I__12813 (
            .O(N__56904),
            .I(N__56896));
    InMux I__12812 (
            .O(N__56903),
            .I(N__56891));
    InMux I__12811 (
            .O(N__56902),
            .I(N__56891));
    Span4Mux_h I__12810 (
            .O(N__56899),
            .I(N__56888));
    LocalMux I__12809 (
            .O(N__56896),
            .I(\c0.data_in_frame_10_5 ));
    LocalMux I__12808 (
            .O(N__56891),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__12807 (
            .O(N__56888),
            .I(\c0.data_in_frame_10_5 ));
    CascadeMux I__12806 (
            .O(N__56881),
            .I(\c0.n19199_cascade_ ));
    CascadeMux I__12805 (
            .O(N__56878),
            .I(N__56875));
    InMux I__12804 (
            .O(N__56875),
            .I(N__56872));
    LocalMux I__12803 (
            .O(N__56872),
            .I(N__56869));
    Span4Mux_h I__12802 (
            .O(N__56869),
            .I(N__56866));
    Span4Mux_h I__12801 (
            .O(N__56866),
            .I(N__56863));
    Odrv4 I__12800 (
            .O(N__56863),
            .I(\c0.n19_adj_3540 ));
    CascadeMux I__12799 (
            .O(N__56860),
            .I(N__56857));
    InMux I__12798 (
            .O(N__56857),
            .I(N__56854));
    LocalMux I__12797 (
            .O(N__56854),
            .I(N__56849));
    InMux I__12796 (
            .O(N__56853),
            .I(N__56843));
    InMux I__12795 (
            .O(N__56852),
            .I(N__56840));
    Span4Mux_h I__12794 (
            .O(N__56849),
            .I(N__56837));
    InMux I__12793 (
            .O(N__56848),
            .I(N__56834));
    InMux I__12792 (
            .O(N__56847),
            .I(N__56831));
    InMux I__12791 (
            .O(N__56846),
            .I(N__56826));
    LocalMux I__12790 (
            .O(N__56843),
            .I(N__56818));
    LocalMux I__12789 (
            .O(N__56840),
            .I(N__56818));
    Span4Mux_h I__12788 (
            .O(N__56837),
            .I(N__56811));
    LocalMux I__12787 (
            .O(N__56834),
            .I(N__56811));
    LocalMux I__12786 (
            .O(N__56831),
            .I(N__56811));
    CascadeMux I__12785 (
            .O(N__56830),
            .I(N__56807));
    CascadeMux I__12784 (
            .O(N__56829),
            .I(N__56804));
    LocalMux I__12783 (
            .O(N__56826),
            .I(N__56797));
    InMux I__12782 (
            .O(N__56825),
            .I(N__56794));
    InMux I__12781 (
            .O(N__56824),
            .I(N__56791));
    InMux I__12780 (
            .O(N__56823),
            .I(N__56788));
    Span4Mux_h I__12779 (
            .O(N__56818),
            .I(N__56783));
    Span4Mux_h I__12778 (
            .O(N__56811),
            .I(N__56783));
    InMux I__12777 (
            .O(N__56810),
            .I(N__56776));
    InMux I__12776 (
            .O(N__56807),
            .I(N__56776));
    InMux I__12775 (
            .O(N__56804),
            .I(N__56776));
    InMux I__12774 (
            .O(N__56803),
            .I(N__56771));
    InMux I__12773 (
            .O(N__56802),
            .I(N__56771));
    InMux I__12772 (
            .O(N__56801),
            .I(N__56768));
    InMux I__12771 (
            .O(N__56800),
            .I(N__56765));
    Span4Mux_h I__12770 (
            .O(N__56797),
            .I(N__56758));
    LocalMux I__12769 (
            .O(N__56794),
            .I(N__56758));
    LocalMux I__12768 (
            .O(N__56791),
            .I(N__56758));
    LocalMux I__12767 (
            .O(N__56788),
            .I(data_in_frame_0_1));
    Odrv4 I__12766 (
            .O(N__56783),
            .I(data_in_frame_0_1));
    LocalMux I__12765 (
            .O(N__56776),
            .I(data_in_frame_0_1));
    LocalMux I__12764 (
            .O(N__56771),
            .I(data_in_frame_0_1));
    LocalMux I__12763 (
            .O(N__56768),
            .I(data_in_frame_0_1));
    LocalMux I__12762 (
            .O(N__56765),
            .I(data_in_frame_0_1));
    Odrv4 I__12761 (
            .O(N__56758),
            .I(data_in_frame_0_1));
    InMux I__12760 (
            .O(N__56743),
            .I(N__56740));
    LocalMux I__12759 (
            .O(N__56740),
            .I(N__56737));
    Span4Mux_h I__12758 (
            .O(N__56737),
            .I(N__56734));
    Odrv4 I__12757 (
            .O(N__56734),
            .I(\c0.n17_adj_3544 ));
    CascadeMux I__12756 (
            .O(N__56731),
            .I(N__56728));
    InMux I__12755 (
            .O(N__56728),
            .I(N__56723));
    InMux I__12754 (
            .O(N__56727),
            .I(N__56720));
    InMux I__12753 (
            .O(N__56726),
            .I(N__56716));
    LocalMux I__12752 (
            .O(N__56723),
            .I(N__56711));
    LocalMux I__12751 (
            .O(N__56720),
            .I(N__56711));
    InMux I__12750 (
            .O(N__56719),
            .I(N__56708));
    LocalMux I__12749 (
            .O(N__56716),
            .I(N__56704));
    Span4Mux_h I__12748 (
            .O(N__56711),
            .I(N__56700));
    LocalMux I__12747 (
            .O(N__56708),
            .I(N__56697));
    InMux I__12746 (
            .O(N__56707),
            .I(N__56694));
    Span4Mux_h I__12745 (
            .O(N__56704),
            .I(N__56691));
    InMux I__12744 (
            .O(N__56703),
            .I(N__56688));
    Span4Mux_h I__12743 (
            .O(N__56700),
            .I(N__56685));
    Span4Mux_h I__12742 (
            .O(N__56697),
            .I(N__56682));
    LocalMux I__12741 (
            .O(N__56694),
            .I(\c0.data_in_frame_9_1 ));
    Odrv4 I__12740 (
            .O(N__56691),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__12739 (
            .O(N__56688),
            .I(\c0.data_in_frame_9_1 ));
    Odrv4 I__12738 (
            .O(N__56685),
            .I(\c0.data_in_frame_9_1 ));
    Odrv4 I__12737 (
            .O(N__56682),
            .I(\c0.data_in_frame_9_1 ));
    CascadeMux I__12736 (
            .O(N__56671),
            .I(\c0.n11858_cascade_ ));
    InMux I__12735 (
            .O(N__56668),
            .I(N__56665));
    LocalMux I__12734 (
            .O(N__56665),
            .I(N__56662));
    Span4Mux_v I__12733 (
            .O(N__56662),
            .I(N__56659));
    Odrv4 I__12732 (
            .O(N__56659),
            .I(\c0.n19446 ));
    CascadeMux I__12731 (
            .O(N__56656),
            .I(\c0.n19446_cascade_ ));
    InMux I__12730 (
            .O(N__56653),
            .I(N__56647));
    InMux I__12729 (
            .O(N__56652),
            .I(N__56643));
    InMux I__12728 (
            .O(N__56651),
            .I(N__56637));
    InMux I__12727 (
            .O(N__56650),
            .I(N__56637));
    LocalMux I__12726 (
            .O(N__56647),
            .I(N__56634));
    InMux I__12725 (
            .O(N__56646),
            .I(N__56631));
    LocalMux I__12724 (
            .O(N__56643),
            .I(N__56626));
    InMux I__12723 (
            .O(N__56642),
            .I(N__56623));
    LocalMux I__12722 (
            .O(N__56637),
            .I(N__56620));
    Span4Mux_v I__12721 (
            .O(N__56634),
            .I(N__56617));
    LocalMux I__12720 (
            .O(N__56631),
            .I(N__56614));
    InMux I__12719 (
            .O(N__56630),
            .I(N__56611));
    InMux I__12718 (
            .O(N__56629),
            .I(N__56608));
    Span4Mux_v I__12717 (
            .O(N__56626),
            .I(N__56605));
    LocalMux I__12716 (
            .O(N__56623),
            .I(N__56602));
    Span4Mux_v I__12715 (
            .O(N__56620),
            .I(N__56599));
    Span4Mux_h I__12714 (
            .O(N__56617),
            .I(N__56594));
    Span4Mux_v I__12713 (
            .O(N__56614),
            .I(N__56594));
    LocalMux I__12712 (
            .O(N__56611),
            .I(N__56591));
    LocalMux I__12711 (
            .O(N__56608),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    Odrv4 I__12710 (
            .O(N__56605),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    Odrv4 I__12709 (
            .O(N__56602),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    Odrv4 I__12708 (
            .O(N__56599),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    Odrv4 I__12707 (
            .O(N__56594),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    Odrv12 I__12706 (
            .O(N__56591),
            .I(\c0.data_out_frame_0__7__N_1537 ));
    InMux I__12705 (
            .O(N__56578),
            .I(N__56575));
    LocalMux I__12704 (
            .O(N__56575),
            .I(N__56572));
    Odrv12 I__12703 (
            .O(N__56572),
            .I(\c0.n11982 ));
    CascadeMux I__12702 (
            .O(N__56569),
            .I(\c0.n33_adj_3209_cascade_ ));
    InMux I__12701 (
            .O(N__56566),
            .I(N__56563));
    LocalMux I__12700 (
            .O(N__56563),
            .I(N__56557));
    InMux I__12699 (
            .O(N__56562),
            .I(N__56552));
    InMux I__12698 (
            .O(N__56561),
            .I(N__56552));
    InMux I__12697 (
            .O(N__56560),
            .I(N__56549));
    Span4Mux_v I__12696 (
            .O(N__56557),
            .I(N__56546));
    LocalMux I__12695 (
            .O(N__56552),
            .I(N__56543));
    LocalMux I__12694 (
            .O(N__56549),
            .I(N__56540));
    Odrv4 I__12693 (
            .O(N__56546),
            .I(\c0.n5598 ));
    Odrv4 I__12692 (
            .O(N__56543),
            .I(\c0.n5598 ));
    Odrv4 I__12691 (
            .O(N__56540),
            .I(\c0.n5598 ));
    CascadeMux I__12690 (
            .O(N__56533),
            .I(N__56530));
    InMux I__12689 (
            .O(N__56530),
            .I(N__56525));
    InMux I__12688 (
            .O(N__56529),
            .I(N__56521));
    InMux I__12687 (
            .O(N__56528),
            .I(N__56518));
    LocalMux I__12686 (
            .O(N__56525),
            .I(N__56515));
    CascadeMux I__12685 (
            .O(N__56524),
            .I(N__56512));
    LocalMux I__12684 (
            .O(N__56521),
            .I(N__56509));
    LocalMux I__12683 (
            .O(N__56518),
            .I(N__56504));
    Span4Mux_h I__12682 (
            .O(N__56515),
            .I(N__56504));
    InMux I__12681 (
            .O(N__56512),
            .I(N__56501));
    Span12Mux_h I__12680 (
            .O(N__56509),
            .I(N__56498));
    Span4Mux_v I__12679 (
            .O(N__56504),
            .I(N__56495));
    LocalMux I__12678 (
            .O(N__56501),
            .I(\c0.data_in_frame_17_7 ));
    Odrv12 I__12677 (
            .O(N__56498),
            .I(\c0.data_in_frame_17_7 ));
    Odrv4 I__12676 (
            .O(N__56495),
            .I(\c0.data_in_frame_17_7 ));
    InMux I__12675 (
            .O(N__56488),
            .I(N__56485));
    LocalMux I__12674 (
            .O(N__56485),
            .I(N__56481));
    InMux I__12673 (
            .O(N__56484),
            .I(N__56478));
    Span4Mux_v I__12672 (
            .O(N__56481),
            .I(N__56475));
    LocalMux I__12671 (
            .O(N__56478),
            .I(\c0.n9_adj_3350 ));
    Odrv4 I__12670 (
            .O(N__56475),
            .I(\c0.n9_adj_3350 ));
    InMux I__12669 (
            .O(N__56470),
            .I(N__56467));
    LocalMux I__12668 (
            .O(N__56467),
            .I(N__56464));
    Span4Mux_v I__12667 (
            .O(N__56464),
            .I(N__56461));
    Odrv4 I__12666 (
            .O(N__56461),
            .I(\c0.n29_adj_3533 ));
    InMux I__12665 (
            .O(N__56458),
            .I(N__56455));
    LocalMux I__12664 (
            .O(N__56455),
            .I(\c0.n33_adj_3209 ));
    CascadeMux I__12663 (
            .O(N__56452),
            .I(N__56447));
    InMux I__12662 (
            .O(N__56451),
            .I(N__56442));
    InMux I__12661 (
            .O(N__56450),
            .I(N__56442));
    InMux I__12660 (
            .O(N__56447),
            .I(N__56437));
    LocalMux I__12659 (
            .O(N__56442),
            .I(N__56434));
    InMux I__12658 (
            .O(N__56441),
            .I(N__56429));
    InMux I__12657 (
            .O(N__56440),
            .I(N__56429));
    LocalMux I__12656 (
            .O(N__56437),
            .I(N__56426));
    Span4Mux_h I__12655 (
            .O(N__56434),
            .I(N__56421));
    LocalMux I__12654 (
            .O(N__56429),
            .I(N__56421));
    Span4Mux_v I__12653 (
            .O(N__56426),
            .I(N__56418));
    Span4Mux_v I__12652 (
            .O(N__56421),
            .I(N__56413));
    Span4Mux_h I__12651 (
            .O(N__56418),
            .I(N__56413));
    Odrv4 I__12650 (
            .O(N__56413),
            .I(\c0.n12209 ));
    InMux I__12649 (
            .O(N__56410),
            .I(N__56406));
    InMux I__12648 (
            .O(N__56409),
            .I(N__56403));
    LocalMux I__12647 (
            .O(N__56406),
            .I(N__56400));
    LocalMux I__12646 (
            .O(N__56403),
            .I(N__56393));
    Span4Mux_h I__12645 (
            .O(N__56400),
            .I(N__56393));
    InMux I__12644 (
            .O(N__56399),
            .I(N__56390));
    InMux I__12643 (
            .O(N__56398),
            .I(N__56387));
    Span4Mux_v I__12642 (
            .O(N__56393),
            .I(N__56384));
    LocalMux I__12641 (
            .O(N__56390),
            .I(N__56379));
    LocalMux I__12640 (
            .O(N__56387),
            .I(N__56379));
    Span4Mux_v I__12639 (
            .O(N__56384),
            .I(N__56373));
    Span4Mux_v I__12638 (
            .O(N__56379),
            .I(N__56373));
    InMux I__12637 (
            .O(N__56378),
            .I(N__56370));
    Odrv4 I__12636 (
            .O(N__56373),
            .I(\c0.n9_adj_3027 ));
    LocalMux I__12635 (
            .O(N__56370),
            .I(\c0.n9_adj_3027 ));
    InMux I__12634 (
            .O(N__56365),
            .I(N__56362));
    LocalMux I__12633 (
            .O(N__56362),
            .I(\c0.n45_adj_3224 ));
    CascadeMux I__12632 (
            .O(N__56359),
            .I(N__56356));
    InMux I__12631 (
            .O(N__56356),
            .I(N__56353));
    LocalMux I__12630 (
            .O(N__56353),
            .I(N__56348));
    InMux I__12629 (
            .O(N__56352),
            .I(N__56345));
    CascadeMux I__12628 (
            .O(N__56351),
            .I(N__56342));
    Span4Mux_h I__12627 (
            .O(N__56348),
            .I(N__56338));
    LocalMux I__12626 (
            .O(N__56345),
            .I(N__56335));
    InMux I__12625 (
            .O(N__56342),
            .I(N__56332));
    InMux I__12624 (
            .O(N__56341),
            .I(N__56329));
    Span4Mux_h I__12623 (
            .O(N__56338),
            .I(N__56326));
    Span4Mux_h I__12622 (
            .O(N__56335),
            .I(N__56323));
    LocalMux I__12621 (
            .O(N__56332),
            .I(\c0.data_in_frame_7_6 ));
    LocalMux I__12620 (
            .O(N__56329),
            .I(\c0.data_in_frame_7_6 ));
    Odrv4 I__12619 (
            .O(N__56326),
            .I(\c0.data_in_frame_7_6 ));
    Odrv4 I__12618 (
            .O(N__56323),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__12617 (
            .O(N__56314),
            .I(N__56308));
    InMux I__12616 (
            .O(N__56313),
            .I(N__56308));
    LocalMux I__12615 (
            .O(N__56308),
            .I(N__56305));
    Sp12to4 I__12614 (
            .O(N__56305),
            .I(N__56302));
    Odrv12 I__12613 (
            .O(N__56302),
            .I(\c0.n15 ));
    InMux I__12612 (
            .O(N__56299),
            .I(N__56296));
    LocalMux I__12611 (
            .O(N__56296),
            .I(N__56292));
    InMux I__12610 (
            .O(N__56295),
            .I(N__56287));
    Span4Mux_h I__12609 (
            .O(N__56292),
            .I(N__56284));
    InMux I__12608 (
            .O(N__56291),
            .I(N__56279));
    InMux I__12607 (
            .O(N__56290),
            .I(N__56279));
    LocalMux I__12606 (
            .O(N__56287),
            .I(\c0.n23 ));
    Odrv4 I__12605 (
            .O(N__56284),
            .I(\c0.n23 ));
    LocalMux I__12604 (
            .O(N__56279),
            .I(\c0.n23 ));
    InMux I__12603 (
            .O(N__56272),
            .I(N__56269));
    LocalMux I__12602 (
            .O(N__56269),
            .I(\c0.n51_adj_3426 ));
    InMux I__12601 (
            .O(N__56266),
            .I(N__56263));
    LocalMux I__12600 (
            .O(N__56263),
            .I(N__56260));
    Span4Mux_v I__12599 (
            .O(N__56260),
            .I(N__56256));
    InMux I__12598 (
            .O(N__56259),
            .I(N__56253));
    Span4Mux_h I__12597 (
            .O(N__56256),
            .I(N__56248));
    LocalMux I__12596 (
            .O(N__56253),
            .I(N__56248));
    Span4Mux_h I__12595 (
            .O(N__56248),
            .I(N__56245));
    Span4Mux_v I__12594 (
            .O(N__56245),
            .I(N__56242));
    Odrv4 I__12593 (
            .O(N__56242),
            .I(n15645));
    CascadeMux I__12592 (
            .O(N__56239),
            .I(N__56233));
    CascadeMux I__12591 (
            .O(N__56238),
            .I(N__56230));
    CascadeMux I__12590 (
            .O(N__56237),
            .I(N__56227));
    CascadeMux I__12589 (
            .O(N__56236),
            .I(N__56221));
    InMux I__12588 (
            .O(N__56233),
            .I(N__56214));
    InMux I__12587 (
            .O(N__56230),
            .I(N__56214));
    InMux I__12586 (
            .O(N__56227),
            .I(N__56214));
    CascadeMux I__12585 (
            .O(N__56226),
            .I(N__56210));
    CascadeMux I__12584 (
            .O(N__56225),
            .I(N__56207));
    CascadeMux I__12583 (
            .O(N__56224),
            .I(N__56204));
    InMux I__12582 (
            .O(N__56221),
            .I(N__56201));
    LocalMux I__12581 (
            .O(N__56214),
            .I(N__56197));
    InMux I__12580 (
            .O(N__56213),
            .I(N__56194));
    InMux I__12579 (
            .O(N__56210),
            .I(N__56188));
    InMux I__12578 (
            .O(N__56207),
            .I(N__56188));
    InMux I__12577 (
            .O(N__56204),
            .I(N__56185));
    LocalMux I__12576 (
            .O(N__56201),
            .I(N__56182));
    InMux I__12575 (
            .O(N__56200),
            .I(N__56179));
    Span4Mux_h I__12574 (
            .O(N__56197),
            .I(N__56176));
    LocalMux I__12573 (
            .O(N__56194),
            .I(N__56173));
    InMux I__12572 (
            .O(N__56193),
            .I(N__56170));
    LocalMux I__12571 (
            .O(N__56188),
            .I(N__56167));
    LocalMux I__12570 (
            .O(N__56185),
            .I(N__56164));
    Sp12to4 I__12569 (
            .O(N__56182),
            .I(N__56161));
    LocalMux I__12568 (
            .O(N__56179),
            .I(N__56158));
    Span4Mux_v I__12567 (
            .O(N__56176),
            .I(N__56155));
    Span4Mux_h I__12566 (
            .O(N__56173),
            .I(N__56149));
    LocalMux I__12565 (
            .O(N__56170),
            .I(N__56149));
    Span4Mux_v I__12564 (
            .O(N__56167),
            .I(N__56146));
    Span4Mux_v I__12563 (
            .O(N__56164),
            .I(N__56143));
    Span12Mux_s10_v I__12562 (
            .O(N__56161),
            .I(N__56140));
    Span4Mux_v I__12561 (
            .O(N__56158),
            .I(N__56135));
    Span4Mux_v I__12560 (
            .O(N__56155),
            .I(N__56135));
    InMux I__12559 (
            .O(N__56154),
            .I(N__56132));
    Span4Mux_v I__12558 (
            .O(N__56149),
            .I(N__56127));
    Span4Mux_h I__12557 (
            .O(N__56146),
            .I(N__56127));
    Sp12to4 I__12556 (
            .O(N__56143),
            .I(N__56123));
    Span12Mux_h I__12555 (
            .O(N__56140),
            .I(N__56120));
    Span4Mux_h I__12554 (
            .O(N__56135),
            .I(N__56117));
    LocalMux I__12553 (
            .O(N__56132),
            .I(N__56114));
    Sp12to4 I__12552 (
            .O(N__56127),
            .I(N__56111));
    InMux I__12551 (
            .O(N__56126),
            .I(N__56108));
    Span12Mux_s9_v I__12550 (
            .O(N__56123),
            .I(N__56103));
    Span12Mux_v I__12549 (
            .O(N__56120),
            .I(N__56103));
    Span4Mux_v I__12548 (
            .O(N__56117),
            .I(N__56098));
    Span4Mux_h I__12547 (
            .O(N__56114),
            .I(N__56098));
    Span12Mux_h I__12546 (
            .O(N__56111),
            .I(N__56093));
    LocalMux I__12545 (
            .O(N__56108),
            .I(N__56093));
    Odrv12 I__12544 (
            .O(N__56103),
            .I(r_Rx_Data));
    Odrv4 I__12543 (
            .O(N__56098),
            .I(r_Rx_Data));
    Odrv12 I__12542 (
            .O(N__56093),
            .I(r_Rx_Data));
    InMux I__12541 (
            .O(N__56086),
            .I(N__56081));
    InMux I__12540 (
            .O(N__56085),
            .I(N__56077));
    InMux I__12539 (
            .O(N__56084),
            .I(N__56074));
    LocalMux I__12538 (
            .O(N__56081),
            .I(N__56071));
    CascadeMux I__12537 (
            .O(N__56080),
            .I(N__56068));
    LocalMux I__12536 (
            .O(N__56077),
            .I(N__56065));
    LocalMux I__12535 (
            .O(N__56074),
            .I(N__56062));
    Span4Mux_h I__12534 (
            .O(N__56071),
            .I(N__56059));
    InMux I__12533 (
            .O(N__56068),
            .I(N__56056));
    Span4Mux_v I__12532 (
            .O(N__56065),
            .I(N__56053));
    Span4Mux_h I__12531 (
            .O(N__56062),
            .I(N__56048));
    Span4Mux_h I__12530 (
            .O(N__56059),
            .I(N__56048));
    LocalMux I__12529 (
            .O(N__56056),
            .I(N__56043));
    Span4Mux_h I__12528 (
            .O(N__56053),
            .I(N__56043));
    Span4Mux_v I__12527 (
            .O(N__56048),
            .I(N__56040));
    Span4Mux_h I__12526 (
            .O(N__56043),
            .I(N__56035));
    Span4Mux_v I__12525 (
            .O(N__56040),
            .I(N__56035));
    Odrv4 I__12524 (
            .O(N__56035),
            .I(n11466));
    InMux I__12523 (
            .O(N__56032),
            .I(N__56029));
    LocalMux I__12522 (
            .O(N__56029),
            .I(N__56024));
    InMux I__12521 (
            .O(N__56028),
            .I(N__56021));
    InMux I__12520 (
            .O(N__56027),
            .I(N__56018));
    Span4Mux_v I__12519 (
            .O(N__56024),
            .I(N__56014));
    LocalMux I__12518 (
            .O(N__56021),
            .I(N__56011));
    LocalMux I__12517 (
            .O(N__56018),
            .I(N__56008));
    CascadeMux I__12516 (
            .O(N__56017),
            .I(N__56005));
    Span4Mux_v I__12515 (
            .O(N__56014),
            .I(N__56002));
    Span4Mux_h I__12514 (
            .O(N__56011),
            .I(N__55999));
    Span4Mux_h I__12513 (
            .O(N__56008),
            .I(N__55996));
    InMux I__12512 (
            .O(N__56005),
            .I(N__55993));
    Span4Mux_h I__12511 (
            .O(N__56002),
            .I(N__55988));
    Span4Mux_v I__12510 (
            .O(N__55999),
            .I(N__55988));
    Span4Mux_h I__12509 (
            .O(N__55996),
            .I(N__55985));
    LocalMux I__12508 (
            .O(N__55993),
            .I(\c0.data_in_frame_13_7 ));
    Odrv4 I__12507 (
            .O(N__55988),
            .I(\c0.data_in_frame_13_7 ));
    Odrv4 I__12506 (
            .O(N__55985),
            .I(\c0.data_in_frame_13_7 ));
    CascadeMux I__12505 (
            .O(N__55978),
            .I(N__55975));
    InMux I__12504 (
            .O(N__55975),
            .I(N__55972));
    LocalMux I__12503 (
            .O(N__55972),
            .I(N__55969));
    Span4Mux_v I__12502 (
            .O(N__55969),
            .I(N__55966));
    Span4Mux_v I__12501 (
            .O(N__55966),
            .I(N__55963));
    Odrv4 I__12500 (
            .O(N__55963),
            .I(\c0.n13_adj_3541 ));
    InMux I__12499 (
            .O(N__55960),
            .I(N__55956));
    CascadeMux I__12498 (
            .O(N__55959),
            .I(N__55953));
    LocalMux I__12497 (
            .O(N__55956),
            .I(N__55948));
    InMux I__12496 (
            .O(N__55953),
            .I(N__55945));
    InMux I__12495 (
            .O(N__55952),
            .I(N__55942));
    CascadeMux I__12494 (
            .O(N__55951),
            .I(N__55939));
    Span4Mux_v I__12493 (
            .O(N__55948),
            .I(N__55932));
    LocalMux I__12492 (
            .O(N__55945),
            .I(N__55932));
    LocalMux I__12491 (
            .O(N__55942),
            .I(N__55932));
    InMux I__12490 (
            .O(N__55939),
            .I(N__55929));
    Span4Mux_v I__12489 (
            .O(N__55932),
            .I(N__55926));
    LocalMux I__12488 (
            .O(N__55929),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__12487 (
            .O(N__55926),
            .I(\c0.data_in_frame_13_2 ));
    InMux I__12486 (
            .O(N__55921),
            .I(N__55916));
    CascadeMux I__12485 (
            .O(N__55920),
            .I(N__55913));
    InMux I__12484 (
            .O(N__55919),
            .I(N__55910));
    LocalMux I__12483 (
            .O(N__55916),
            .I(N__55907));
    InMux I__12482 (
            .O(N__55913),
            .I(N__55904));
    LocalMux I__12481 (
            .O(N__55910),
            .I(N__55901));
    Span4Mux_h I__12480 (
            .O(N__55907),
            .I(N__55898));
    LocalMux I__12479 (
            .O(N__55904),
            .I(N__55893));
    Span4Mux_v I__12478 (
            .O(N__55901),
            .I(N__55893));
    Odrv4 I__12477 (
            .O(N__55898),
            .I(\c0.data_in_frame_9_5 ));
    Odrv4 I__12476 (
            .O(N__55893),
            .I(\c0.data_in_frame_9_5 ));
    InMux I__12475 (
            .O(N__55888),
            .I(N__55880));
    InMux I__12474 (
            .O(N__55887),
            .I(N__55877));
    CascadeMux I__12473 (
            .O(N__55886),
            .I(N__55869));
    InMux I__12472 (
            .O(N__55885),
            .I(N__55862));
    InMux I__12471 (
            .O(N__55884),
            .I(N__55862));
    InMux I__12470 (
            .O(N__55883),
            .I(N__55859));
    LocalMux I__12469 (
            .O(N__55880),
            .I(N__55854));
    LocalMux I__12468 (
            .O(N__55877),
            .I(N__55854));
    InMux I__12467 (
            .O(N__55876),
            .I(N__55849));
    InMux I__12466 (
            .O(N__55875),
            .I(N__55849));
    InMux I__12465 (
            .O(N__55874),
            .I(N__55842));
    InMux I__12464 (
            .O(N__55873),
            .I(N__55842));
    InMux I__12463 (
            .O(N__55872),
            .I(N__55842));
    InMux I__12462 (
            .O(N__55869),
            .I(N__55839));
    CascadeMux I__12461 (
            .O(N__55868),
            .I(N__55836));
    InMux I__12460 (
            .O(N__55867),
            .I(N__55833));
    LocalMux I__12459 (
            .O(N__55862),
            .I(N__55828));
    LocalMux I__12458 (
            .O(N__55859),
            .I(N__55828));
    Span4Mux_h I__12457 (
            .O(N__55854),
            .I(N__55825));
    LocalMux I__12456 (
            .O(N__55849),
            .I(N__55820));
    LocalMux I__12455 (
            .O(N__55842),
            .I(N__55820));
    LocalMux I__12454 (
            .O(N__55839),
            .I(N__55816));
    InMux I__12453 (
            .O(N__55836),
            .I(N__55813));
    LocalMux I__12452 (
            .O(N__55833),
            .I(N__55809));
    Span4Mux_v I__12451 (
            .O(N__55828),
            .I(N__55806));
    Span4Mux_h I__12450 (
            .O(N__55825),
            .I(N__55801));
    Span4Mux_v I__12449 (
            .O(N__55820),
            .I(N__55801));
    CascadeMux I__12448 (
            .O(N__55819),
            .I(N__55797));
    Span4Mux_v I__12447 (
            .O(N__55816),
            .I(N__55792));
    LocalMux I__12446 (
            .O(N__55813),
            .I(N__55789));
    InMux I__12445 (
            .O(N__55812),
            .I(N__55786));
    Span4Mux_h I__12444 (
            .O(N__55809),
            .I(N__55783));
    Span4Mux_h I__12443 (
            .O(N__55806),
            .I(N__55778));
    Span4Mux_v I__12442 (
            .O(N__55801),
            .I(N__55778));
    InMux I__12441 (
            .O(N__55800),
            .I(N__55775));
    InMux I__12440 (
            .O(N__55797),
            .I(N__55768));
    InMux I__12439 (
            .O(N__55796),
            .I(N__55768));
    InMux I__12438 (
            .O(N__55795),
            .I(N__55768));
    Span4Mux_v I__12437 (
            .O(N__55792),
            .I(N__55765));
    Span4Mux_v I__12436 (
            .O(N__55789),
            .I(N__55762));
    LocalMux I__12435 (
            .O(N__55786),
            .I(N__55757));
    Span4Mux_v I__12434 (
            .O(N__55783),
            .I(N__55757));
    Span4Mux_h I__12433 (
            .O(N__55778),
            .I(N__55754));
    LocalMux I__12432 (
            .O(N__55775),
            .I(N__55747));
    LocalMux I__12431 (
            .O(N__55768),
            .I(N__55747));
    Sp12to4 I__12430 (
            .O(N__55765),
            .I(N__55747));
    Span4Mux_h I__12429 (
            .O(N__55762),
            .I(N__55742));
    Span4Mux_v I__12428 (
            .O(N__55757),
            .I(N__55742));
    Sp12to4 I__12427 (
            .O(N__55754),
            .I(N__55737));
    Span12Mux_v I__12426 (
            .O(N__55747),
            .I(N__55737));
    Odrv4 I__12425 (
            .O(N__55742),
            .I(\c0.n9_adj_3211 ));
    Odrv12 I__12424 (
            .O(N__55737),
            .I(\c0.n9_adj_3211 ));
    InMux I__12423 (
            .O(N__55732),
            .I(N__55729));
    LocalMux I__12422 (
            .O(N__55729),
            .I(N__55726));
    Span4Mux_h I__12421 (
            .O(N__55726),
            .I(N__55721));
    InMux I__12420 (
            .O(N__55725),
            .I(N__55718));
    InMux I__12419 (
            .O(N__55724),
            .I(N__55715));
    Odrv4 I__12418 (
            .O(N__55721),
            .I(\c0.n6_adj_3019 ));
    LocalMux I__12417 (
            .O(N__55718),
            .I(\c0.n6_adj_3019 ));
    LocalMux I__12416 (
            .O(N__55715),
            .I(\c0.n6_adj_3019 ));
    CascadeMux I__12415 (
            .O(N__55708),
            .I(N__55705));
    InMux I__12414 (
            .O(N__55705),
            .I(N__55701));
    InMux I__12413 (
            .O(N__55704),
            .I(N__55698));
    LocalMux I__12412 (
            .O(N__55701),
            .I(N__55693));
    LocalMux I__12411 (
            .O(N__55698),
            .I(N__55690));
    InMux I__12410 (
            .O(N__55697),
            .I(N__55685));
    InMux I__12409 (
            .O(N__55696),
            .I(N__55685));
    Odrv4 I__12408 (
            .O(N__55693),
            .I(\c0.data_in_frame_7_5 ));
    Odrv4 I__12407 (
            .O(N__55690),
            .I(\c0.data_in_frame_7_5 ));
    LocalMux I__12406 (
            .O(N__55685),
            .I(\c0.data_in_frame_7_5 ));
    CascadeMux I__12405 (
            .O(N__55678),
            .I(\c0.n6_adj_3019_cascade_ ));
    CascadeMux I__12404 (
            .O(N__55675),
            .I(N__55672));
    InMux I__12403 (
            .O(N__55672),
            .I(N__55665));
    CascadeMux I__12402 (
            .O(N__55671),
            .I(N__55662));
    InMux I__12401 (
            .O(N__55670),
            .I(N__55659));
    InMux I__12400 (
            .O(N__55669),
            .I(N__55656));
    InMux I__12399 (
            .O(N__55668),
            .I(N__55653));
    LocalMux I__12398 (
            .O(N__55665),
            .I(N__55650));
    InMux I__12397 (
            .O(N__55662),
            .I(N__55647));
    LocalMux I__12396 (
            .O(N__55659),
            .I(N__55642));
    LocalMux I__12395 (
            .O(N__55656),
            .I(N__55642));
    LocalMux I__12394 (
            .O(N__55653),
            .I(N__55639));
    Span4Mux_v I__12393 (
            .O(N__55650),
            .I(N__55636));
    LocalMux I__12392 (
            .O(N__55647),
            .I(N__55631));
    Span4Mux_v I__12391 (
            .O(N__55642),
            .I(N__55631));
    Span12Mux_h I__12390 (
            .O(N__55639),
            .I(N__55628));
    Span4Mux_v I__12389 (
            .O(N__55636),
            .I(N__55623));
    Span4Mux_h I__12388 (
            .O(N__55631),
            .I(N__55623));
    Odrv12 I__12387 (
            .O(N__55628),
            .I(\c0.n20386 ));
    Odrv4 I__12386 (
            .O(N__55623),
            .I(\c0.n20386 ));
    InMux I__12385 (
            .O(N__55618),
            .I(N__55615));
    LocalMux I__12384 (
            .O(N__55615),
            .I(N__55611));
    CascadeMux I__12383 (
            .O(N__55614),
            .I(N__55607));
    Span4Mux_h I__12382 (
            .O(N__55611),
            .I(N__55604));
    InMux I__12381 (
            .O(N__55610),
            .I(N__55601));
    InMux I__12380 (
            .O(N__55607),
            .I(N__55598));
    Span4Mux_v I__12379 (
            .O(N__55604),
            .I(N__55593));
    LocalMux I__12378 (
            .O(N__55601),
            .I(N__55593));
    LocalMux I__12377 (
            .O(N__55598),
            .I(\c0.data_in_frame_9_6 ));
    Odrv4 I__12376 (
            .O(N__55593),
            .I(\c0.data_in_frame_9_6 ));
    InMux I__12375 (
            .O(N__55588),
            .I(N__55580));
    InMux I__12374 (
            .O(N__55587),
            .I(N__55575));
    InMux I__12373 (
            .O(N__55586),
            .I(N__55575));
    InMux I__12372 (
            .O(N__55585),
            .I(N__55572));
    InMux I__12371 (
            .O(N__55584),
            .I(N__55569));
    InMux I__12370 (
            .O(N__55583),
            .I(N__55566));
    LocalMux I__12369 (
            .O(N__55580),
            .I(N__55559));
    LocalMux I__12368 (
            .O(N__55575),
            .I(N__55559));
    LocalMux I__12367 (
            .O(N__55572),
            .I(N__55559));
    LocalMux I__12366 (
            .O(N__55569),
            .I(N__55556));
    LocalMux I__12365 (
            .O(N__55566),
            .I(\c0.data_in_frame_3_7 ));
    Odrv12 I__12364 (
            .O(N__55559),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__12363 (
            .O(N__55556),
            .I(\c0.data_in_frame_3_7 ));
    InMux I__12362 (
            .O(N__55549),
            .I(N__55545));
    CascadeMux I__12361 (
            .O(N__55548),
            .I(N__55541));
    LocalMux I__12360 (
            .O(N__55545),
            .I(N__55537));
    InMux I__12359 (
            .O(N__55544),
            .I(N__55532));
    InMux I__12358 (
            .O(N__55541),
            .I(N__55532));
    InMux I__12357 (
            .O(N__55540),
            .I(N__55529));
    Span12Mux_h I__12356 (
            .O(N__55537),
            .I(N__55526));
    LocalMux I__12355 (
            .O(N__55532),
            .I(N__55523));
    LocalMux I__12354 (
            .O(N__55529),
            .I(\c0.data_in_frame_5_5 ));
    Odrv12 I__12353 (
            .O(N__55526),
            .I(\c0.data_in_frame_5_5 ));
    Odrv4 I__12352 (
            .O(N__55523),
            .I(\c0.data_in_frame_5_5 ));
    InMux I__12351 (
            .O(N__55516),
            .I(N__55512));
    CascadeMux I__12350 (
            .O(N__55515),
            .I(N__55506));
    LocalMux I__12349 (
            .O(N__55512),
            .I(N__55502));
    InMux I__12348 (
            .O(N__55511),
            .I(N__55499));
    InMux I__12347 (
            .O(N__55510),
            .I(N__55496));
    InMux I__12346 (
            .O(N__55509),
            .I(N__55493));
    InMux I__12345 (
            .O(N__55506),
            .I(N__55490));
    InMux I__12344 (
            .O(N__55505),
            .I(N__55487));
    Span4Mux_h I__12343 (
            .O(N__55502),
            .I(N__55484));
    LocalMux I__12342 (
            .O(N__55499),
            .I(N__55477));
    LocalMux I__12341 (
            .O(N__55496),
            .I(N__55477));
    LocalMux I__12340 (
            .O(N__55493),
            .I(N__55477));
    LocalMux I__12339 (
            .O(N__55490),
            .I(\c0.data_in_frame_5_3 ));
    LocalMux I__12338 (
            .O(N__55487),
            .I(\c0.data_in_frame_5_3 ));
    Odrv4 I__12337 (
            .O(N__55484),
            .I(\c0.data_in_frame_5_3 ));
    Odrv12 I__12336 (
            .O(N__55477),
            .I(\c0.data_in_frame_5_3 ));
    InMux I__12335 (
            .O(N__55468),
            .I(N__55462));
    InMux I__12334 (
            .O(N__55467),
            .I(N__55459));
    InMux I__12333 (
            .O(N__55466),
            .I(N__55454));
    InMux I__12332 (
            .O(N__55465),
            .I(N__55454));
    LocalMux I__12331 (
            .O(N__55462),
            .I(N__55451));
    LocalMux I__12330 (
            .O(N__55459),
            .I(N__55448));
    LocalMux I__12329 (
            .O(N__55454),
            .I(N__55445));
    Span4Mux_h I__12328 (
            .O(N__55451),
            .I(N__55442));
    Span4Mux_v I__12327 (
            .O(N__55448),
            .I(N__55439));
    Span4Mux_v I__12326 (
            .O(N__55445),
            .I(N__55436));
    Sp12to4 I__12325 (
            .O(N__55442),
            .I(N__55433));
    Span4Mux_v I__12324 (
            .O(N__55439),
            .I(N__55430));
    Sp12to4 I__12323 (
            .O(N__55436),
            .I(N__55425));
    Span12Mux_v I__12322 (
            .O(N__55433),
            .I(N__55425));
    Odrv4 I__12321 (
            .O(N__55430),
            .I(n11461));
    Odrv12 I__12320 (
            .O(N__55425),
            .I(n11461));
    InMux I__12319 (
            .O(N__55420),
            .I(N__55417));
    LocalMux I__12318 (
            .O(N__55417),
            .I(N__55414));
    Odrv4 I__12317 (
            .O(N__55414),
            .I(\c0.n11626 ));
    InMux I__12316 (
            .O(N__55411),
            .I(N__55408));
    LocalMux I__12315 (
            .O(N__55408),
            .I(N__55405));
    Odrv12 I__12314 (
            .O(N__55405),
            .I(\c0.n21_adj_3205 ));
    CascadeMux I__12313 (
            .O(N__55402),
            .I(N__55399));
    InMux I__12312 (
            .O(N__55399),
            .I(N__55396));
    LocalMux I__12311 (
            .O(N__55396),
            .I(N__55393));
    Span4Mux_v I__12310 (
            .O(N__55393),
            .I(N__55390));
    Span4Mux_h I__12309 (
            .O(N__55390),
            .I(N__55387));
    Odrv4 I__12308 (
            .O(N__55387),
            .I(\c0.n28_adj_3428 ));
    InMux I__12307 (
            .O(N__55384),
            .I(N__55379));
    InMux I__12306 (
            .O(N__55383),
            .I(N__55374));
    InMux I__12305 (
            .O(N__55382),
            .I(N__55371));
    LocalMux I__12304 (
            .O(N__55379),
            .I(N__55368));
    InMux I__12303 (
            .O(N__55378),
            .I(N__55365));
    InMux I__12302 (
            .O(N__55377),
            .I(N__55361));
    LocalMux I__12301 (
            .O(N__55374),
            .I(N__55358));
    LocalMux I__12300 (
            .O(N__55371),
            .I(N__55355));
    Span4Mux_h I__12299 (
            .O(N__55368),
            .I(N__55350));
    LocalMux I__12298 (
            .O(N__55365),
            .I(N__55350));
    InMux I__12297 (
            .O(N__55364),
            .I(N__55346));
    LocalMux I__12296 (
            .O(N__55361),
            .I(N__55341));
    Span4Mux_v I__12295 (
            .O(N__55358),
            .I(N__55338));
    Span4Mux_v I__12294 (
            .O(N__55355),
            .I(N__55333));
    Span4Mux_v I__12293 (
            .O(N__55350),
            .I(N__55333));
    InMux I__12292 (
            .O(N__55349),
            .I(N__55330));
    LocalMux I__12291 (
            .O(N__55346),
            .I(N__55327));
    InMux I__12290 (
            .O(N__55345),
            .I(N__55322));
    InMux I__12289 (
            .O(N__55344),
            .I(N__55322));
    Odrv4 I__12288 (
            .O(N__55341),
            .I(data_in_frame_1_5));
    Odrv4 I__12287 (
            .O(N__55338),
            .I(data_in_frame_1_5));
    Odrv4 I__12286 (
            .O(N__55333),
            .I(data_in_frame_1_5));
    LocalMux I__12285 (
            .O(N__55330),
            .I(data_in_frame_1_5));
    Odrv12 I__12284 (
            .O(N__55327),
            .I(data_in_frame_1_5));
    LocalMux I__12283 (
            .O(N__55322),
            .I(data_in_frame_1_5));
    CascadeMux I__12282 (
            .O(N__55309),
            .I(N__55305));
    InMux I__12281 (
            .O(N__55308),
            .I(N__55300));
    InMux I__12280 (
            .O(N__55305),
            .I(N__55300));
    LocalMux I__12279 (
            .O(N__55300),
            .I(N__55297));
    Odrv12 I__12278 (
            .O(N__55297),
            .I(\c0.n7_adj_3509 ));
    CascadeMux I__12277 (
            .O(N__55294),
            .I(\c0.n7_adj_3509_cascade_ ));
    CascadeMux I__12276 (
            .O(N__55291),
            .I(N__55288));
    InMux I__12275 (
            .O(N__55288),
            .I(N__55285));
    LocalMux I__12274 (
            .O(N__55285),
            .I(N__55281));
    InMux I__12273 (
            .O(N__55284),
            .I(N__55278));
    Span4Mux_v I__12272 (
            .O(N__55281),
            .I(N__55272));
    LocalMux I__12271 (
            .O(N__55278),
            .I(N__55272));
    InMux I__12270 (
            .O(N__55277),
            .I(N__55269));
    Odrv4 I__12269 (
            .O(N__55272),
            .I(\c0.n10_adj_3012 ));
    LocalMux I__12268 (
            .O(N__55269),
            .I(\c0.n10_adj_3012 ));
    InMux I__12267 (
            .O(N__55264),
            .I(N__55260));
    InMux I__12266 (
            .O(N__55263),
            .I(N__55257));
    LocalMux I__12265 (
            .O(N__55260),
            .I(N__55254));
    LocalMux I__12264 (
            .O(N__55257),
            .I(N__55251));
    Span4Mux_h I__12263 (
            .O(N__55254),
            .I(N__55248));
    Span4Mux_h I__12262 (
            .O(N__55251),
            .I(N__55245));
    Odrv4 I__12261 (
            .O(N__55248),
            .I(\c0.n45 ));
    Odrv4 I__12260 (
            .O(N__55245),
            .I(\c0.n45 ));
    InMux I__12259 (
            .O(N__55240),
            .I(N__55236));
    InMux I__12258 (
            .O(N__55239),
            .I(N__55231));
    LocalMux I__12257 (
            .O(N__55236),
            .I(N__55228));
    InMux I__12256 (
            .O(N__55235),
            .I(N__55225));
    CascadeMux I__12255 (
            .O(N__55234),
            .I(N__55222));
    LocalMux I__12254 (
            .O(N__55231),
            .I(N__55219));
    Span4Mux_v I__12253 (
            .O(N__55228),
            .I(N__55214));
    LocalMux I__12252 (
            .O(N__55225),
            .I(N__55214));
    InMux I__12251 (
            .O(N__55222),
            .I(N__55209));
    Span4Mux_v I__12250 (
            .O(N__55219),
            .I(N__55206));
    Span4Mux_h I__12249 (
            .O(N__55214),
            .I(N__55203));
    InMux I__12248 (
            .O(N__55213),
            .I(N__55200));
    InMux I__12247 (
            .O(N__55212),
            .I(N__55197));
    LocalMux I__12246 (
            .O(N__55209),
            .I(\c0.data_in_frame_4_1 ));
    Odrv4 I__12245 (
            .O(N__55206),
            .I(\c0.data_in_frame_4_1 ));
    Odrv4 I__12244 (
            .O(N__55203),
            .I(\c0.data_in_frame_4_1 ));
    LocalMux I__12243 (
            .O(N__55200),
            .I(\c0.data_in_frame_4_1 ));
    LocalMux I__12242 (
            .O(N__55197),
            .I(\c0.data_in_frame_4_1 ));
    CascadeMux I__12241 (
            .O(N__55186),
            .I(N__55175));
    InMux I__12240 (
            .O(N__55185),
            .I(N__55172));
    InMux I__12239 (
            .O(N__55184),
            .I(N__55169));
    InMux I__12238 (
            .O(N__55183),
            .I(N__55166));
    InMux I__12237 (
            .O(N__55182),
            .I(N__55157));
    InMux I__12236 (
            .O(N__55181),
            .I(N__55157));
    InMux I__12235 (
            .O(N__55180),
            .I(N__55154));
    InMux I__12234 (
            .O(N__55179),
            .I(N__55151));
    CascadeMux I__12233 (
            .O(N__55178),
            .I(N__55148));
    InMux I__12232 (
            .O(N__55175),
            .I(N__55144));
    LocalMux I__12231 (
            .O(N__55172),
            .I(N__55137));
    LocalMux I__12230 (
            .O(N__55169),
            .I(N__55137));
    LocalMux I__12229 (
            .O(N__55166),
            .I(N__55137));
    InMux I__12228 (
            .O(N__55165),
            .I(N__55130));
    InMux I__12227 (
            .O(N__55164),
            .I(N__55130));
    InMux I__12226 (
            .O(N__55163),
            .I(N__55130));
    CascadeMux I__12225 (
            .O(N__55162),
            .I(N__55124));
    LocalMux I__12224 (
            .O(N__55157),
            .I(N__55121));
    LocalMux I__12223 (
            .O(N__55154),
            .I(N__55118));
    LocalMux I__12222 (
            .O(N__55151),
            .I(N__55115));
    InMux I__12221 (
            .O(N__55148),
            .I(N__55110));
    InMux I__12220 (
            .O(N__55147),
            .I(N__55110));
    LocalMux I__12219 (
            .O(N__55144),
            .I(N__55105));
    Span4Mux_v I__12218 (
            .O(N__55137),
            .I(N__55100));
    LocalMux I__12217 (
            .O(N__55130),
            .I(N__55100));
    InMux I__12216 (
            .O(N__55129),
            .I(N__55095));
    InMux I__12215 (
            .O(N__55128),
            .I(N__55095));
    InMux I__12214 (
            .O(N__55127),
            .I(N__55092));
    InMux I__12213 (
            .O(N__55124),
            .I(N__55089));
    Span4Mux_v I__12212 (
            .O(N__55121),
            .I(N__55080));
    Span4Mux_v I__12211 (
            .O(N__55118),
            .I(N__55080));
    Span4Mux_h I__12210 (
            .O(N__55115),
            .I(N__55080));
    LocalMux I__12209 (
            .O(N__55110),
            .I(N__55080));
    InMux I__12208 (
            .O(N__55109),
            .I(N__55077));
    InMux I__12207 (
            .O(N__55108),
            .I(N__55074));
    Span4Mux_v I__12206 (
            .O(N__55105),
            .I(N__55069));
    Span4Mux_h I__12205 (
            .O(N__55100),
            .I(N__55069));
    LocalMux I__12204 (
            .O(N__55095),
            .I(data_in_frame_0_6));
    LocalMux I__12203 (
            .O(N__55092),
            .I(data_in_frame_0_6));
    LocalMux I__12202 (
            .O(N__55089),
            .I(data_in_frame_0_6));
    Odrv4 I__12201 (
            .O(N__55080),
            .I(data_in_frame_0_6));
    LocalMux I__12200 (
            .O(N__55077),
            .I(data_in_frame_0_6));
    LocalMux I__12199 (
            .O(N__55074),
            .I(data_in_frame_0_6));
    Odrv4 I__12198 (
            .O(N__55069),
            .I(data_in_frame_0_6));
    InMux I__12197 (
            .O(N__55054),
            .I(N__55049));
    InMux I__12196 (
            .O(N__55053),
            .I(N__55046));
    InMux I__12195 (
            .O(N__55052),
            .I(N__55043));
    LocalMux I__12194 (
            .O(N__55049),
            .I(N__55040));
    LocalMux I__12193 (
            .O(N__55046),
            .I(N__55035));
    LocalMux I__12192 (
            .O(N__55043),
            .I(N__55035));
    Span4Mux_h I__12191 (
            .O(N__55040),
            .I(N__55028));
    Span4Mux_h I__12190 (
            .O(N__55035),
            .I(N__55025));
    InMux I__12189 (
            .O(N__55034),
            .I(N__55022));
    InMux I__12188 (
            .O(N__55033),
            .I(N__55017));
    InMux I__12187 (
            .O(N__55032),
            .I(N__55017));
    CascadeMux I__12186 (
            .O(N__55031),
            .I(N__55011));
    Span4Mux_h I__12185 (
            .O(N__55028),
            .I(N__55007));
    Span4Mux_v I__12184 (
            .O(N__55025),
            .I(N__55000));
    LocalMux I__12183 (
            .O(N__55022),
            .I(N__55000));
    LocalMux I__12182 (
            .O(N__55017),
            .I(N__55000));
    InMux I__12181 (
            .O(N__55016),
            .I(N__54995));
    InMux I__12180 (
            .O(N__55015),
            .I(N__54995));
    InMux I__12179 (
            .O(N__55014),
            .I(N__54992));
    InMux I__12178 (
            .O(N__55011),
            .I(N__54987));
    InMux I__12177 (
            .O(N__55010),
            .I(N__54987));
    Odrv4 I__12176 (
            .O(N__55007),
            .I(data_in_frame_1_0));
    Odrv4 I__12175 (
            .O(N__55000),
            .I(data_in_frame_1_0));
    LocalMux I__12174 (
            .O(N__54995),
            .I(data_in_frame_1_0));
    LocalMux I__12173 (
            .O(N__54992),
            .I(data_in_frame_1_0));
    LocalMux I__12172 (
            .O(N__54987),
            .I(data_in_frame_1_0));
    InMux I__12171 (
            .O(N__54976),
            .I(N__54973));
    LocalMux I__12170 (
            .O(N__54973),
            .I(N__54970));
    Span4Mux_v I__12169 (
            .O(N__54970),
            .I(N__54967));
    Span4Mux_h I__12168 (
            .O(N__54967),
            .I(N__54962));
    InMux I__12167 (
            .O(N__54966),
            .I(N__54957));
    InMux I__12166 (
            .O(N__54965),
            .I(N__54957));
    Odrv4 I__12165 (
            .O(N__54962),
            .I(\c0.n20341 ));
    LocalMux I__12164 (
            .O(N__54957),
            .I(\c0.n20341 ));
    InMux I__12163 (
            .O(N__54952),
            .I(N__54949));
    LocalMux I__12162 (
            .O(N__54949),
            .I(N__54946));
    Odrv4 I__12161 (
            .O(N__54946),
            .I(\c0.n58_adj_3497 ));
    InMux I__12160 (
            .O(N__54943),
            .I(N__54940));
    LocalMux I__12159 (
            .O(N__54940),
            .I(\c0.n56_adj_3505 ));
    InMux I__12158 (
            .O(N__54937),
            .I(N__54934));
    LocalMux I__12157 (
            .O(N__54934),
            .I(N__54931));
    Span4Mux_h I__12156 (
            .O(N__54931),
            .I(N__54928));
    Odrv4 I__12155 (
            .O(N__54928),
            .I(\c0.n64_adj_3506 ));
    InMux I__12154 (
            .O(N__54925),
            .I(N__54922));
    LocalMux I__12153 (
            .O(N__54922),
            .I(N__54919));
    Span12Mux_s10_h I__12152 (
            .O(N__54919),
            .I(N__54916));
    Odrv12 I__12151 (
            .O(N__54916),
            .I(\c0.n19217 ));
    CascadeMux I__12150 (
            .O(N__54913),
            .I(\c0.n4_adj_3036_cascade_ ));
    InMux I__12149 (
            .O(N__54910),
            .I(N__54907));
    LocalMux I__12148 (
            .O(N__54907),
            .I(\c0.n57_adj_3499 ));
    CascadeMux I__12147 (
            .O(N__54904),
            .I(\c0.n11478_cascade_ ));
    InMux I__12146 (
            .O(N__54901),
            .I(N__54898));
    LocalMux I__12145 (
            .O(N__54898),
            .I(\c0.n81 ));
    InMux I__12144 (
            .O(N__54895),
            .I(N__54889));
    CascadeMux I__12143 (
            .O(N__54894),
            .I(N__54884));
    InMux I__12142 (
            .O(N__54893),
            .I(N__54881));
    InMux I__12141 (
            .O(N__54892),
            .I(N__54877));
    LocalMux I__12140 (
            .O(N__54889),
            .I(N__54873));
    InMux I__12139 (
            .O(N__54888),
            .I(N__54868));
    InMux I__12138 (
            .O(N__54887),
            .I(N__54868));
    InMux I__12137 (
            .O(N__54884),
            .I(N__54865));
    LocalMux I__12136 (
            .O(N__54881),
            .I(N__54862));
    InMux I__12135 (
            .O(N__54880),
            .I(N__54859));
    LocalMux I__12134 (
            .O(N__54877),
            .I(N__54855));
    InMux I__12133 (
            .O(N__54876),
            .I(N__54852));
    Span4Mux_h I__12132 (
            .O(N__54873),
            .I(N__54846));
    LocalMux I__12131 (
            .O(N__54868),
            .I(N__54846));
    LocalMux I__12130 (
            .O(N__54865),
            .I(N__54843));
    Span4Mux_h I__12129 (
            .O(N__54862),
            .I(N__54837));
    LocalMux I__12128 (
            .O(N__54859),
            .I(N__54837));
    CascadeMux I__12127 (
            .O(N__54858),
            .I(N__54831));
    Span12Mux_h I__12126 (
            .O(N__54855),
            .I(N__54828));
    LocalMux I__12125 (
            .O(N__54852),
            .I(N__54825));
    InMux I__12124 (
            .O(N__54851),
            .I(N__54822));
    Span4Mux_v I__12123 (
            .O(N__54846),
            .I(N__54819));
    Span4Mux_h I__12122 (
            .O(N__54843),
            .I(N__54816));
    InMux I__12121 (
            .O(N__54842),
            .I(N__54813));
    Span4Mux_h I__12120 (
            .O(N__54837),
            .I(N__54810));
    InMux I__12119 (
            .O(N__54836),
            .I(N__54807));
    InMux I__12118 (
            .O(N__54835),
            .I(N__54800));
    InMux I__12117 (
            .O(N__54834),
            .I(N__54800));
    InMux I__12116 (
            .O(N__54831),
            .I(N__54800));
    Odrv12 I__12115 (
            .O(N__54828),
            .I(data_in_frame_1_6));
    Odrv12 I__12114 (
            .O(N__54825),
            .I(data_in_frame_1_6));
    LocalMux I__12113 (
            .O(N__54822),
            .I(data_in_frame_1_6));
    Odrv4 I__12112 (
            .O(N__54819),
            .I(data_in_frame_1_6));
    Odrv4 I__12111 (
            .O(N__54816),
            .I(data_in_frame_1_6));
    LocalMux I__12110 (
            .O(N__54813),
            .I(data_in_frame_1_6));
    Odrv4 I__12109 (
            .O(N__54810),
            .I(data_in_frame_1_6));
    LocalMux I__12108 (
            .O(N__54807),
            .I(data_in_frame_1_6));
    LocalMux I__12107 (
            .O(N__54800),
            .I(data_in_frame_1_6));
    InMux I__12106 (
            .O(N__54781),
            .I(N__54778));
    LocalMux I__12105 (
            .O(N__54778),
            .I(\c0.n11526 ));
    CascadeMux I__12104 (
            .O(N__54775),
            .I(N__54772));
    InMux I__12103 (
            .O(N__54772),
            .I(N__54767));
    InMux I__12102 (
            .O(N__54771),
            .I(N__54762));
    InMux I__12101 (
            .O(N__54770),
            .I(N__54762));
    LocalMux I__12100 (
            .O(N__54767),
            .I(\c0.data_in_frame_6_5 ));
    LocalMux I__12099 (
            .O(N__54762),
            .I(\c0.data_in_frame_6_5 ));
    CascadeMux I__12098 (
            .O(N__54757),
            .I(N__54754));
    InMux I__12097 (
            .O(N__54754),
            .I(N__54751));
    LocalMux I__12096 (
            .O(N__54751),
            .I(N__54747));
    InMux I__12095 (
            .O(N__54750),
            .I(N__54744));
    Span4Mux_h I__12094 (
            .O(N__54747),
            .I(N__54741));
    LocalMux I__12093 (
            .O(N__54744),
            .I(N__54738));
    Odrv4 I__12092 (
            .O(N__54741),
            .I(\c0.n11549 ));
    Odrv4 I__12091 (
            .O(N__54738),
            .I(\c0.n11549 ));
    InMux I__12090 (
            .O(N__54733),
            .I(N__54728));
    InMux I__12089 (
            .O(N__54732),
            .I(N__54722));
    InMux I__12088 (
            .O(N__54731),
            .I(N__54722));
    LocalMux I__12087 (
            .O(N__54728),
            .I(N__54719));
    InMux I__12086 (
            .O(N__54727),
            .I(N__54716));
    LocalMux I__12085 (
            .O(N__54722),
            .I(N__54713));
    Odrv12 I__12084 (
            .O(N__54719),
            .I(\c0.n11651 ));
    LocalMux I__12083 (
            .O(N__54716),
            .I(\c0.n11651 ));
    Odrv4 I__12082 (
            .O(N__54713),
            .I(\c0.n11651 ));
    InMux I__12081 (
            .O(N__54706),
            .I(N__54703));
    LocalMux I__12080 (
            .O(N__54703),
            .I(N__54700));
    Span4Mux_h I__12079 (
            .O(N__54700),
            .I(N__54697));
    Span4Mux_h I__12078 (
            .O(N__54697),
            .I(N__54694));
    Odrv4 I__12077 (
            .O(N__54694),
            .I(\c0.n27_adj_3457 ));
    InMux I__12076 (
            .O(N__54691),
            .I(N__54688));
    LocalMux I__12075 (
            .O(N__54688),
            .I(N__54685));
    Span4Mux_h I__12074 (
            .O(N__54685),
            .I(N__54681));
    CascadeMux I__12073 (
            .O(N__54684),
            .I(N__54677));
    Span4Mux_v I__12072 (
            .O(N__54681),
            .I(N__54668));
    InMux I__12071 (
            .O(N__54680),
            .I(N__54665));
    InMux I__12070 (
            .O(N__54677),
            .I(N__54658));
    InMux I__12069 (
            .O(N__54676),
            .I(N__54658));
    InMux I__12068 (
            .O(N__54675),
            .I(N__54658));
    InMux I__12067 (
            .O(N__54674),
            .I(N__54655));
    InMux I__12066 (
            .O(N__54673),
            .I(N__54652));
    InMux I__12065 (
            .O(N__54672),
            .I(N__54647));
    InMux I__12064 (
            .O(N__54671),
            .I(N__54647));
    Odrv4 I__12063 (
            .O(N__54668),
            .I(data_in_frame_1_7));
    LocalMux I__12062 (
            .O(N__54665),
            .I(data_in_frame_1_7));
    LocalMux I__12061 (
            .O(N__54658),
            .I(data_in_frame_1_7));
    LocalMux I__12060 (
            .O(N__54655),
            .I(data_in_frame_1_7));
    LocalMux I__12059 (
            .O(N__54652),
            .I(data_in_frame_1_7));
    LocalMux I__12058 (
            .O(N__54647),
            .I(data_in_frame_1_7));
    InMux I__12057 (
            .O(N__54634),
            .I(N__54631));
    LocalMux I__12056 (
            .O(N__54631),
            .I(\c0.n12_adj_3378 ));
    CascadeMux I__12055 (
            .O(N__54628),
            .I(N__54624));
    CascadeMux I__12054 (
            .O(N__54627),
            .I(N__54620));
    InMux I__12053 (
            .O(N__54624),
            .I(N__54617));
    InMux I__12052 (
            .O(N__54623),
            .I(N__54614));
    InMux I__12051 (
            .O(N__54620),
            .I(N__54609));
    LocalMux I__12050 (
            .O(N__54617),
            .I(N__54606));
    LocalMux I__12049 (
            .O(N__54614),
            .I(N__54603));
    InMux I__12048 (
            .O(N__54613),
            .I(N__54598));
    InMux I__12047 (
            .O(N__54612),
            .I(N__54598));
    LocalMux I__12046 (
            .O(N__54609),
            .I(\c0.data_in_frame_2_1 ));
    Odrv12 I__12045 (
            .O(N__54606),
            .I(\c0.data_in_frame_2_1 ));
    Odrv12 I__12044 (
            .O(N__54603),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__12043 (
            .O(N__54598),
            .I(\c0.data_in_frame_2_1 ));
    InMux I__12042 (
            .O(N__54589),
            .I(N__54586));
    LocalMux I__12041 (
            .O(N__54586),
            .I(N__54583));
    Odrv12 I__12040 (
            .O(N__54583),
            .I(\c0.n34_adj_3326 ));
    CascadeMux I__12039 (
            .O(N__54580),
            .I(N__54576));
    InMux I__12038 (
            .O(N__54579),
            .I(N__54571));
    InMux I__12037 (
            .O(N__54576),
            .I(N__54571));
    LocalMux I__12036 (
            .O(N__54571),
            .I(\c0.n13_adj_3344 ));
    InMux I__12035 (
            .O(N__54568),
            .I(N__54564));
    CascadeMux I__12034 (
            .O(N__54567),
            .I(N__54561));
    LocalMux I__12033 (
            .O(N__54564),
            .I(N__54557));
    InMux I__12032 (
            .O(N__54561),
            .I(N__54553));
    InMux I__12031 (
            .O(N__54560),
            .I(N__54550));
    Span12Mux_h I__12030 (
            .O(N__54557),
            .I(N__54547));
    InMux I__12029 (
            .O(N__54556),
            .I(N__54544));
    LocalMux I__12028 (
            .O(N__54553),
            .I(N__54541));
    LocalMux I__12027 (
            .O(N__54550),
            .I(\c0.n23_adj_3076 ));
    Odrv12 I__12026 (
            .O(N__54547),
            .I(\c0.n23_adj_3076 ));
    LocalMux I__12025 (
            .O(N__54544),
            .I(\c0.n23_adj_3076 ));
    Odrv4 I__12024 (
            .O(N__54541),
            .I(\c0.n23_adj_3076 ));
    InMux I__12023 (
            .O(N__54532),
            .I(N__54525));
    InMux I__12022 (
            .O(N__54531),
            .I(N__54525));
    InMux I__12021 (
            .O(N__54530),
            .I(N__54522));
    LocalMux I__12020 (
            .O(N__54525),
            .I(N__54519));
    LocalMux I__12019 (
            .O(N__54522),
            .I(N__54515));
    Span4Mux_v I__12018 (
            .O(N__54519),
            .I(N__54512));
    InMux I__12017 (
            .O(N__54518),
            .I(N__54509));
    Odrv4 I__12016 (
            .O(N__54515),
            .I(\c0.n19424 ));
    Odrv4 I__12015 (
            .O(N__54512),
            .I(\c0.n19424 ));
    LocalMux I__12014 (
            .O(N__54509),
            .I(\c0.n19424 ));
    CascadeMux I__12013 (
            .O(N__54502),
            .I(N__54499));
    InMux I__12012 (
            .O(N__54499),
            .I(N__54496));
    LocalMux I__12011 (
            .O(N__54496),
            .I(N__54493));
    Span4Mux_v I__12010 (
            .O(N__54493),
            .I(N__54489));
    InMux I__12009 (
            .O(N__54492),
            .I(N__54486));
    Odrv4 I__12008 (
            .O(N__54489),
            .I(\c0.n7_adj_3029 ));
    LocalMux I__12007 (
            .O(N__54486),
            .I(\c0.n7_adj_3029 ));
    CascadeMux I__12006 (
            .O(N__54481),
            .I(N__54476));
    InMux I__12005 (
            .O(N__54480),
            .I(N__54473));
    CascadeMux I__12004 (
            .O(N__54479),
            .I(N__54469));
    InMux I__12003 (
            .O(N__54476),
            .I(N__54463));
    LocalMux I__12002 (
            .O(N__54473),
            .I(N__54456));
    CascadeMux I__12001 (
            .O(N__54472),
            .I(N__54453));
    InMux I__12000 (
            .O(N__54469),
            .I(N__54449));
    InMux I__11999 (
            .O(N__54468),
            .I(N__54446));
    InMux I__11998 (
            .O(N__54467),
            .I(N__54443));
    InMux I__11997 (
            .O(N__54466),
            .I(N__54439));
    LocalMux I__11996 (
            .O(N__54463),
            .I(N__54436));
    InMux I__11995 (
            .O(N__54462),
            .I(N__54431));
    InMux I__11994 (
            .O(N__54461),
            .I(N__54431));
    InMux I__11993 (
            .O(N__54460),
            .I(N__54428));
    CascadeMux I__11992 (
            .O(N__54459),
            .I(N__54424));
    Span4Mux_v I__11991 (
            .O(N__54456),
            .I(N__54418));
    InMux I__11990 (
            .O(N__54453),
            .I(N__54415));
    InMux I__11989 (
            .O(N__54452),
            .I(N__54412));
    LocalMux I__11988 (
            .O(N__54449),
            .I(N__54405));
    LocalMux I__11987 (
            .O(N__54446),
            .I(N__54405));
    LocalMux I__11986 (
            .O(N__54443),
            .I(N__54402));
    InMux I__11985 (
            .O(N__54442),
            .I(N__54399));
    LocalMux I__11984 (
            .O(N__54439),
            .I(N__54396));
    Span4Mux_h I__11983 (
            .O(N__54436),
            .I(N__54388));
    LocalMux I__11982 (
            .O(N__54431),
            .I(N__54388));
    LocalMux I__11981 (
            .O(N__54428),
            .I(N__54388));
    InMux I__11980 (
            .O(N__54427),
            .I(N__54385));
    InMux I__11979 (
            .O(N__54424),
            .I(N__54378));
    InMux I__11978 (
            .O(N__54423),
            .I(N__54378));
    InMux I__11977 (
            .O(N__54422),
            .I(N__54373));
    InMux I__11976 (
            .O(N__54421),
            .I(N__54373));
    Span4Mux_h I__11975 (
            .O(N__54418),
            .I(N__54370));
    LocalMux I__11974 (
            .O(N__54415),
            .I(N__54365));
    LocalMux I__11973 (
            .O(N__54412),
            .I(N__54365));
    InMux I__11972 (
            .O(N__54411),
            .I(N__54360));
    InMux I__11971 (
            .O(N__54410),
            .I(N__54360));
    Span4Mux_h I__11970 (
            .O(N__54405),
            .I(N__54351));
    Span4Mux_v I__11969 (
            .O(N__54402),
            .I(N__54351));
    LocalMux I__11968 (
            .O(N__54399),
            .I(N__54351));
    Span4Mux_h I__11967 (
            .O(N__54396),
            .I(N__54351));
    InMux I__11966 (
            .O(N__54395),
            .I(N__54348));
    Span4Mux_h I__11965 (
            .O(N__54388),
            .I(N__54343));
    LocalMux I__11964 (
            .O(N__54385),
            .I(N__54343));
    InMux I__11963 (
            .O(N__54384),
            .I(N__54340));
    InMux I__11962 (
            .O(N__54383),
            .I(N__54337));
    LocalMux I__11961 (
            .O(N__54378),
            .I(data_in_frame_0_4));
    LocalMux I__11960 (
            .O(N__54373),
            .I(data_in_frame_0_4));
    Odrv4 I__11959 (
            .O(N__54370),
            .I(data_in_frame_0_4));
    Odrv12 I__11958 (
            .O(N__54365),
            .I(data_in_frame_0_4));
    LocalMux I__11957 (
            .O(N__54360),
            .I(data_in_frame_0_4));
    Odrv4 I__11956 (
            .O(N__54351),
            .I(data_in_frame_0_4));
    LocalMux I__11955 (
            .O(N__54348),
            .I(data_in_frame_0_4));
    Odrv4 I__11954 (
            .O(N__54343),
            .I(data_in_frame_0_4));
    LocalMux I__11953 (
            .O(N__54340),
            .I(data_in_frame_0_4));
    LocalMux I__11952 (
            .O(N__54337),
            .I(data_in_frame_0_4));
    CascadeMux I__11951 (
            .O(N__54316),
            .I(N__54312));
    InMux I__11950 (
            .O(N__54315),
            .I(N__54309));
    InMux I__11949 (
            .O(N__54312),
            .I(N__54305));
    LocalMux I__11948 (
            .O(N__54309),
            .I(N__54302));
    InMux I__11947 (
            .O(N__54308),
            .I(N__54299));
    LocalMux I__11946 (
            .O(N__54305),
            .I(N__54291));
    Span4Mux_h I__11945 (
            .O(N__54302),
            .I(N__54291));
    LocalMux I__11944 (
            .O(N__54299),
            .I(N__54288));
    InMux I__11943 (
            .O(N__54298),
            .I(N__54285));
    InMux I__11942 (
            .O(N__54297),
            .I(N__54280));
    InMux I__11941 (
            .O(N__54296),
            .I(N__54280));
    Odrv4 I__11940 (
            .O(N__54291),
            .I(\c0.data_in_frame_2_3 ));
    Odrv12 I__11939 (
            .O(N__54288),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__11938 (
            .O(N__54285),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__11937 (
            .O(N__54280),
            .I(\c0.data_in_frame_2_3 ));
    InMux I__11936 (
            .O(N__54271),
            .I(N__54268));
    LocalMux I__11935 (
            .O(N__54268),
            .I(N__54263));
    InMux I__11934 (
            .O(N__54267),
            .I(N__54258));
    CascadeMux I__11933 (
            .O(N__54266),
            .I(N__54255));
    Span4Mux_v I__11932 (
            .O(N__54263),
            .I(N__54251));
    InMux I__11931 (
            .O(N__54262),
            .I(N__54246));
    InMux I__11930 (
            .O(N__54261),
            .I(N__54246));
    LocalMux I__11929 (
            .O(N__54258),
            .I(N__54243));
    InMux I__11928 (
            .O(N__54255),
            .I(N__54239));
    InMux I__11927 (
            .O(N__54254),
            .I(N__54236));
    Span4Mux_h I__11926 (
            .O(N__54251),
            .I(N__54233));
    LocalMux I__11925 (
            .O(N__54246),
            .I(N__54230));
    Span4Mux_h I__11924 (
            .O(N__54243),
            .I(N__54227));
    InMux I__11923 (
            .O(N__54242),
            .I(N__54224));
    LocalMux I__11922 (
            .O(N__54239),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__11921 (
            .O(N__54236),
            .I(\c0.data_in_frame_4_4 ));
    Odrv4 I__11920 (
            .O(N__54233),
            .I(\c0.data_in_frame_4_4 ));
    Odrv4 I__11919 (
            .O(N__54230),
            .I(\c0.data_in_frame_4_4 ));
    Odrv4 I__11918 (
            .O(N__54227),
            .I(\c0.data_in_frame_4_4 ));
    LocalMux I__11917 (
            .O(N__54224),
            .I(\c0.data_in_frame_4_4 ));
    InMux I__11916 (
            .O(N__54211),
            .I(N__54205));
    InMux I__11915 (
            .O(N__54210),
            .I(N__54205));
    LocalMux I__11914 (
            .O(N__54205),
            .I(N__54202));
    Odrv4 I__11913 (
            .O(N__54202),
            .I(\c0.n8_adj_3345 ));
    InMux I__11912 (
            .O(N__54199),
            .I(N__54195));
    InMux I__11911 (
            .O(N__54198),
            .I(N__54192));
    LocalMux I__11910 (
            .O(N__54195),
            .I(\c0.n7_adj_3520 ));
    LocalMux I__11909 (
            .O(N__54192),
            .I(\c0.n7_adj_3520 ));
    InMux I__11908 (
            .O(N__54187),
            .I(N__54178));
    InMux I__11907 (
            .O(N__54186),
            .I(N__54178));
    InMux I__11906 (
            .O(N__54185),
            .I(N__54178));
    LocalMux I__11905 (
            .O(N__54178),
            .I(N__54175));
    Odrv4 I__11904 (
            .O(N__54175),
            .I(\c0.n9_adj_3346 ));
    CascadeMux I__11903 (
            .O(N__54172),
            .I(\c0.n8_adj_3345_cascade_ ));
    CascadeMux I__11902 (
            .O(N__54169),
            .I(\c0.n11626_cascade_ ));
    InMux I__11901 (
            .O(N__54166),
            .I(N__54163));
    LocalMux I__11900 (
            .O(N__54163),
            .I(N__54159));
    CascadeMux I__11899 (
            .O(N__54162),
            .I(N__54156));
    Span4Mux_h I__11898 (
            .O(N__54159),
            .I(N__54152));
    InMux I__11897 (
            .O(N__54156),
            .I(N__54149));
    InMux I__11896 (
            .O(N__54155),
            .I(N__54146));
    Span4Mux_v I__11895 (
            .O(N__54152),
            .I(N__54143));
    LocalMux I__11894 (
            .O(N__54149),
            .I(\c0.data_in_frame_8_7 ));
    LocalMux I__11893 (
            .O(N__54146),
            .I(\c0.data_in_frame_8_7 ));
    Odrv4 I__11892 (
            .O(N__54143),
            .I(\c0.data_in_frame_8_7 ));
    InMux I__11891 (
            .O(N__54136),
            .I(N__54131));
    InMux I__11890 (
            .O(N__54135),
            .I(N__54127));
    InMux I__11889 (
            .O(N__54134),
            .I(N__54123));
    LocalMux I__11888 (
            .O(N__54131),
            .I(N__54119));
    InMux I__11887 (
            .O(N__54130),
            .I(N__54116));
    LocalMux I__11886 (
            .O(N__54127),
            .I(N__54112));
    InMux I__11885 (
            .O(N__54126),
            .I(N__54109));
    LocalMux I__11884 (
            .O(N__54123),
            .I(N__54106));
    InMux I__11883 (
            .O(N__54122),
            .I(N__54103));
    Span4Mux_v I__11882 (
            .O(N__54119),
            .I(N__54098));
    LocalMux I__11881 (
            .O(N__54116),
            .I(N__54098));
    InMux I__11880 (
            .O(N__54115),
            .I(N__54091));
    Span4Mux_h I__11879 (
            .O(N__54112),
            .I(N__54088));
    LocalMux I__11878 (
            .O(N__54109),
            .I(N__54079));
    Span4Mux_h I__11877 (
            .O(N__54106),
            .I(N__54079));
    LocalMux I__11876 (
            .O(N__54103),
            .I(N__54079));
    Span4Mux_v I__11875 (
            .O(N__54098),
            .I(N__54079));
    InMux I__11874 (
            .O(N__54097),
            .I(N__54070));
    InMux I__11873 (
            .O(N__54096),
            .I(N__54070));
    InMux I__11872 (
            .O(N__54095),
            .I(N__54070));
    InMux I__11871 (
            .O(N__54094),
            .I(N__54070));
    LocalMux I__11870 (
            .O(N__54091),
            .I(N__54067));
    Odrv4 I__11869 (
            .O(N__54088),
            .I(data_in_frame_1_1));
    Odrv4 I__11868 (
            .O(N__54079),
            .I(data_in_frame_1_1));
    LocalMux I__11867 (
            .O(N__54070),
            .I(data_in_frame_1_1));
    Odrv4 I__11866 (
            .O(N__54067),
            .I(data_in_frame_1_1));
    InMux I__11865 (
            .O(N__54058),
            .I(N__54055));
    LocalMux I__11864 (
            .O(N__54055),
            .I(N__54051));
    InMux I__11863 (
            .O(N__54054),
            .I(N__54048));
    Span4Mux_v I__11862 (
            .O(N__54051),
            .I(N__54045));
    LocalMux I__11861 (
            .O(N__54048),
            .I(N__54042));
    Span4Mux_h I__11860 (
            .O(N__54045),
            .I(N__54039));
    Span4Mux_v I__11859 (
            .O(N__54042),
            .I(N__54036));
    Odrv4 I__11858 (
            .O(N__54039),
            .I(\c0.n19970 ));
    Odrv4 I__11857 (
            .O(N__54036),
            .I(\c0.n19970 ));
    InMux I__11856 (
            .O(N__54031),
            .I(N__54028));
    LocalMux I__11855 (
            .O(N__54028),
            .I(N__54025));
    Odrv12 I__11854 (
            .O(N__54025),
            .I(\c0.n6_adj_3501 ));
    CascadeMux I__11853 (
            .O(N__54022),
            .I(N__54017));
    InMux I__11852 (
            .O(N__54021),
            .I(N__54014));
    CascadeMux I__11851 (
            .O(N__54020),
            .I(N__54011));
    InMux I__11850 (
            .O(N__54017),
            .I(N__54008));
    LocalMux I__11849 (
            .O(N__54014),
            .I(N__54005));
    InMux I__11848 (
            .O(N__54011),
            .I(N__54002));
    LocalMux I__11847 (
            .O(N__54008),
            .I(N__53999));
    Span4Mux_v I__11846 (
            .O(N__54005),
            .I(N__53996));
    LocalMux I__11845 (
            .O(N__54002),
            .I(N__53993));
    Odrv12 I__11844 (
            .O(N__53999),
            .I(\c0.data_in_frame_6_3 ));
    Odrv4 I__11843 (
            .O(N__53996),
            .I(\c0.data_in_frame_6_3 ));
    Odrv4 I__11842 (
            .O(N__53993),
            .I(\c0.data_in_frame_6_3 ));
    InMux I__11841 (
            .O(N__53986),
            .I(N__53983));
    LocalMux I__11840 (
            .O(N__53983),
            .I(N__53980));
    Span4Mux_v I__11839 (
            .O(N__53980),
            .I(N__53977));
    Odrv4 I__11838 (
            .O(N__53977),
            .I(\c0.n25_adj_3048 ));
    InMux I__11837 (
            .O(N__53974),
            .I(N__53970));
    InMux I__11836 (
            .O(N__53973),
            .I(N__53967));
    LocalMux I__11835 (
            .O(N__53970),
            .I(N__53964));
    LocalMux I__11834 (
            .O(N__53967),
            .I(N__53960));
    Span4Mux_v I__11833 (
            .O(N__53964),
            .I(N__53957));
    InMux I__11832 (
            .O(N__53963),
            .I(N__53954));
    Odrv4 I__11831 (
            .O(N__53960),
            .I(\c0.n19312 ));
    Odrv4 I__11830 (
            .O(N__53957),
            .I(\c0.n19312 ));
    LocalMux I__11829 (
            .O(N__53954),
            .I(\c0.n19312 ));
    InMux I__11828 (
            .O(N__53947),
            .I(N__53944));
    LocalMux I__11827 (
            .O(N__53944),
            .I(N__53939));
    InMux I__11826 (
            .O(N__53943),
            .I(N__53936));
    InMux I__11825 (
            .O(N__53942),
            .I(N__53933));
    Span4Mux_h I__11824 (
            .O(N__53939),
            .I(N__53930));
    LocalMux I__11823 (
            .O(N__53936),
            .I(N__53927));
    LocalMux I__11822 (
            .O(N__53933),
            .I(N__53924));
    Span4Mux_v I__11821 (
            .O(N__53930),
            .I(N__53921));
    Span4Mux_h I__11820 (
            .O(N__53927),
            .I(N__53918));
    Odrv12 I__11819 (
            .O(N__53924),
            .I(\c0.n20512 ));
    Odrv4 I__11818 (
            .O(N__53921),
            .I(\c0.n20512 ));
    Odrv4 I__11817 (
            .O(N__53918),
            .I(\c0.n20512 ));
    InMux I__11816 (
            .O(N__53911),
            .I(N__53908));
    LocalMux I__11815 (
            .O(N__53908),
            .I(N__53904));
    InMux I__11814 (
            .O(N__53907),
            .I(N__53901));
    Span4Mux_v I__11813 (
            .O(N__53904),
            .I(N__53898));
    LocalMux I__11812 (
            .O(N__53901),
            .I(N__53895));
    Span4Mux_v I__11811 (
            .O(N__53898),
            .I(N__53892));
    Span4Mux_v I__11810 (
            .O(N__53895),
            .I(N__53889));
    Odrv4 I__11809 (
            .O(N__53892),
            .I(\c0.n19202 ));
    Odrv4 I__11808 (
            .O(N__53889),
            .I(\c0.n19202 ));
    CascadeMux I__11807 (
            .O(N__53884),
            .I(\c0.n12_adj_3210_cascade_ ));
    InMux I__11806 (
            .O(N__53881),
            .I(N__53878));
    LocalMux I__11805 (
            .O(N__53878),
            .I(N__53875));
    Span4Mux_h I__11804 (
            .O(N__53875),
            .I(N__53871));
    InMux I__11803 (
            .O(N__53874),
            .I(N__53865));
    Span4Mux_v I__11802 (
            .O(N__53871),
            .I(N__53862));
    InMux I__11801 (
            .O(N__53870),
            .I(N__53859));
    InMux I__11800 (
            .O(N__53869),
            .I(N__53854));
    InMux I__11799 (
            .O(N__53868),
            .I(N__53854));
    LocalMux I__11798 (
            .O(N__53865),
            .I(N__53851));
    Odrv4 I__11797 (
            .O(N__53862),
            .I(\c0.n18433 ));
    LocalMux I__11796 (
            .O(N__53859),
            .I(\c0.n18433 ));
    LocalMux I__11795 (
            .O(N__53854),
            .I(\c0.n18433 ));
    Odrv4 I__11794 (
            .O(N__53851),
            .I(\c0.n18433 ));
    InMux I__11793 (
            .O(N__53842),
            .I(N__53839));
    LocalMux I__11792 (
            .O(N__53839),
            .I(N__53834));
    InMux I__11791 (
            .O(N__53838),
            .I(N__53829));
    InMux I__11790 (
            .O(N__53837),
            .I(N__53829));
    Odrv4 I__11789 (
            .O(N__53834),
            .I(\c0.n17834 ));
    LocalMux I__11788 (
            .O(N__53829),
            .I(\c0.n17834 ));
    CascadeMux I__11787 (
            .O(N__53824),
            .I(N__53821));
    InMux I__11786 (
            .O(N__53821),
            .I(N__53818));
    LocalMux I__11785 (
            .O(N__53818),
            .I(N__53815));
    Span4Mux_h I__11784 (
            .O(N__53815),
            .I(N__53812));
    Odrv4 I__11783 (
            .O(N__53812),
            .I(\c0.n21767 ));
    InMux I__11782 (
            .O(N__53809),
            .I(N__53805));
    InMux I__11781 (
            .O(N__53808),
            .I(N__53801));
    LocalMux I__11780 (
            .O(N__53805),
            .I(N__53798));
    InMux I__11779 (
            .O(N__53804),
            .I(N__53795));
    LocalMux I__11778 (
            .O(N__53801),
            .I(N__53791));
    Span4Mux_v I__11777 (
            .O(N__53798),
            .I(N__53786));
    LocalMux I__11776 (
            .O(N__53795),
            .I(N__53786));
    InMux I__11775 (
            .O(N__53794),
            .I(N__53783));
    Span12Mux_v I__11774 (
            .O(N__53791),
            .I(N__53780));
    Span4Mux_v I__11773 (
            .O(N__53786),
            .I(N__53777));
    LocalMux I__11772 (
            .O(N__53783),
            .I(data_in_frame_22_6));
    Odrv12 I__11771 (
            .O(N__53780),
            .I(data_in_frame_22_6));
    Odrv4 I__11770 (
            .O(N__53777),
            .I(data_in_frame_22_6));
    InMux I__11769 (
            .O(N__53770),
            .I(N__53765));
    InMux I__11768 (
            .O(N__53769),
            .I(N__53760));
    InMux I__11767 (
            .O(N__53768),
            .I(N__53760));
    LocalMux I__11766 (
            .O(N__53765),
            .I(data_in_frame_23_0));
    LocalMux I__11765 (
            .O(N__53760),
            .I(data_in_frame_23_0));
    InMux I__11764 (
            .O(N__53755),
            .I(N__53752));
    LocalMux I__11763 (
            .O(N__53752),
            .I(N__53748));
    InMux I__11762 (
            .O(N__53751),
            .I(N__53745));
    Span4Mux_v I__11761 (
            .O(N__53748),
            .I(N__53741));
    LocalMux I__11760 (
            .O(N__53745),
            .I(N__53738));
    InMux I__11759 (
            .O(N__53744),
            .I(N__53735));
    Span4Mux_h I__11758 (
            .O(N__53741),
            .I(N__53732));
    Span4Mux_v I__11757 (
            .O(N__53738),
            .I(N__53729));
    LocalMux I__11756 (
            .O(N__53735),
            .I(data_in_frame_23_4));
    Odrv4 I__11755 (
            .O(N__53732),
            .I(data_in_frame_23_4));
    Odrv4 I__11754 (
            .O(N__53729),
            .I(data_in_frame_23_4));
    InMux I__11753 (
            .O(N__53722),
            .I(N__53715));
    InMux I__11752 (
            .O(N__53721),
            .I(N__53715));
    InMux I__11751 (
            .O(N__53720),
            .I(N__53711));
    LocalMux I__11750 (
            .O(N__53715),
            .I(N__53706));
    InMux I__11749 (
            .O(N__53714),
            .I(N__53703));
    LocalMux I__11748 (
            .O(N__53711),
            .I(N__53699));
    InMux I__11747 (
            .O(N__53710),
            .I(N__53694));
    InMux I__11746 (
            .O(N__53709),
            .I(N__53694));
    Span4Mux_v I__11745 (
            .O(N__53706),
            .I(N__53688));
    LocalMux I__11744 (
            .O(N__53703),
            .I(N__53688));
    InMux I__11743 (
            .O(N__53702),
            .I(N__53685));
    Span12Mux_v I__11742 (
            .O(N__53699),
            .I(N__53682));
    LocalMux I__11741 (
            .O(N__53694),
            .I(N__53679));
    InMux I__11740 (
            .O(N__53693),
            .I(N__53676));
    Span4Mux_h I__11739 (
            .O(N__53688),
            .I(N__53671));
    LocalMux I__11738 (
            .O(N__53685),
            .I(N__53671));
    Odrv12 I__11737 (
            .O(N__53682),
            .I(n19126));
    Odrv12 I__11736 (
            .O(N__53679),
            .I(n19126));
    LocalMux I__11735 (
            .O(N__53676),
            .I(n19126));
    Odrv4 I__11734 (
            .O(N__53671),
            .I(n19126));
    CascadeMux I__11733 (
            .O(N__53662),
            .I(N__53659));
    InMux I__11732 (
            .O(N__53659),
            .I(N__53654));
    CascadeMux I__11731 (
            .O(N__53658),
            .I(N__53651));
    CascadeMux I__11730 (
            .O(N__53657),
            .I(N__53648));
    LocalMux I__11729 (
            .O(N__53654),
            .I(N__53645));
    InMux I__11728 (
            .O(N__53651),
            .I(N__53642));
    InMux I__11727 (
            .O(N__53648),
            .I(N__53639));
    Span4Mux_h I__11726 (
            .O(N__53645),
            .I(N__53636));
    LocalMux I__11725 (
            .O(N__53642),
            .I(N__53633));
    LocalMux I__11724 (
            .O(N__53639),
            .I(\c0.data_in_frame_11_0 ));
    Odrv4 I__11723 (
            .O(N__53636),
            .I(\c0.data_in_frame_11_0 ));
    Odrv4 I__11722 (
            .O(N__53633),
            .I(\c0.data_in_frame_11_0 ));
    InMux I__11721 (
            .O(N__53626),
            .I(N__53623));
    LocalMux I__11720 (
            .O(N__53623),
            .I(N__53619));
    InMux I__11719 (
            .O(N__53622),
            .I(N__53615));
    Span4Mux_v I__11718 (
            .O(N__53619),
            .I(N__53612));
    InMux I__11717 (
            .O(N__53618),
            .I(N__53609));
    LocalMux I__11716 (
            .O(N__53615),
            .I(data_in_frame_24_7));
    Odrv4 I__11715 (
            .O(N__53612),
            .I(data_in_frame_24_7));
    LocalMux I__11714 (
            .O(N__53609),
            .I(data_in_frame_24_7));
    InMux I__11713 (
            .O(N__53602),
            .I(N__53598));
    InMux I__11712 (
            .O(N__53601),
            .I(N__53595));
    LocalMux I__11711 (
            .O(N__53598),
            .I(N__53592));
    LocalMux I__11710 (
            .O(N__53595),
            .I(\c0.n12206 ));
    Odrv4 I__11709 (
            .O(N__53592),
            .I(\c0.n12206 ));
    InMux I__11708 (
            .O(N__53587),
            .I(N__53582));
    InMux I__11707 (
            .O(N__53586),
            .I(N__53579));
    InMux I__11706 (
            .O(N__53585),
            .I(N__53576));
    LocalMux I__11705 (
            .O(N__53582),
            .I(N__53573));
    LocalMux I__11704 (
            .O(N__53579),
            .I(N__53570));
    LocalMux I__11703 (
            .O(N__53576),
            .I(\c0.n19268 ));
    Odrv4 I__11702 (
            .O(N__53573),
            .I(\c0.n19268 ));
    Odrv12 I__11701 (
            .O(N__53570),
            .I(\c0.n19268 ));
    CascadeMux I__11700 (
            .O(N__53563),
            .I(\c0.n19268_cascade_ ));
    InMux I__11699 (
            .O(N__53560),
            .I(N__53557));
    LocalMux I__11698 (
            .O(N__53557),
            .I(N__53553));
    InMux I__11697 (
            .O(N__53556),
            .I(N__53550));
    Span4Mux_v I__11696 (
            .O(N__53553),
            .I(N__53545));
    LocalMux I__11695 (
            .O(N__53550),
            .I(N__53545));
    Span4Mux_h I__11694 (
            .O(N__53545),
            .I(N__53542));
    Odrv4 I__11693 (
            .O(N__53542),
            .I(\c0.n20_adj_3301 ));
    InMux I__11692 (
            .O(N__53539),
            .I(N__53532));
    InMux I__11691 (
            .O(N__53538),
            .I(N__53532));
    InMux I__11690 (
            .O(N__53537),
            .I(N__53529));
    LocalMux I__11689 (
            .O(N__53532),
            .I(N__53526));
    LocalMux I__11688 (
            .O(N__53529),
            .I(N__53523));
    Span4Mux_v I__11687 (
            .O(N__53526),
            .I(N__53520));
    Span4Mux_v I__11686 (
            .O(N__53523),
            .I(N__53517));
    Odrv4 I__11685 (
            .O(N__53520),
            .I(\c0.n7_adj_3054 ));
    Odrv4 I__11684 (
            .O(N__53517),
            .I(\c0.n7_adj_3054 ));
    InMux I__11683 (
            .O(N__53512),
            .I(N__53507));
    InMux I__11682 (
            .O(N__53511),
            .I(N__53501));
    InMux I__11681 (
            .O(N__53510),
            .I(N__53501));
    LocalMux I__11680 (
            .O(N__53507),
            .I(N__53498));
    InMux I__11679 (
            .O(N__53506),
            .I(N__53495));
    LocalMux I__11678 (
            .O(N__53501),
            .I(N__53491));
    Span4Mux_v I__11677 (
            .O(N__53498),
            .I(N__53488));
    LocalMux I__11676 (
            .O(N__53495),
            .I(N__53485));
    InMux I__11675 (
            .O(N__53494),
            .I(N__53482));
    Odrv4 I__11674 (
            .O(N__53491),
            .I(\c0.n11601 ));
    Odrv4 I__11673 (
            .O(N__53488),
            .I(\c0.n11601 ));
    Odrv4 I__11672 (
            .O(N__53485),
            .I(\c0.n11601 ));
    LocalMux I__11671 (
            .O(N__53482),
            .I(\c0.n11601 ));
    InMux I__11670 (
            .O(N__53473),
            .I(N__53470));
    LocalMux I__11669 (
            .O(N__53470),
            .I(N__53466));
    InMux I__11668 (
            .O(N__53469),
            .I(N__53463));
    Span4Mux_v I__11667 (
            .O(N__53466),
            .I(N__53460));
    LocalMux I__11666 (
            .O(N__53463),
            .I(N__53456));
    Span4Mux_h I__11665 (
            .O(N__53460),
            .I(N__53453));
    InMux I__11664 (
            .O(N__53459),
            .I(N__53450));
    Odrv12 I__11663 (
            .O(N__53456),
            .I(\c0.n19764 ));
    Odrv4 I__11662 (
            .O(N__53453),
            .I(\c0.n19764 ));
    LocalMux I__11661 (
            .O(N__53450),
            .I(\c0.n19764 ));
    InMux I__11660 (
            .O(N__53443),
            .I(N__53439));
    InMux I__11659 (
            .O(N__53442),
            .I(N__53436));
    LocalMux I__11658 (
            .O(N__53439),
            .I(N__53433));
    LocalMux I__11657 (
            .O(N__53436),
            .I(N__53430));
    Odrv4 I__11656 (
            .O(N__53433),
            .I(\c0.n42_adj_3055 ));
    Odrv12 I__11655 (
            .O(N__53430),
            .I(\c0.n42_adj_3055 ));
    InMux I__11654 (
            .O(N__53425),
            .I(N__53422));
    LocalMux I__11653 (
            .O(N__53422),
            .I(N__53418));
    InMux I__11652 (
            .O(N__53421),
            .I(N__53415));
    Span4Mux_v I__11651 (
            .O(N__53418),
            .I(N__53409));
    LocalMux I__11650 (
            .O(N__53415),
            .I(N__53409));
    InMux I__11649 (
            .O(N__53414),
            .I(N__53406));
    Span4Mux_v I__11648 (
            .O(N__53409),
            .I(N__53403));
    LocalMux I__11647 (
            .O(N__53406),
            .I(N__53400));
    Odrv4 I__11646 (
            .O(N__53403),
            .I(\c0.n11815 ));
    Odrv4 I__11645 (
            .O(N__53400),
            .I(\c0.n11815 ));
    CascadeMux I__11644 (
            .O(N__53395),
            .I(N__53392));
    InMux I__11643 (
            .O(N__53392),
            .I(N__53386));
    InMux I__11642 (
            .O(N__53391),
            .I(N__53386));
    LocalMux I__11641 (
            .O(N__53386),
            .I(\c0.n4_adj_3100 ));
    InMux I__11640 (
            .O(N__53383),
            .I(N__53380));
    LocalMux I__11639 (
            .O(N__53380),
            .I(N__53376));
    CascadeMux I__11638 (
            .O(N__53379),
            .I(N__53372));
    Span4Mux_v I__11637 (
            .O(N__53376),
            .I(N__53369));
    InMux I__11636 (
            .O(N__53375),
            .I(N__53366));
    InMux I__11635 (
            .O(N__53372),
            .I(N__53363));
    Sp12to4 I__11634 (
            .O(N__53369),
            .I(N__53358));
    LocalMux I__11633 (
            .O(N__53366),
            .I(N__53358));
    LocalMux I__11632 (
            .O(N__53363),
            .I(\c0.data_in_frame_25_0 ));
    Odrv12 I__11631 (
            .O(N__53358),
            .I(\c0.data_in_frame_25_0 ));
    InMux I__11630 (
            .O(N__53353),
            .I(N__53350));
    LocalMux I__11629 (
            .O(N__53350),
            .I(N__53347));
    Odrv4 I__11628 (
            .O(N__53347),
            .I(\c0.n19436 ));
    InMux I__11627 (
            .O(N__53344),
            .I(N__53339));
    InMux I__11626 (
            .O(N__53343),
            .I(N__53334));
    InMux I__11625 (
            .O(N__53342),
            .I(N__53334));
    LocalMux I__11624 (
            .O(N__53339),
            .I(N__53330));
    LocalMux I__11623 (
            .O(N__53334),
            .I(N__53327));
    InMux I__11622 (
            .O(N__53333),
            .I(N__53322));
    Span4Mux_v I__11621 (
            .O(N__53330),
            .I(N__53319));
    Span4Mux_h I__11620 (
            .O(N__53327),
            .I(N__53316));
    InMux I__11619 (
            .O(N__53326),
            .I(N__53311));
    InMux I__11618 (
            .O(N__53325),
            .I(N__53311));
    LocalMux I__11617 (
            .O(N__53322),
            .I(data_in_frame_22_4));
    Odrv4 I__11616 (
            .O(N__53319),
            .I(data_in_frame_22_4));
    Odrv4 I__11615 (
            .O(N__53316),
            .I(data_in_frame_22_4));
    LocalMux I__11614 (
            .O(N__53311),
            .I(data_in_frame_22_4));
    CascadeMux I__11613 (
            .O(N__53302),
            .I(\c0.n19436_cascade_ ));
    InMux I__11612 (
            .O(N__53299),
            .I(N__53294));
    InMux I__11611 (
            .O(N__53298),
            .I(N__53289));
    InMux I__11610 (
            .O(N__53297),
            .I(N__53289));
    LocalMux I__11609 (
            .O(N__53294),
            .I(\c0.n11776 ));
    LocalMux I__11608 (
            .O(N__53289),
            .I(\c0.n11776 ));
    CascadeMux I__11607 (
            .O(N__53284),
            .I(N__53281));
    InMux I__11606 (
            .O(N__53281),
            .I(N__53275));
    InMux I__11605 (
            .O(N__53280),
            .I(N__53275));
    LocalMux I__11604 (
            .O(N__53275),
            .I(\c0.n6_adj_3112 ));
    InMux I__11603 (
            .O(N__53272),
            .I(N__53266));
    InMux I__11602 (
            .O(N__53271),
            .I(N__53266));
    LocalMux I__11601 (
            .O(N__53266),
            .I(\c0.n19151 ));
    InMux I__11600 (
            .O(N__53263),
            .I(N__53260));
    LocalMux I__11599 (
            .O(N__53260),
            .I(N__53256));
    InMux I__11598 (
            .O(N__53259),
            .I(N__53252));
    Span4Mux_h I__11597 (
            .O(N__53256),
            .I(N__53249));
    InMux I__11596 (
            .O(N__53255),
            .I(N__53246));
    LocalMux I__11595 (
            .O(N__53252),
            .I(N__53243));
    Span4Mux_h I__11594 (
            .O(N__53249),
            .I(N__53238));
    LocalMux I__11593 (
            .O(N__53246),
            .I(N__53238));
    Span12Mux_h I__11592 (
            .O(N__53243),
            .I(N__53235));
    Odrv4 I__11591 (
            .O(N__53238),
            .I(\c0.n20933 ));
    Odrv12 I__11590 (
            .O(N__53235),
            .I(\c0.n20933 ));
    InMux I__11589 (
            .O(N__53230),
            .I(N__53212));
    InMux I__11588 (
            .O(N__53229),
            .I(N__53205));
    InMux I__11587 (
            .O(N__53228),
            .I(N__53202));
    InMux I__11586 (
            .O(N__53227),
            .I(N__53199));
    InMux I__11585 (
            .O(N__53226),
            .I(N__53196));
    InMux I__11584 (
            .O(N__53225),
            .I(N__53192));
    CascadeMux I__11583 (
            .O(N__53224),
            .I(N__53189));
    InMux I__11582 (
            .O(N__53223),
            .I(N__53180));
    InMux I__11581 (
            .O(N__53222),
            .I(N__53180));
    InMux I__11580 (
            .O(N__53221),
            .I(N__53180));
    InMux I__11579 (
            .O(N__53220),
            .I(N__53165));
    InMux I__11578 (
            .O(N__53219),
            .I(N__53165));
    InMux I__11577 (
            .O(N__53218),
            .I(N__53165));
    InMux I__11576 (
            .O(N__53217),
            .I(N__53160));
    InMux I__11575 (
            .O(N__53216),
            .I(N__53160));
    InMux I__11574 (
            .O(N__53215),
            .I(N__53157));
    LocalMux I__11573 (
            .O(N__53212),
            .I(N__53154));
    InMux I__11572 (
            .O(N__53211),
            .I(N__53145));
    InMux I__11571 (
            .O(N__53210),
            .I(N__53145));
    InMux I__11570 (
            .O(N__53209),
            .I(N__53145));
    InMux I__11569 (
            .O(N__53208),
            .I(N__53145));
    LocalMux I__11568 (
            .O(N__53205),
            .I(N__53136));
    LocalMux I__11567 (
            .O(N__53202),
            .I(N__53136));
    LocalMux I__11566 (
            .O(N__53199),
            .I(N__53136));
    LocalMux I__11565 (
            .O(N__53196),
            .I(N__53136));
    InMux I__11564 (
            .O(N__53195),
            .I(N__53132));
    LocalMux I__11563 (
            .O(N__53192),
            .I(N__53129));
    InMux I__11562 (
            .O(N__53189),
            .I(N__53122));
    InMux I__11561 (
            .O(N__53188),
            .I(N__53122));
    InMux I__11560 (
            .O(N__53187),
            .I(N__53122));
    LocalMux I__11559 (
            .O(N__53180),
            .I(N__53119));
    InMux I__11558 (
            .O(N__53179),
            .I(N__53115));
    InMux I__11557 (
            .O(N__53178),
            .I(N__53112));
    InMux I__11556 (
            .O(N__53177),
            .I(N__53109));
    InMux I__11555 (
            .O(N__53176),
            .I(N__53106));
    InMux I__11554 (
            .O(N__53175),
            .I(N__53103));
    InMux I__11553 (
            .O(N__53174),
            .I(N__53100));
    InMux I__11552 (
            .O(N__53173),
            .I(N__53095));
    InMux I__11551 (
            .O(N__53172),
            .I(N__53095));
    LocalMux I__11550 (
            .O(N__53165),
            .I(N__53092));
    LocalMux I__11549 (
            .O(N__53160),
            .I(N__53087));
    LocalMux I__11548 (
            .O(N__53157),
            .I(N__53087));
    Span4Mux_h I__11547 (
            .O(N__53154),
            .I(N__53080));
    LocalMux I__11546 (
            .O(N__53145),
            .I(N__53080));
    Span4Mux_v I__11545 (
            .O(N__53136),
            .I(N__53080));
    InMux I__11544 (
            .O(N__53135),
            .I(N__53076));
    LocalMux I__11543 (
            .O(N__53132),
            .I(N__53071));
    Span4Mux_h I__11542 (
            .O(N__53129),
            .I(N__53071));
    LocalMux I__11541 (
            .O(N__53122),
            .I(N__53066));
    Span4Mux_v I__11540 (
            .O(N__53119),
            .I(N__53066));
    CascadeMux I__11539 (
            .O(N__53118),
            .I(N__53063));
    LocalMux I__11538 (
            .O(N__53115),
            .I(N__53060));
    LocalMux I__11537 (
            .O(N__53112),
            .I(N__53055));
    LocalMux I__11536 (
            .O(N__53109),
            .I(N__53055));
    LocalMux I__11535 (
            .O(N__53106),
            .I(N__53040));
    LocalMux I__11534 (
            .O(N__53103),
            .I(N__53040));
    LocalMux I__11533 (
            .O(N__53100),
            .I(N__53040));
    LocalMux I__11532 (
            .O(N__53095),
            .I(N__53040));
    Span4Mux_h I__11531 (
            .O(N__53092),
            .I(N__53040));
    Span4Mux_v I__11530 (
            .O(N__53087),
            .I(N__53040));
    Span4Mux_h I__11529 (
            .O(N__53080),
            .I(N__53040));
    InMux I__11528 (
            .O(N__53079),
            .I(N__53037));
    LocalMux I__11527 (
            .O(N__53076),
            .I(N__53033));
    Span4Mux_v I__11526 (
            .O(N__53071),
            .I(N__53030));
    Span4Mux_v I__11525 (
            .O(N__53066),
            .I(N__53027));
    InMux I__11524 (
            .O(N__53063),
            .I(N__53024));
    Span4Mux_h I__11523 (
            .O(N__53060),
            .I(N__53015));
    Span4Mux_v I__11522 (
            .O(N__53055),
            .I(N__53015));
    Span4Mux_v I__11521 (
            .O(N__53040),
            .I(N__53015));
    LocalMux I__11520 (
            .O(N__53037),
            .I(N__53015));
    CascadeMux I__11519 (
            .O(N__53036),
            .I(N__53012));
    Sp12to4 I__11518 (
            .O(N__53033),
            .I(N__53008));
    Span4Mux_v I__11517 (
            .O(N__53030),
            .I(N__53005));
    Span4Mux_v I__11516 (
            .O(N__53027),
            .I(N__53000));
    LocalMux I__11515 (
            .O(N__53024),
            .I(N__53000));
    Span4Mux_v I__11514 (
            .O(N__53015),
            .I(N__52997));
    InMux I__11513 (
            .O(N__53012),
            .I(N__52993));
    InMux I__11512 (
            .O(N__53011),
            .I(N__52990));
    Span12Mux_v I__11511 (
            .O(N__53008),
            .I(N__52987));
    Span4Mux_v I__11510 (
            .O(N__53005),
            .I(N__52984));
    Span4Mux_v I__11509 (
            .O(N__53000),
            .I(N__52981));
    Span4Mux_v I__11508 (
            .O(N__52997),
            .I(N__52978));
    InMux I__11507 (
            .O(N__52996),
            .I(N__52975));
    LocalMux I__11506 (
            .O(N__52993),
            .I(rx_data_ready));
    LocalMux I__11505 (
            .O(N__52990),
            .I(rx_data_ready));
    Odrv12 I__11504 (
            .O(N__52987),
            .I(rx_data_ready));
    Odrv4 I__11503 (
            .O(N__52984),
            .I(rx_data_ready));
    Odrv4 I__11502 (
            .O(N__52981),
            .I(rx_data_ready));
    Odrv4 I__11501 (
            .O(N__52978),
            .I(rx_data_ready));
    LocalMux I__11500 (
            .O(N__52975),
            .I(rx_data_ready));
    InMux I__11499 (
            .O(N__52960),
            .I(N__52957));
    LocalMux I__11498 (
            .O(N__52957),
            .I(N__52953));
    CascadeMux I__11497 (
            .O(N__52956),
            .I(N__52950));
    Span4Mux_h I__11496 (
            .O(N__52953),
            .I(N__52946));
    InMux I__11495 (
            .O(N__52950),
            .I(N__52943));
    InMux I__11494 (
            .O(N__52949),
            .I(N__52939));
    Span4Mux_h I__11493 (
            .O(N__52946),
            .I(N__52936));
    LocalMux I__11492 (
            .O(N__52943),
            .I(N__52933));
    InMux I__11491 (
            .O(N__52942),
            .I(N__52930));
    LocalMux I__11490 (
            .O(N__52939),
            .I(data_in_3_6));
    Odrv4 I__11489 (
            .O(N__52936),
            .I(data_in_3_6));
    Odrv4 I__11488 (
            .O(N__52933),
            .I(data_in_3_6));
    LocalMux I__11487 (
            .O(N__52930),
            .I(data_in_3_6));
    CascadeMux I__11486 (
            .O(N__52921),
            .I(N__52916));
    InMux I__11485 (
            .O(N__52920),
            .I(N__52913));
    InMux I__11484 (
            .O(N__52919),
            .I(N__52910));
    InMux I__11483 (
            .O(N__52916),
            .I(N__52907));
    LocalMux I__11482 (
            .O(N__52913),
            .I(N__52904));
    LocalMux I__11481 (
            .O(N__52910),
            .I(N__52900));
    LocalMux I__11480 (
            .O(N__52907),
            .I(N__52895));
    Span4Mux_h I__11479 (
            .O(N__52904),
            .I(N__52895));
    InMux I__11478 (
            .O(N__52903),
            .I(N__52892));
    Span12Mux_h I__11477 (
            .O(N__52900),
            .I(N__52889));
    Span4Mux_h I__11476 (
            .O(N__52895),
            .I(N__52886));
    LocalMux I__11475 (
            .O(N__52892),
            .I(data_in_2_6));
    Odrv12 I__11474 (
            .O(N__52889),
            .I(data_in_2_6));
    Odrv4 I__11473 (
            .O(N__52886),
            .I(data_in_2_6));
    InMux I__11472 (
            .O(N__52879),
            .I(N__52876));
    LocalMux I__11471 (
            .O(N__52876),
            .I(N__52872));
    InMux I__11470 (
            .O(N__52875),
            .I(N__52869));
    Odrv4 I__11469 (
            .O(N__52872),
            .I(\c0.n24_adj_3427 ));
    LocalMux I__11468 (
            .O(N__52869),
            .I(\c0.n24_adj_3427 ));
    InMux I__11467 (
            .O(N__52864),
            .I(N__52859));
    InMux I__11466 (
            .O(N__52863),
            .I(N__52854));
    InMux I__11465 (
            .O(N__52862),
            .I(N__52854));
    LocalMux I__11464 (
            .O(N__52859),
            .I(N__52849));
    LocalMux I__11463 (
            .O(N__52854),
            .I(N__52849));
    Span4Mux_v I__11462 (
            .O(N__52849),
            .I(N__52846));
    Odrv4 I__11461 (
            .O(N__52846),
            .I(\c0.n11714 ));
    InMux I__11460 (
            .O(N__52843),
            .I(N__52840));
    LocalMux I__11459 (
            .O(N__52840),
            .I(N__52837));
    Span4Mux_h I__11458 (
            .O(N__52837),
            .I(N__52834));
    Odrv4 I__11457 (
            .O(N__52834),
            .I(\c0.n22_adj_3296 ));
    CascadeMux I__11456 (
            .O(N__52831),
            .I(\c0.n19159_cascade_ ));
    InMux I__11455 (
            .O(N__52828),
            .I(N__52824));
    InMux I__11454 (
            .O(N__52827),
            .I(N__52821));
    LocalMux I__11453 (
            .O(N__52824),
            .I(N__52818));
    LocalMux I__11452 (
            .O(N__52821),
            .I(N__52815));
    Span4Mux_v I__11451 (
            .O(N__52818),
            .I(N__52812));
    Span4Mux_h I__11450 (
            .O(N__52815),
            .I(N__52809));
    Odrv4 I__11449 (
            .O(N__52812),
            .I(\c0.n11632 ));
    Odrv4 I__11448 (
            .O(N__52809),
            .I(\c0.n11632 ));
    InMux I__11447 (
            .O(N__52804),
            .I(N__52801));
    LocalMux I__11446 (
            .O(N__52801),
            .I(\c0.n19159 ));
    CascadeMux I__11445 (
            .O(N__52798),
            .I(N__52795));
    InMux I__11444 (
            .O(N__52795),
            .I(N__52791));
    CascadeMux I__11443 (
            .O(N__52794),
            .I(N__52788));
    LocalMux I__11442 (
            .O(N__52791),
            .I(N__52785));
    InMux I__11441 (
            .O(N__52788),
            .I(N__52782));
    Span4Mux_v I__11440 (
            .O(N__52785),
            .I(N__52779));
    LocalMux I__11439 (
            .O(N__52782),
            .I(\c0.data_in_frame_28_7 ));
    Odrv4 I__11438 (
            .O(N__52779),
            .I(\c0.data_in_frame_28_7 ));
    InMux I__11437 (
            .O(N__52774),
            .I(N__52771));
    LocalMux I__11436 (
            .O(N__52771),
            .I(N__52768));
    Span4Mux_h I__11435 (
            .O(N__52768),
            .I(N__52765));
    Odrv4 I__11434 (
            .O(N__52765),
            .I(\c0.n79 ));
    InMux I__11433 (
            .O(N__52762),
            .I(N__52759));
    LocalMux I__11432 (
            .O(N__52759),
            .I(N__52755));
    InMux I__11431 (
            .O(N__52758),
            .I(N__52752));
    Span12Mux_h I__11430 (
            .O(N__52755),
            .I(N__52749));
    LocalMux I__11429 (
            .O(N__52752),
            .I(N__52746));
    Span12Mux_v I__11428 (
            .O(N__52749),
            .I(N__52743));
    Span4Mux_v I__11427 (
            .O(N__52746),
            .I(N__52740));
    Odrv12 I__11426 (
            .O(N__52743),
            .I(\c0.n10_adj_3207 ));
    Odrv4 I__11425 (
            .O(N__52740),
            .I(\c0.n10_adj_3207 ));
    InMux I__11424 (
            .O(N__52735),
            .I(N__52729));
    InMux I__11423 (
            .O(N__52734),
            .I(N__52729));
    LocalMux I__11422 (
            .O(N__52729),
            .I(N__52726));
    Span4Mux_v I__11421 (
            .O(N__52726),
            .I(N__52723));
    Span4Mux_h I__11420 (
            .O(N__52723),
            .I(N__52719));
    InMux I__11419 (
            .O(N__52722),
            .I(N__52716));
    Odrv4 I__11418 (
            .O(N__52719),
            .I(\c0.n11_adj_3206 ));
    LocalMux I__11417 (
            .O(N__52716),
            .I(\c0.n11_adj_3206 ));
    CascadeMux I__11416 (
            .O(N__52711),
            .I(\c0.n11776_cascade_ ));
    InMux I__11415 (
            .O(N__52708),
            .I(N__52703));
    InMux I__11414 (
            .O(N__52707),
            .I(N__52698));
    InMux I__11413 (
            .O(N__52706),
            .I(N__52698));
    LocalMux I__11412 (
            .O(N__52703),
            .I(\c0.n6_adj_3319 ));
    LocalMux I__11411 (
            .O(N__52698),
            .I(\c0.n6_adj_3319 ));
    CascadeMux I__11410 (
            .O(N__52693),
            .I(\c0.n70_adj_3087_cascade_ ));
    InMux I__11409 (
            .O(N__52690),
            .I(N__52686));
    InMux I__11408 (
            .O(N__52689),
            .I(N__52683));
    LocalMux I__11407 (
            .O(N__52686),
            .I(N__52678));
    LocalMux I__11406 (
            .O(N__52683),
            .I(N__52678));
    Span4Mux_v I__11405 (
            .O(N__52678),
            .I(N__52675));
    Odrv4 I__11404 (
            .O(N__52675),
            .I(\c0.n20339 ));
    InMux I__11403 (
            .O(N__52672),
            .I(N__52668));
    InMux I__11402 (
            .O(N__52671),
            .I(N__52665));
    LocalMux I__11401 (
            .O(N__52668),
            .I(N__52662));
    LocalMux I__11400 (
            .O(N__52665),
            .I(N__52657));
    Span4Mux_h I__11399 (
            .O(N__52662),
            .I(N__52657));
    Span4Mux_h I__11398 (
            .O(N__52657),
            .I(N__52654));
    Odrv4 I__11397 (
            .O(N__52654),
            .I(\c0.n27_adj_3311 ));
    InMux I__11396 (
            .O(N__52651),
            .I(N__52648));
    LocalMux I__11395 (
            .O(N__52648),
            .I(N__52642));
    InMux I__11394 (
            .O(N__52647),
            .I(N__52637));
    InMux I__11393 (
            .O(N__52646),
            .I(N__52637));
    InMux I__11392 (
            .O(N__52645),
            .I(N__52634));
    Span4Mux_v I__11391 (
            .O(N__52642),
            .I(N__52629));
    LocalMux I__11390 (
            .O(N__52637),
            .I(N__52629));
    LocalMux I__11389 (
            .O(N__52634),
            .I(N__52626));
    Span4Mux_h I__11388 (
            .O(N__52629),
            .I(N__52623));
    Span4Mux_v I__11387 (
            .O(N__52626),
            .I(N__52620));
    Odrv4 I__11386 (
            .O(N__52623),
            .I(\c0.n7_adj_3094 ));
    Odrv4 I__11385 (
            .O(N__52620),
            .I(\c0.n7_adj_3094 ));
    InMux I__11384 (
            .O(N__52615),
            .I(N__52612));
    LocalMux I__11383 (
            .O(N__52612),
            .I(N__52609));
    Odrv4 I__11382 (
            .O(N__52609),
            .I(\c0.n20_adj_3293 ));
    InMux I__11381 (
            .O(N__52606),
            .I(N__52603));
    LocalMux I__11380 (
            .O(N__52603),
            .I(N__52600));
    Span4Mux_h I__11379 (
            .O(N__52600),
            .I(N__52596));
    InMux I__11378 (
            .O(N__52599),
            .I(N__52593));
    Odrv4 I__11377 (
            .O(N__52596),
            .I(\c0.n33_adj_3279 ));
    LocalMux I__11376 (
            .O(N__52593),
            .I(\c0.n33_adj_3279 ));
    InMux I__11375 (
            .O(N__52588),
            .I(N__52585));
    LocalMux I__11374 (
            .O(N__52585),
            .I(\c0.n30_adj_3295 ));
    CascadeMux I__11373 (
            .O(N__52582),
            .I(\c0.n32_adj_3294_cascade_ ));
    InMux I__11372 (
            .O(N__52579),
            .I(N__52576));
    LocalMux I__11371 (
            .O(N__52576),
            .I(N__52573));
    Span4Mux_v I__11370 (
            .O(N__52573),
            .I(N__52570));
    Odrv4 I__11369 (
            .O(N__52570),
            .I(\c0.n21075 ));
    InMux I__11368 (
            .O(N__52567),
            .I(N__52564));
    LocalMux I__11367 (
            .O(N__52564),
            .I(N__52560));
    InMux I__11366 (
            .O(N__52563),
            .I(N__52556));
    Span4Mux_h I__11365 (
            .O(N__52560),
            .I(N__52553));
    InMux I__11364 (
            .O(N__52559),
            .I(N__52550));
    LocalMux I__11363 (
            .O(N__52556),
            .I(N__52547));
    Span4Mux_v I__11362 (
            .O(N__52553),
            .I(N__52544));
    LocalMux I__11361 (
            .O(N__52550),
            .I(N__52540));
    Span4Mux_v I__11360 (
            .O(N__52547),
            .I(N__52535));
    Span4Mux_h I__11359 (
            .O(N__52544),
            .I(N__52535));
    InMux I__11358 (
            .O(N__52543),
            .I(N__52532));
    Odrv4 I__11357 (
            .O(N__52540),
            .I(\c0.n7_adj_3079 ));
    Odrv4 I__11356 (
            .O(N__52535),
            .I(\c0.n7_adj_3079 ));
    LocalMux I__11355 (
            .O(N__52532),
            .I(\c0.n7_adj_3079 ));
    InMux I__11354 (
            .O(N__52525),
            .I(N__52522));
    LocalMux I__11353 (
            .O(N__52522),
            .I(\c0.n29_adj_3299 ));
    InMux I__11352 (
            .O(N__52519),
            .I(N__52516));
    LocalMux I__11351 (
            .O(N__52516),
            .I(N__52513));
    Span4Mux_v I__11350 (
            .O(N__52513),
            .I(N__52510));
    Odrv4 I__11349 (
            .O(N__52510),
            .I(\c0.n19_adj_3320 ));
    InMux I__11348 (
            .O(N__52507),
            .I(N__52500));
    InMux I__11347 (
            .O(N__52506),
            .I(N__52500));
    InMux I__11346 (
            .O(N__52505),
            .I(N__52497));
    LocalMux I__11345 (
            .O(N__52500),
            .I(\c0.n20336 ));
    LocalMux I__11344 (
            .O(N__52497),
            .I(\c0.n20336 ));
    CascadeMux I__11343 (
            .O(N__52492),
            .I(N__52486));
    InMux I__11342 (
            .O(N__52491),
            .I(N__52483));
    CascadeMux I__11341 (
            .O(N__52490),
            .I(N__52479));
    CascadeMux I__11340 (
            .O(N__52489),
            .I(N__52476));
    InMux I__11339 (
            .O(N__52486),
            .I(N__52473));
    LocalMux I__11338 (
            .O(N__52483),
            .I(N__52470));
    InMux I__11337 (
            .O(N__52482),
            .I(N__52467));
    InMux I__11336 (
            .O(N__52479),
            .I(N__52462));
    InMux I__11335 (
            .O(N__52476),
            .I(N__52462));
    LocalMux I__11334 (
            .O(N__52473),
            .I(N__52459));
    Span4Mux_h I__11333 (
            .O(N__52470),
            .I(N__52454));
    LocalMux I__11332 (
            .O(N__52467),
            .I(N__52454));
    LocalMux I__11331 (
            .O(N__52462),
            .I(\c0.n18379 ));
    Odrv4 I__11330 (
            .O(N__52459),
            .I(\c0.n18379 ));
    Odrv4 I__11329 (
            .O(N__52454),
            .I(\c0.n18379 ));
    InMux I__11328 (
            .O(N__52447),
            .I(N__52441));
    InMux I__11327 (
            .O(N__52446),
            .I(N__52438));
    InMux I__11326 (
            .O(N__52445),
            .I(N__52435));
    InMux I__11325 (
            .O(N__52444),
            .I(N__52432));
    LocalMux I__11324 (
            .O(N__52441),
            .I(\c0.n21034 ));
    LocalMux I__11323 (
            .O(N__52438),
            .I(\c0.n21034 ));
    LocalMux I__11322 (
            .O(N__52435),
            .I(\c0.n21034 ));
    LocalMux I__11321 (
            .O(N__52432),
            .I(\c0.n21034 ));
    InMux I__11320 (
            .O(N__52423),
            .I(N__52420));
    LocalMux I__11319 (
            .O(N__52420),
            .I(N__52417));
    Span4Mux_h I__11318 (
            .O(N__52417),
            .I(N__52413));
    InMux I__11317 (
            .O(N__52416),
            .I(N__52410));
    Odrv4 I__11316 (
            .O(N__52413),
            .I(\c0.n57 ));
    LocalMux I__11315 (
            .O(N__52410),
            .I(\c0.n57 ));
    InMux I__11314 (
            .O(N__52405),
            .I(N__52402));
    LocalMux I__11313 (
            .O(N__52402),
            .I(\c0.n32_adj_3465 ));
    CascadeMux I__11312 (
            .O(N__52399),
            .I(N__52394));
    InMux I__11311 (
            .O(N__52398),
            .I(N__52391));
    InMux I__11310 (
            .O(N__52397),
            .I(N__52388));
    InMux I__11309 (
            .O(N__52394),
            .I(N__52385));
    LocalMux I__11308 (
            .O(N__52391),
            .I(\c0.n33_adj_3315 ));
    LocalMux I__11307 (
            .O(N__52388),
            .I(\c0.n33_adj_3315 ));
    LocalMux I__11306 (
            .O(N__52385),
            .I(\c0.n33_adj_3315 ));
    InMux I__11305 (
            .O(N__52378),
            .I(N__52375));
    LocalMux I__11304 (
            .O(N__52375),
            .I(N__52372));
    Span4Mux_h I__11303 (
            .O(N__52372),
            .I(N__52369));
    Odrv4 I__11302 (
            .O(N__52369),
            .I(\c0.n49_adj_3316 ));
    InMux I__11301 (
            .O(N__52366),
            .I(N__52363));
    LocalMux I__11300 (
            .O(N__52363),
            .I(N__52359));
    InMux I__11299 (
            .O(N__52362),
            .I(N__52356));
    Odrv4 I__11298 (
            .O(N__52359),
            .I(\c0.n35_adj_3317 ));
    LocalMux I__11297 (
            .O(N__52356),
            .I(\c0.n35_adj_3317 ));
    InMux I__11296 (
            .O(N__52351),
            .I(N__52347));
    InMux I__11295 (
            .O(N__52350),
            .I(N__52342));
    LocalMux I__11294 (
            .O(N__52347),
            .I(N__52339));
    InMux I__11293 (
            .O(N__52346),
            .I(N__52335));
    InMux I__11292 (
            .O(N__52345),
            .I(N__52332));
    LocalMux I__11291 (
            .O(N__52342),
            .I(N__52328));
    Span4Mux_h I__11290 (
            .O(N__52339),
            .I(N__52325));
    InMux I__11289 (
            .O(N__52338),
            .I(N__52322));
    LocalMux I__11288 (
            .O(N__52335),
            .I(N__52319));
    LocalMux I__11287 (
            .O(N__52332),
            .I(N__52316));
    CascadeMux I__11286 (
            .O(N__52331),
            .I(N__52313));
    Span4Mux_h I__11285 (
            .O(N__52328),
            .I(N__52308));
    Span4Mux_v I__11284 (
            .O(N__52325),
            .I(N__52308));
    LocalMux I__11283 (
            .O(N__52322),
            .I(N__52305));
    Span4Mux_h I__11282 (
            .O(N__52319),
            .I(N__52300));
    Span4Mux_h I__11281 (
            .O(N__52316),
            .I(N__52300));
    InMux I__11280 (
            .O(N__52313),
            .I(N__52297));
    Span4Mux_v I__11279 (
            .O(N__52308),
            .I(N__52294));
    Span4Mux_h I__11278 (
            .O(N__52305),
            .I(N__52289));
    Span4Mux_v I__11277 (
            .O(N__52300),
            .I(N__52289));
    LocalMux I__11276 (
            .O(N__52297),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__11275 (
            .O(N__52294),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__11274 (
            .O(N__52289),
            .I(\c0.data_in_frame_17_1 ));
    InMux I__11273 (
            .O(N__52282),
            .I(N__52279));
    LocalMux I__11272 (
            .O(N__52279),
            .I(N__52276));
    Span4Mux_v I__11271 (
            .O(N__52276),
            .I(N__52272));
    InMux I__11270 (
            .O(N__52275),
            .I(N__52269));
    Span4Mux_h I__11269 (
            .O(N__52272),
            .I(N__52264));
    LocalMux I__11268 (
            .O(N__52269),
            .I(N__52264));
    Odrv4 I__11267 (
            .O(N__52264),
            .I(\c0.n17871 ));
    InMux I__11266 (
            .O(N__52261),
            .I(N__52258));
    LocalMux I__11265 (
            .O(N__52258),
            .I(N__52255));
    Odrv4 I__11264 (
            .O(N__52255),
            .I(\c0.n22_adj_3363 ));
    CascadeMux I__11263 (
            .O(N__52252),
            .I(\c0.n22_adj_3363_cascade_ ));
    InMux I__11262 (
            .O(N__52249),
            .I(N__52246));
    LocalMux I__11261 (
            .O(N__52246),
            .I(N__52243));
    Odrv4 I__11260 (
            .O(N__52243),
            .I(\c0.n30_adj_3468 ));
    InMux I__11259 (
            .O(N__52240),
            .I(N__52237));
    LocalMux I__11258 (
            .O(N__52237),
            .I(N__52234));
    Odrv12 I__11257 (
            .O(N__52234),
            .I(\c0.n65 ));
    InMux I__11256 (
            .O(N__52231),
            .I(N__52228));
    LocalMux I__11255 (
            .O(N__52228),
            .I(N__52225));
    Sp12to4 I__11254 (
            .O(N__52225),
            .I(N__52222));
    Span12Mux_v I__11253 (
            .O(N__52222),
            .I(N__52219));
    Odrv12 I__11252 (
            .O(N__52219),
            .I(\c0.n19223 ));
    InMux I__11251 (
            .O(N__52216),
            .I(N__52213));
    LocalMux I__11250 (
            .O(N__52213),
            .I(N__52210));
    Span4Mux_h I__11249 (
            .O(N__52210),
            .I(N__52207));
    Span4Mux_v I__11248 (
            .O(N__52207),
            .I(N__52203));
    InMux I__11247 (
            .O(N__52206),
            .I(N__52200));
    Odrv4 I__11246 (
            .O(N__52203),
            .I(\c0.n12218 ));
    LocalMux I__11245 (
            .O(N__52200),
            .I(\c0.n12218 ));
    CascadeMux I__11244 (
            .O(N__52195),
            .I(\c0.n7_adj_3047_cascade_ ));
    CascadeMux I__11243 (
            .O(N__52192),
            .I(\c0.n28_adj_3059_cascade_ ));
    InMux I__11242 (
            .O(N__52189),
            .I(N__52186));
    LocalMux I__11241 (
            .O(N__52186),
            .I(N__52181));
    InMux I__11240 (
            .O(N__52185),
            .I(N__52176));
    InMux I__11239 (
            .O(N__52184),
            .I(N__52176));
    Odrv4 I__11238 (
            .O(N__52181),
            .I(\c0.n36_adj_3452 ));
    LocalMux I__11237 (
            .O(N__52176),
            .I(\c0.n36_adj_3452 ));
    InMux I__11236 (
            .O(N__52171),
            .I(N__52168));
    LocalMux I__11235 (
            .O(N__52168),
            .I(N__52163));
    InMux I__11234 (
            .O(N__52167),
            .I(N__52160));
    InMux I__11233 (
            .O(N__52166),
            .I(N__52155));
    Span4Mux_h I__11232 (
            .O(N__52163),
            .I(N__52152));
    LocalMux I__11231 (
            .O(N__52160),
            .I(N__52149));
    InMux I__11230 (
            .O(N__52159),
            .I(N__52144));
    InMux I__11229 (
            .O(N__52158),
            .I(N__52144));
    LocalMux I__11228 (
            .O(N__52155),
            .I(\c0.n47 ));
    Odrv4 I__11227 (
            .O(N__52152),
            .I(\c0.n47 ));
    Odrv4 I__11226 (
            .O(N__52149),
            .I(\c0.n47 ));
    LocalMux I__11225 (
            .O(N__52144),
            .I(\c0.n47 ));
    InMux I__11224 (
            .O(N__52135),
            .I(N__52131));
    InMux I__11223 (
            .O(N__52134),
            .I(N__52127));
    LocalMux I__11222 (
            .O(N__52131),
            .I(N__52124));
    InMux I__11221 (
            .O(N__52130),
            .I(N__52121));
    LocalMux I__11220 (
            .O(N__52127),
            .I(N__52118));
    Span4Mux_h I__11219 (
            .O(N__52124),
            .I(N__52115));
    LocalMux I__11218 (
            .O(N__52121),
            .I(\c0.n17819 ));
    Odrv4 I__11217 (
            .O(N__52118),
            .I(\c0.n17819 ));
    Odrv4 I__11216 (
            .O(N__52115),
            .I(\c0.n17819 ));
    InMux I__11215 (
            .O(N__52108),
            .I(N__52104));
    InMux I__11214 (
            .O(N__52107),
            .I(N__52100));
    LocalMux I__11213 (
            .O(N__52104),
            .I(N__52097));
    InMux I__11212 (
            .O(N__52103),
            .I(N__52094));
    LocalMux I__11211 (
            .O(N__52100),
            .I(N__52089));
    Span4Mux_h I__11210 (
            .O(N__52097),
            .I(N__52084));
    LocalMux I__11209 (
            .O(N__52094),
            .I(N__52084));
    InMux I__11208 (
            .O(N__52093),
            .I(N__52081));
    InMux I__11207 (
            .O(N__52092),
            .I(N__52078));
    Span4Mux_h I__11206 (
            .O(N__52089),
            .I(N__52075));
    Span4Mux_v I__11205 (
            .O(N__52084),
            .I(N__52070));
    LocalMux I__11204 (
            .O(N__52081),
            .I(N__52070));
    LocalMux I__11203 (
            .O(N__52078),
            .I(N__52067));
    Odrv4 I__11202 (
            .O(N__52075),
            .I(\c0.n20321 ));
    Odrv4 I__11201 (
            .O(N__52070),
            .I(\c0.n20321 ));
    Odrv4 I__11200 (
            .O(N__52067),
            .I(\c0.n20321 ));
    InMux I__11199 (
            .O(N__52060),
            .I(N__52057));
    LocalMux I__11198 (
            .O(N__52057),
            .I(\c0.n19824 ));
    InMux I__11197 (
            .O(N__52054),
            .I(N__52050));
    InMux I__11196 (
            .O(N__52053),
            .I(N__52047));
    LocalMux I__11195 (
            .O(N__52050),
            .I(N__52044));
    LocalMux I__11194 (
            .O(N__52047),
            .I(N__52041));
    Span4Mux_v I__11193 (
            .O(N__52044),
            .I(N__52037));
    Span4Mux_v I__11192 (
            .O(N__52041),
            .I(N__52034));
    InMux I__11191 (
            .O(N__52040),
            .I(N__52031));
    Odrv4 I__11190 (
            .O(N__52037),
            .I(\c0.n12_adj_3469 ));
    Odrv4 I__11189 (
            .O(N__52034),
            .I(\c0.n12_adj_3469 ));
    LocalMux I__11188 (
            .O(N__52031),
            .I(\c0.n12_adj_3469 ));
    CascadeMux I__11187 (
            .O(N__52024),
            .I(\c0.n29_adj_3461_cascade_ ));
    InMux I__11186 (
            .O(N__52021),
            .I(N__52016));
    InMux I__11185 (
            .O(N__52020),
            .I(N__52012));
    InMux I__11184 (
            .O(N__52019),
            .I(N__52009));
    LocalMux I__11183 (
            .O(N__52016),
            .I(N__52006));
    InMux I__11182 (
            .O(N__52015),
            .I(N__52003));
    LocalMux I__11181 (
            .O(N__52012),
            .I(N__52000));
    LocalMux I__11180 (
            .O(N__52009),
            .I(N__51997));
    Span4Mux_v I__11179 (
            .O(N__52006),
            .I(N__51992));
    LocalMux I__11178 (
            .O(N__52003),
            .I(N__51992));
    Span4Mux_v I__11177 (
            .O(N__52000),
            .I(N__51986));
    Span4Mux_v I__11176 (
            .O(N__51997),
            .I(N__51986));
    Span4Mux_h I__11175 (
            .O(N__51992),
            .I(N__51983));
    InMux I__11174 (
            .O(N__51991),
            .I(N__51980));
    Odrv4 I__11173 (
            .O(N__51986),
            .I(\c0.n25_adj_3035 ));
    Odrv4 I__11172 (
            .O(N__51983),
            .I(\c0.n25_adj_3035 ));
    LocalMux I__11171 (
            .O(N__51980),
            .I(\c0.n25_adj_3035 ));
    InMux I__11170 (
            .O(N__51973),
            .I(N__51969));
    InMux I__11169 (
            .O(N__51972),
            .I(N__51966));
    LocalMux I__11168 (
            .O(N__51969),
            .I(N__51963));
    LocalMux I__11167 (
            .O(N__51966),
            .I(N__51960));
    Sp12to4 I__11166 (
            .O(N__51963),
            .I(N__51957));
    Span4Mux_v I__11165 (
            .O(N__51960),
            .I(N__51954));
    Span12Mux_h I__11164 (
            .O(N__51957),
            .I(N__51951));
    Odrv4 I__11163 (
            .O(N__51954),
            .I(\c0.n23_adj_3364 ));
    Odrv12 I__11162 (
            .O(N__51951),
            .I(\c0.n23_adj_3364 ));
    InMux I__11161 (
            .O(N__51946),
            .I(N__51943));
    LocalMux I__11160 (
            .O(N__51943),
            .I(N__51939));
    InMux I__11159 (
            .O(N__51942),
            .I(N__51936));
    Span4Mux_v I__11158 (
            .O(N__51939),
            .I(N__51933));
    LocalMux I__11157 (
            .O(N__51936),
            .I(N__51930));
    Span4Mux_h I__11156 (
            .O(N__51933),
            .I(N__51927));
    Span4Mux_v I__11155 (
            .O(N__51930),
            .I(N__51924));
    Odrv4 I__11154 (
            .O(N__51927),
            .I(\c0.n24_adj_3335 ));
    Odrv4 I__11153 (
            .O(N__51924),
            .I(\c0.n24_adj_3335 ));
    CascadeMux I__11152 (
            .O(N__51919),
            .I(\c0.n36_adj_3470_cascade_ ));
    InMux I__11151 (
            .O(N__51916),
            .I(N__51913));
    LocalMux I__11150 (
            .O(N__51913),
            .I(N__51909));
    InMux I__11149 (
            .O(N__51912),
            .I(N__51906));
    Span4Mux_v I__11148 (
            .O(N__51909),
            .I(N__51903));
    LocalMux I__11147 (
            .O(N__51906),
            .I(N__51900));
    Odrv4 I__11146 (
            .O(N__51903),
            .I(\c0.n22_adj_3341 ));
    Odrv4 I__11145 (
            .O(N__51900),
            .I(\c0.n22_adj_3341 ));
    CascadeMux I__11144 (
            .O(N__51895),
            .I(\c0.n11_adj_3124_cascade_ ));
    InMux I__11143 (
            .O(N__51892),
            .I(N__51889));
    LocalMux I__11142 (
            .O(N__51889),
            .I(N__51886));
    Span4Mux_h I__11141 (
            .O(N__51886),
            .I(N__51882));
    InMux I__11140 (
            .O(N__51885),
            .I(N__51879));
    Odrv4 I__11139 (
            .O(N__51882),
            .I(\c0.n22_adj_3287 ));
    LocalMux I__11138 (
            .O(N__51879),
            .I(\c0.n22_adj_3287 ));
    CascadeMux I__11137 (
            .O(N__51874),
            .I(\c0.n47_adj_3286_cascade_ ));
    InMux I__11136 (
            .O(N__51871),
            .I(N__51868));
    LocalMux I__11135 (
            .O(N__51868),
            .I(\c0.n51_adj_3290 ));
    CascadeMux I__11134 (
            .O(N__51865),
            .I(\c0.n52_adj_3288_cascade_ ));
    InMux I__11133 (
            .O(N__51862),
            .I(N__51859));
    LocalMux I__11132 (
            .O(N__51859),
            .I(N__51856));
    Span4Mux_h I__11131 (
            .O(N__51856),
            .I(N__51853));
    Span4Mux_v I__11130 (
            .O(N__51853),
            .I(N__51850));
    Odrv4 I__11129 (
            .O(N__51850),
            .I(\c0.n6_adj_3291 ));
    CascadeMux I__11128 (
            .O(N__51847),
            .I(N__51843));
    CascadeMux I__11127 (
            .O(N__51846),
            .I(N__51840));
    InMux I__11126 (
            .O(N__51843),
            .I(N__51837));
    InMux I__11125 (
            .O(N__51840),
            .I(N__51834));
    LocalMux I__11124 (
            .O(N__51837),
            .I(N__51830));
    LocalMux I__11123 (
            .O(N__51834),
            .I(N__51827));
    InMux I__11122 (
            .O(N__51833),
            .I(N__51824));
    Span4Mux_h I__11121 (
            .O(N__51830),
            .I(N__51821));
    Span4Mux_h I__11120 (
            .O(N__51827),
            .I(N__51818));
    LocalMux I__11119 (
            .O(N__51824),
            .I(\c0.data_in_frame_11_6 ));
    Odrv4 I__11118 (
            .O(N__51821),
            .I(\c0.data_in_frame_11_6 ));
    Odrv4 I__11117 (
            .O(N__51818),
            .I(\c0.data_in_frame_11_6 ));
    CascadeMux I__11116 (
            .O(N__51811),
            .I(\c0.n19909_cascade_ ));
    InMux I__11115 (
            .O(N__51808),
            .I(N__51804));
    InMux I__11114 (
            .O(N__51807),
            .I(N__51801));
    LocalMux I__11113 (
            .O(N__51804),
            .I(N__51798));
    LocalMux I__11112 (
            .O(N__51801),
            .I(N__51795));
    Span4Mux_h I__11111 (
            .O(N__51798),
            .I(N__51792));
    Odrv4 I__11110 (
            .O(N__51795),
            .I(\c0.n87 ));
    Odrv4 I__11109 (
            .O(N__51792),
            .I(\c0.n87 ));
    InMux I__11108 (
            .O(N__51787),
            .I(N__51782));
    InMux I__11107 (
            .O(N__51786),
            .I(N__51777));
    InMux I__11106 (
            .O(N__51785),
            .I(N__51777));
    LocalMux I__11105 (
            .O(N__51782),
            .I(N__51770));
    LocalMux I__11104 (
            .O(N__51777),
            .I(N__51770));
    InMux I__11103 (
            .O(N__51776),
            .I(N__51765));
    InMux I__11102 (
            .O(N__51775),
            .I(N__51765));
    Odrv12 I__11101 (
            .O(N__51770),
            .I(\c0.n6_adj_3137 ));
    LocalMux I__11100 (
            .O(N__51765),
            .I(\c0.n6_adj_3137 ));
    InMux I__11099 (
            .O(N__51760),
            .I(N__51756));
    CascadeMux I__11098 (
            .O(N__51759),
            .I(N__51753));
    LocalMux I__11097 (
            .O(N__51756),
            .I(N__51750));
    InMux I__11096 (
            .O(N__51753),
            .I(N__51747));
    Span4Mux_v I__11095 (
            .O(N__51750),
            .I(N__51744));
    LocalMux I__11094 (
            .O(N__51747),
            .I(N__51741));
    Span4Mux_h I__11093 (
            .O(N__51744),
            .I(N__51736));
    Span4Mux_h I__11092 (
            .O(N__51741),
            .I(N__51736));
    Span4Mux_v I__11091 (
            .O(N__51736),
            .I(N__51733));
    Odrv4 I__11090 (
            .O(N__51733),
            .I(\c0.n35_adj_3098 ));
    InMux I__11089 (
            .O(N__51730),
            .I(N__51726));
    InMux I__11088 (
            .O(N__51729),
            .I(N__51723));
    LocalMux I__11087 (
            .O(N__51726),
            .I(\c0.n19909 ));
    LocalMux I__11086 (
            .O(N__51723),
            .I(\c0.n19909 ));
    CascadeMux I__11085 (
            .O(N__51718),
            .I(N__51715));
    InMux I__11084 (
            .O(N__51715),
            .I(N__51712));
    LocalMux I__11083 (
            .O(N__51712),
            .I(N__51708));
    InMux I__11082 (
            .O(N__51711),
            .I(N__51703));
    Span4Mux_h I__11081 (
            .O(N__51708),
            .I(N__51700));
    InMux I__11080 (
            .O(N__51707),
            .I(N__51695));
    InMux I__11079 (
            .O(N__51706),
            .I(N__51695));
    LocalMux I__11078 (
            .O(N__51703),
            .I(\c0.data_in_frame_13_5 ));
    Odrv4 I__11077 (
            .O(N__51700),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__11076 (
            .O(N__51695),
            .I(\c0.data_in_frame_13_5 ));
    InMux I__11075 (
            .O(N__51688),
            .I(N__51682));
    InMux I__11074 (
            .O(N__51687),
            .I(N__51675));
    InMux I__11073 (
            .O(N__51686),
            .I(N__51675));
    InMux I__11072 (
            .O(N__51685),
            .I(N__51675));
    LocalMux I__11071 (
            .O(N__51682),
            .I(N__51669));
    LocalMux I__11070 (
            .O(N__51675),
            .I(N__51666));
    InMux I__11069 (
            .O(N__51674),
            .I(N__51663));
    InMux I__11068 (
            .O(N__51673),
            .I(N__51658));
    InMux I__11067 (
            .O(N__51672),
            .I(N__51658));
    Odrv4 I__11066 (
            .O(N__51669),
            .I(\c0.n20826 ));
    Odrv4 I__11065 (
            .O(N__51666),
            .I(\c0.n20826 ));
    LocalMux I__11064 (
            .O(N__51663),
            .I(\c0.n20826 ));
    LocalMux I__11063 (
            .O(N__51658),
            .I(\c0.n20826 ));
    InMux I__11062 (
            .O(N__51649),
            .I(N__51646));
    LocalMux I__11061 (
            .O(N__51646),
            .I(N__51643));
    Odrv12 I__11060 (
            .O(N__51643),
            .I(\c0.n54_adj_3234 ));
    CascadeMux I__11059 (
            .O(N__51640),
            .I(\c0.n43_adj_3232_cascade_ ));
    InMux I__11058 (
            .O(N__51637),
            .I(N__51633));
    InMux I__11057 (
            .O(N__51636),
            .I(N__51630));
    LocalMux I__11056 (
            .O(N__51633),
            .I(N__51627));
    LocalMux I__11055 (
            .O(N__51630),
            .I(N__51624));
    Span4Mux_v I__11054 (
            .O(N__51627),
            .I(N__51618));
    Span4Mux_h I__11053 (
            .O(N__51624),
            .I(N__51618));
    InMux I__11052 (
            .O(N__51623),
            .I(N__51614));
    Span4Mux_h I__11051 (
            .O(N__51618),
            .I(N__51611));
    InMux I__11050 (
            .O(N__51617),
            .I(N__51608));
    LocalMux I__11049 (
            .O(N__51614),
            .I(\c0.n17849 ));
    Odrv4 I__11048 (
            .O(N__51611),
            .I(\c0.n17849 ));
    LocalMux I__11047 (
            .O(N__51608),
            .I(\c0.n17849 ));
    InMux I__11046 (
            .O(N__51601),
            .I(N__51598));
    LocalMux I__11045 (
            .O(N__51598),
            .I(\c0.n49_adj_3237 ));
    CascadeMux I__11044 (
            .O(N__51595),
            .I(\c0.n7_adj_3225_cascade_ ));
    CascadeMux I__11043 (
            .O(N__51592),
            .I(N__51589));
    InMux I__11042 (
            .O(N__51589),
            .I(N__51583));
    InMux I__11041 (
            .O(N__51588),
            .I(N__51583));
    LocalMux I__11040 (
            .O(N__51583),
            .I(N__51579));
    CascadeMux I__11039 (
            .O(N__51582),
            .I(N__51576));
    Span4Mux_h I__11038 (
            .O(N__51579),
            .I(N__51573));
    InMux I__11037 (
            .O(N__51576),
            .I(N__51570));
    Span4Mux_h I__11036 (
            .O(N__51573),
            .I(N__51567));
    LocalMux I__11035 (
            .O(N__51570),
            .I(N__51562));
    Span4Mux_v I__11034 (
            .O(N__51567),
            .I(N__51562));
    Odrv4 I__11033 (
            .O(N__51562),
            .I(\c0.data_in_frame_15_4 ));
    InMux I__11032 (
            .O(N__51559),
            .I(N__51556));
    LocalMux I__11031 (
            .O(N__51556),
            .I(\c0.n7_adj_3225 ));
    InMux I__11030 (
            .O(N__51553),
            .I(N__51550));
    LocalMux I__11029 (
            .O(N__51550),
            .I(N__51547));
    Odrv4 I__11028 (
            .O(N__51547),
            .I(\c0.n44_adj_3226 ));
    InMux I__11027 (
            .O(N__51544),
            .I(N__51541));
    LocalMux I__11026 (
            .O(N__51541),
            .I(N__51535));
    InMux I__11025 (
            .O(N__51540),
            .I(N__51532));
    InMux I__11024 (
            .O(N__51539),
            .I(N__51527));
    InMux I__11023 (
            .O(N__51538),
            .I(N__51527));
    Odrv12 I__11022 (
            .O(N__51535),
            .I(\c0.data_in_frame_10_4 ));
    LocalMux I__11021 (
            .O(N__51532),
            .I(\c0.data_in_frame_10_4 ));
    LocalMux I__11020 (
            .O(N__51527),
            .I(\c0.data_in_frame_10_4 ));
    CascadeMux I__11019 (
            .O(N__51520),
            .I(N__51515));
    CascadeMux I__11018 (
            .O(N__51519),
            .I(N__51510));
    CascadeMux I__11017 (
            .O(N__51518),
            .I(N__51507));
    InMux I__11016 (
            .O(N__51515),
            .I(N__51504));
    InMux I__11015 (
            .O(N__51514),
            .I(N__51501));
    InMux I__11014 (
            .O(N__51513),
            .I(N__51498));
    InMux I__11013 (
            .O(N__51510),
            .I(N__51495));
    InMux I__11012 (
            .O(N__51507),
            .I(N__51492));
    LocalMux I__11011 (
            .O(N__51504),
            .I(N__51489));
    LocalMux I__11010 (
            .O(N__51501),
            .I(N__51484));
    LocalMux I__11009 (
            .O(N__51498),
            .I(N__51484));
    LocalMux I__11008 (
            .O(N__51495),
            .I(N__51479));
    LocalMux I__11007 (
            .O(N__51492),
            .I(N__51479));
    Span4Mux_v I__11006 (
            .O(N__51489),
            .I(N__51475));
    Span4Mux_v I__11005 (
            .O(N__51484),
            .I(N__51472));
    Span4Mux_v I__11004 (
            .O(N__51479),
            .I(N__51469));
    InMux I__11003 (
            .O(N__51478),
            .I(N__51466));
    Odrv4 I__11002 (
            .O(N__51475),
            .I(\c0.data_in_frame_8_1 ));
    Odrv4 I__11001 (
            .O(N__51472),
            .I(\c0.data_in_frame_8_1 ));
    Odrv4 I__11000 (
            .O(N__51469),
            .I(\c0.data_in_frame_8_1 ));
    LocalMux I__10999 (
            .O(N__51466),
            .I(\c0.data_in_frame_8_1 ));
    CascadeMux I__10998 (
            .O(N__51457),
            .I(N__51453));
    CascadeMux I__10997 (
            .O(N__51456),
            .I(N__51450));
    InMux I__10996 (
            .O(N__51453),
            .I(N__51445));
    InMux I__10995 (
            .O(N__51450),
            .I(N__51445));
    LocalMux I__10994 (
            .O(N__51445),
            .I(N__51442));
    Span4Mux_h I__10993 (
            .O(N__51442),
            .I(N__51439));
    Odrv4 I__10992 (
            .O(N__51439),
            .I(\c0.n41_adj_3365 ));
    InMux I__10991 (
            .O(N__51436),
            .I(N__51433));
    LocalMux I__10990 (
            .O(N__51433),
            .I(N__51429));
    InMux I__10989 (
            .O(N__51432),
            .I(N__51426));
    Odrv4 I__10988 (
            .O(N__51429),
            .I(\c0.n16_adj_3218 ));
    LocalMux I__10987 (
            .O(N__51426),
            .I(\c0.n16_adj_3218 ));
    InMux I__10986 (
            .O(N__51421),
            .I(N__51418));
    LocalMux I__10985 (
            .O(N__51418),
            .I(\c0.n48 ));
    InMux I__10984 (
            .O(N__51415),
            .I(N__51411));
    CascadeMux I__10983 (
            .O(N__51414),
            .I(N__51407));
    LocalMux I__10982 (
            .O(N__51411),
            .I(N__51403));
    InMux I__10981 (
            .O(N__51410),
            .I(N__51400));
    InMux I__10980 (
            .O(N__51407),
            .I(N__51396));
    CascadeMux I__10979 (
            .O(N__51406),
            .I(N__51393));
    Span4Mux_v I__10978 (
            .O(N__51403),
            .I(N__51390));
    LocalMux I__10977 (
            .O(N__51400),
            .I(N__51387));
    InMux I__10976 (
            .O(N__51399),
            .I(N__51383));
    LocalMux I__10975 (
            .O(N__51396),
            .I(N__51380));
    InMux I__10974 (
            .O(N__51393),
            .I(N__51377));
    Span4Mux_h I__10973 (
            .O(N__51390),
            .I(N__51374));
    Span12Mux_s10_v I__10972 (
            .O(N__51387),
            .I(N__51371));
    InMux I__10971 (
            .O(N__51386),
            .I(N__51368));
    LocalMux I__10970 (
            .O(N__51383),
            .I(N__51365));
    Span4Mux_h I__10969 (
            .O(N__51380),
            .I(N__51362));
    LocalMux I__10968 (
            .O(N__51377),
            .I(\c0.data_in_frame_5_1 ));
    Odrv4 I__10967 (
            .O(N__51374),
            .I(\c0.data_in_frame_5_1 ));
    Odrv12 I__10966 (
            .O(N__51371),
            .I(\c0.data_in_frame_5_1 ));
    LocalMux I__10965 (
            .O(N__51368),
            .I(\c0.data_in_frame_5_1 ));
    Odrv4 I__10964 (
            .O(N__51365),
            .I(\c0.data_in_frame_5_1 ));
    Odrv4 I__10963 (
            .O(N__51362),
            .I(\c0.data_in_frame_5_1 ));
    InMux I__10962 (
            .O(N__51349),
            .I(N__51346));
    LocalMux I__10961 (
            .O(N__51346),
            .I(N__51342));
    InMux I__10960 (
            .O(N__51345),
            .I(N__51339));
    Span4Mux_v I__10959 (
            .O(N__51342),
            .I(N__51335));
    LocalMux I__10958 (
            .O(N__51339),
            .I(N__51332));
    InMux I__10957 (
            .O(N__51338),
            .I(N__51327));
    Span4Mux_v I__10956 (
            .O(N__51335),
            .I(N__51324));
    Span4Mux_v I__10955 (
            .O(N__51332),
            .I(N__51321));
    InMux I__10954 (
            .O(N__51331),
            .I(N__51318));
    InMux I__10953 (
            .O(N__51330),
            .I(N__51315));
    LocalMux I__10952 (
            .O(N__51327),
            .I(N__51312));
    Odrv4 I__10951 (
            .O(N__51324),
            .I(\c0.n20224 ));
    Odrv4 I__10950 (
            .O(N__51321),
            .I(\c0.n20224 ));
    LocalMux I__10949 (
            .O(N__51318),
            .I(\c0.n20224 ));
    LocalMux I__10948 (
            .O(N__51315),
            .I(\c0.n20224 ));
    Odrv12 I__10947 (
            .O(N__51312),
            .I(\c0.n20224 ));
    CascadeMux I__10946 (
            .O(N__51301),
            .I(N__51298));
    InMux I__10945 (
            .O(N__51298),
            .I(N__51295));
    LocalMux I__10944 (
            .O(N__51295),
            .I(\c0.n5_adj_3549 ));
    InMux I__10943 (
            .O(N__51292),
            .I(N__51288));
    InMux I__10942 (
            .O(N__51291),
            .I(N__51284));
    LocalMux I__10941 (
            .O(N__51288),
            .I(N__51279));
    InMux I__10940 (
            .O(N__51287),
            .I(N__51276));
    LocalMux I__10939 (
            .O(N__51284),
            .I(N__51273));
    InMux I__10938 (
            .O(N__51283),
            .I(N__51270));
    CascadeMux I__10937 (
            .O(N__51282),
            .I(N__51267));
    Span4Mux_v I__10936 (
            .O(N__51279),
            .I(N__51261));
    LocalMux I__10935 (
            .O(N__51276),
            .I(N__51261));
    Span4Mux_h I__10934 (
            .O(N__51273),
            .I(N__51252));
    LocalMux I__10933 (
            .O(N__51270),
            .I(N__51249));
    InMux I__10932 (
            .O(N__51267),
            .I(N__51244));
    InMux I__10931 (
            .O(N__51266),
            .I(N__51244));
    Span4Mux_h I__10930 (
            .O(N__51261),
            .I(N__51241));
    InMux I__10929 (
            .O(N__51260),
            .I(N__51234));
    InMux I__10928 (
            .O(N__51259),
            .I(N__51234));
    InMux I__10927 (
            .O(N__51258),
            .I(N__51234));
    InMux I__10926 (
            .O(N__51257),
            .I(N__51227));
    InMux I__10925 (
            .O(N__51256),
            .I(N__51227));
    InMux I__10924 (
            .O(N__51255),
            .I(N__51227));
    Odrv4 I__10923 (
            .O(N__51252),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__10922 (
            .O(N__51249),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__10921 (
            .O(N__51244),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__10920 (
            .O(N__51241),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__10919 (
            .O(N__51234),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__10918 (
            .O(N__51227),
            .I(\c0.data_in_frame_4_7 ));
    InMux I__10917 (
            .O(N__51214),
            .I(N__51211));
    LocalMux I__10916 (
            .O(N__51211),
            .I(\c0.n11613 ));
    InMux I__10915 (
            .O(N__51208),
            .I(N__51204));
    InMux I__10914 (
            .O(N__51207),
            .I(N__51201));
    LocalMux I__10913 (
            .O(N__51204),
            .I(N__51197));
    LocalMux I__10912 (
            .O(N__51201),
            .I(N__51194));
    InMux I__10911 (
            .O(N__51200),
            .I(N__51191));
    Span4Mux_h I__10910 (
            .O(N__51197),
            .I(N__51188));
    Span4Mux_h I__10909 (
            .O(N__51194),
            .I(N__51185));
    LocalMux I__10908 (
            .O(N__51191),
            .I(\c0.data_in_frame_17_6 ));
    Odrv4 I__10907 (
            .O(N__51188),
            .I(\c0.data_in_frame_17_6 ));
    Odrv4 I__10906 (
            .O(N__51185),
            .I(\c0.data_in_frame_17_6 ));
    InMux I__10905 (
            .O(N__51178),
            .I(N__51175));
    LocalMux I__10904 (
            .O(N__51175),
            .I(N__51172));
    Span4Mux_v I__10903 (
            .O(N__51172),
            .I(N__51168));
    InMux I__10902 (
            .O(N__51171),
            .I(N__51165));
    Span4Mux_h I__10901 (
            .O(N__51168),
            .I(N__51162));
    LocalMux I__10900 (
            .O(N__51165),
            .I(data_in_frame_18_0));
    Odrv4 I__10899 (
            .O(N__51162),
            .I(data_in_frame_18_0));
    CascadeMux I__10898 (
            .O(N__51157),
            .I(\c0.n11613_cascade_ ));
    InMux I__10897 (
            .O(N__51154),
            .I(N__51150));
    InMux I__10896 (
            .O(N__51153),
            .I(N__51147));
    LocalMux I__10895 (
            .O(N__51150),
            .I(N__51142));
    LocalMux I__10894 (
            .O(N__51147),
            .I(N__51142));
    Odrv4 I__10893 (
            .O(N__51142),
            .I(\c0.n19477 ));
    InMux I__10892 (
            .O(N__51139),
            .I(N__51136));
    LocalMux I__10891 (
            .O(N__51136),
            .I(\c0.n17_adj_3482 ));
    InMux I__10890 (
            .O(N__51133),
            .I(N__51130));
    LocalMux I__10889 (
            .O(N__51130),
            .I(N__51126));
    CascadeMux I__10888 (
            .O(N__51129),
            .I(N__51123));
    Span4Mux_h I__10887 (
            .O(N__51126),
            .I(N__51119));
    InMux I__10886 (
            .O(N__51123),
            .I(N__51114));
    InMux I__10885 (
            .O(N__51122),
            .I(N__51114));
    Odrv4 I__10884 (
            .O(N__51119),
            .I(\c0.data_in_frame_13_6 ));
    LocalMux I__10883 (
            .O(N__51114),
            .I(\c0.data_in_frame_13_6 ));
    InMux I__10882 (
            .O(N__51109),
            .I(N__51105));
    InMux I__10881 (
            .O(N__51108),
            .I(N__51101));
    LocalMux I__10880 (
            .O(N__51105),
            .I(N__51098));
    CascadeMux I__10879 (
            .O(N__51104),
            .I(N__51094));
    LocalMux I__10878 (
            .O(N__51101),
            .I(N__51091));
    Span4Mux_v I__10877 (
            .O(N__51098),
            .I(N__51087));
    InMux I__10876 (
            .O(N__51097),
            .I(N__51084));
    InMux I__10875 (
            .O(N__51094),
            .I(N__51081));
    Span4Mux_h I__10874 (
            .O(N__51091),
            .I(N__51078));
    InMux I__10873 (
            .O(N__51090),
            .I(N__51075));
    Span4Mux_h I__10872 (
            .O(N__51087),
            .I(N__51070));
    LocalMux I__10871 (
            .O(N__51084),
            .I(N__51070));
    LocalMux I__10870 (
            .O(N__51081),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__10869 (
            .O(N__51078),
            .I(\c0.data_in_frame_7_4 ));
    LocalMux I__10868 (
            .O(N__51075),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__10867 (
            .O(N__51070),
            .I(\c0.data_in_frame_7_4 ));
    InMux I__10866 (
            .O(N__51061),
            .I(N__51058));
    LocalMux I__10865 (
            .O(N__51058),
            .I(N__51055));
    Span4Mux_v I__10864 (
            .O(N__51055),
            .I(N__51051));
    InMux I__10863 (
            .O(N__51054),
            .I(N__51048));
    Odrv4 I__10862 (
            .O(N__51051),
            .I(\c0.n20391 ));
    LocalMux I__10861 (
            .O(N__51048),
            .I(\c0.n20391 ));
    InMux I__10860 (
            .O(N__51043),
            .I(N__51040));
    LocalMux I__10859 (
            .O(N__51040),
            .I(\c0.n4 ));
    InMux I__10858 (
            .O(N__51037),
            .I(N__51034));
    LocalMux I__10857 (
            .O(N__51034),
            .I(N__51030));
    InMux I__10856 (
            .O(N__51033),
            .I(N__51027));
    Span4Mux_v I__10855 (
            .O(N__51030),
            .I(N__51022));
    LocalMux I__10854 (
            .O(N__51027),
            .I(N__51022));
    Span4Mux_h I__10853 (
            .O(N__51022),
            .I(N__51019));
    Odrv4 I__10852 (
            .O(N__51019),
            .I(\c0.n12026 ));
    InMux I__10851 (
            .O(N__51016),
            .I(N__51012));
    InMux I__10850 (
            .O(N__51015),
            .I(N__51009));
    LocalMux I__10849 (
            .O(N__51012),
            .I(N__51006));
    LocalMux I__10848 (
            .O(N__51009),
            .I(N__51003));
    Span4Mux_v I__10847 (
            .O(N__51006),
            .I(N__51000));
    Span4Mux_v I__10846 (
            .O(N__51003),
            .I(N__50997));
    Odrv4 I__10845 (
            .O(N__51000),
            .I(\c0.n5 ));
    Odrv4 I__10844 (
            .O(N__50997),
            .I(\c0.n5 ));
    CascadeMux I__10843 (
            .O(N__50992),
            .I(\c0.n4_cascade_ ));
    InMux I__10842 (
            .O(N__50989),
            .I(N__50985));
    InMux I__10841 (
            .O(N__50988),
            .I(N__50981));
    LocalMux I__10840 (
            .O(N__50985),
            .I(N__50978));
    CascadeMux I__10839 (
            .O(N__50984),
            .I(N__50974));
    LocalMux I__10838 (
            .O(N__50981),
            .I(N__50971));
    Span4Mux_h I__10837 (
            .O(N__50978),
            .I(N__50968));
    InMux I__10836 (
            .O(N__50977),
            .I(N__50965));
    InMux I__10835 (
            .O(N__50974),
            .I(N__50962));
    Span4Mux_h I__10834 (
            .O(N__50971),
            .I(N__50959));
    Span4Mux_v I__10833 (
            .O(N__50968),
            .I(N__50956));
    LocalMux I__10832 (
            .O(N__50965),
            .I(N__50953));
    LocalMux I__10831 (
            .O(N__50962),
            .I(\c0.data_in_frame_11_4 ));
    Odrv4 I__10830 (
            .O(N__50959),
            .I(\c0.data_in_frame_11_4 ));
    Odrv4 I__10829 (
            .O(N__50956),
            .I(\c0.data_in_frame_11_4 ));
    Odrv12 I__10828 (
            .O(N__50953),
            .I(\c0.data_in_frame_11_4 ));
    CascadeMux I__10827 (
            .O(N__50944),
            .I(N__50941));
    InMux I__10826 (
            .O(N__50941),
            .I(N__50938));
    LocalMux I__10825 (
            .O(N__50938),
            .I(N__50934));
    CascadeMux I__10824 (
            .O(N__50937),
            .I(N__50930));
    Span4Mux_v I__10823 (
            .O(N__50934),
            .I(N__50927));
    InMux I__10822 (
            .O(N__50933),
            .I(N__50924));
    InMux I__10821 (
            .O(N__50930),
            .I(N__50921));
    Span4Mux_h I__10820 (
            .O(N__50927),
            .I(N__50918));
    LocalMux I__10819 (
            .O(N__50924),
            .I(N__50915));
    LocalMux I__10818 (
            .O(N__50921),
            .I(\c0.data_in_frame_10_0 ));
    Odrv4 I__10817 (
            .O(N__50918),
            .I(\c0.data_in_frame_10_0 ));
    Odrv4 I__10816 (
            .O(N__50915),
            .I(\c0.data_in_frame_10_0 ));
    InMux I__10815 (
            .O(N__50908),
            .I(N__50905));
    LocalMux I__10814 (
            .O(N__50905),
            .I(N__50900));
    InMux I__10813 (
            .O(N__50904),
            .I(N__50897));
    CascadeMux I__10812 (
            .O(N__50903),
            .I(N__50894));
    Span4Mux_v I__10811 (
            .O(N__50900),
            .I(N__50891));
    LocalMux I__10810 (
            .O(N__50897),
            .I(N__50888));
    InMux I__10809 (
            .O(N__50894),
            .I(N__50885));
    Span4Mux_h I__10808 (
            .O(N__50891),
            .I(N__50882));
    Span4Mux_h I__10807 (
            .O(N__50888),
            .I(N__50879));
    LocalMux I__10806 (
            .O(N__50885),
            .I(\c0.data_in_frame_21_0 ));
    Odrv4 I__10805 (
            .O(N__50882),
            .I(\c0.data_in_frame_21_0 ));
    Odrv4 I__10804 (
            .O(N__50879),
            .I(\c0.data_in_frame_21_0 ));
    CascadeMux I__10803 (
            .O(N__50872),
            .I(\c0.n36_adj_3212_cascade_ ));
    InMux I__10802 (
            .O(N__50869),
            .I(N__50866));
    LocalMux I__10801 (
            .O(N__50866),
            .I(\c0.n41_adj_3213 ));
    InMux I__10800 (
            .O(N__50863),
            .I(N__50860));
    LocalMux I__10799 (
            .O(N__50860),
            .I(N__50857));
    Span4Mux_v I__10798 (
            .O(N__50857),
            .I(N__50854));
    Span4Mux_h I__10797 (
            .O(N__50854),
            .I(N__50849));
    InMux I__10796 (
            .O(N__50853),
            .I(N__50844));
    InMux I__10795 (
            .O(N__50852),
            .I(N__50844));
    Odrv4 I__10794 (
            .O(N__50849),
            .I(\c0.n20340 ));
    LocalMux I__10793 (
            .O(N__50844),
            .I(\c0.n20340 ));
    CascadeMux I__10792 (
            .O(N__50839),
            .I(\c0.n11651_cascade_ ));
    InMux I__10791 (
            .O(N__50836),
            .I(N__50833));
    LocalMux I__10790 (
            .O(N__50833),
            .I(\c0.n27_adj_3082 ));
    InMux I__10789 (
            .O(N__50830),
            .I(N__50826));
    InMux I__10788 (
            .O(N__50829),
            .I(N__50823));
    LocalMux I__10787 (
            .O(N__50826),
            .I(N__50819));
    LocalMux I__10786 (
            .O(N__50823),
            .I(N__50816));
    InMux I__10785 (
            .O(N__50822),
            .I(N__50813));
    Span4Mux_h I__10784 (
            .O(N__50819),
            .I(N__50810));
    Span4Mux_h I__10783 (
            .O(N__50816),
            .I(N__50807));
    LocalMux I__10782 (
            .O(N__50813),
            .I(N__50804));
    Odrv4 I__10781 (
            .O(N__50810),
            .I(\c0.n11800 ));
    Odrv4 I__10780 (
            .O(N__50807),
            .I(\c0.n11800 ));
    Odrv4 I__10779 (
            .O(N__50804),
            .I(\c0.n11800 ));
    InMux I__10778 (
            .O(N__50797),
            .I(N__50793));
    InMux I__10777 (
            .O(N__50796),
            .I(N__50790));
    LocalMux I__10776 (
            .O(N__50793),
            .I(\c0.n31 ));
    LocalMux I__10775 (
            .O(N__50790),
            .I(\c0.n31 ));
    CascadeMux I__10774 (
            .O(N__50785),
            .I(N__50781));
    CascadeMux I__10773 (
            .O(N__50784),
            .I(N__50778));
    InMux I__10772 (
            .O(N__50781),
            .I(N__50775));
    InMux I__10771 (
            .O(N__50778),
            .I(N__50772));
    LocalMux I__10770 (
            .O(N__50775),
            .I(N__50769));
    LocalMux I__10769 (
            .O(N__50772),
            .I(N__50766));
    Span4Mux_v I__10768 (
            .O(N__50769),
            .I(N__50763));
    Span4Mux_v I__10767 (
            .O(N__50766),
            .I(N__50760));
    Span4Mux_h I__10766 (
            .O(N__50763),
            .I(N__50757));
    Span4Mux_h I__10765 (
            .O(N__50760),
            .I(N__50754));
    Odrv4 I__10764 (
            .O(N__50757),
            .I(\c0.n37_adj_3153 ));
    Odrv4 I__10763 (
            .O(N__50754),
            .I(\c0.n37_adj_3153 ));
    InMux I__10762 (
            .O(N__50749),
            .I(N__50746));
    LocalMux I__10761 (
            .O(N__50746),
            .I(N__50743));
    Odrv12 I__10760 (
            .O(N__50743),
            .I(\c0.n35_adj_3233 ));
    InMux I__10759 (
            .O(N__50740),
            .I(N__50736));
    InMux I__10758 (
            .O(N__50739),
            .I(N__50733));
    LocalMux I__10757 (
            .O(N__50736),
            .I(N__50730));
    LocalMux I__10756 (
            .O(N__50733),
            .I(N__50727));
    Span4Mux_h I__10755 (
            .O(N__50730),
            .I(N__50722));
    Span4Mux_v I__10754 (
            .O(N__50727),
            .I(N__50722));
    Span4Mux_v I__10753 (
            .O(N__50722),
            .I(N__50719));
    Odrv4 I__10752 (
            .O(N__50719),
            .I(\c0.n60 ));
    CascadeMux I__10751 (
            .O(N__50716),
            .I(\c0.n52_adj_3223_cascade_ ));
    CascadeMux I__10750 (
            .O(N__50713),
            .I(N__50710));
    InMux I__10749 (
            .O(N__50710),
            .I(N__50707));
    LocalMux I__10748 (
            .O(N__50707),
            .I(N__50704));
    Span4Mux_h I__10747 (
            .O(N__50704),
            .I(N__50701));
    Odrv4 I__10746 (
            .O(N__50701),
            .I(\c0.n60_adj_3503 ));
    InMux I__10745 (
            .O(N__50698),
            .I(N__50695));
    LocalMux I__10744 (
            .O(N__50695),
            .I(N__50692));
    Span4Mux_h I__10743 (
            .O(N__50692),
            .I(N__50688));
    InMux I__10742 (
            .O(N__50691),
            .I(N__50685));
    Odrv4 I__10741 (
            .O(N__50688),
            .I(\c0.n52_adj_3402 ));
    LocalMux I__10740 (
            .O(N__50685),
            .I(\c0.n52_adj_3402 ));
    CascadeMux I__10739 (
            .O(N__50680),
            .I(N__50675));
    CascadeMux I__10738 (
            .O(N__50679),
            .I(N__50669));
    InMux I__10737 (
            .O(N__50678),
            .I(N__50666));
    InMux I__10736 (
            .O(N__50675),
            .I(N__50663));
    InMux I__10735 (
            .O(N__50674),
            .I(N__50660));
    InMux I__10734 (
            .O(N__50673),
            .I(N__50654));
    InMux I__10733 (
            .O(N__50672),
            .I(N__50654));
    InMux I__10732 (
            .O(N__50669),
            .I(N__50651));
    LocalMux I__10731 (
            .O(N__50666),
            .I(N__50648));
    LocalMux I__10730 (
            .O(N__50663),
            .I(N__50645));
    LocalMux I__10729 (
            .O(N__50660),
            .I(N__50642));
    InMux I__10728 (
            .O(N__50659),
            .I(N__50636));
    LocalMux I__10727 (
            .O(N__50654),
            .I(N__50633));
    LocalMux I__10726 (
            .O(N__50651),
            .I(N__50624));
    Span4Mux_v I__10725 (
            .O(N__50648),
            .I(N__50624));
    Span4Mux_v I__10724 (
            .O(N__50645),
            .I(N__50624));
    Span4Mux_h I__10723 (
            .O(N__50642),
            .I(N__50624));
    InMux I__10722 (
            .O(N__50641),
            .I(N__50621));
    InMux I__10721 (
            .O(N__50640),
            .I(N__50616));
    InMux I__10720 (
            .O(N__50639),
            .I(N__50616));
    LocalMux I__10719 (
            .O(N__50636),
            .I(\c0.data_in_frame_3_1 ));
    Odrv12 I__10718 (
            .O(N__50633),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__10717 (
            .O(N__50624),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__10716 (
            .O(N__50621),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__10715 (
            .O(N__50616),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__10714 (
            .O(N__50605),
            .I(N__50596));
    InMux I__10713 (
            .O(N__50604),
            .I(N__50593));
    InMux I__10712 (
            .O(N__50603),
            .I(N__50589));
    InMux I__10711 (
            .O(N__50602),
            .I(N__50586));
    InMux I__10710 (
            .O(N__50601),
            .I(N__50583));
    CascadeMux I__10709 (
            .O(N__50600),
            .I(N__50579));
    CascadeMux I__10708 (
            .O(N__50599),
            .I(N__50576));
    LocalMux I__10707 (
            .O(N__50596),
            .I(N__50573));
    LocalMux I__10706 (
            .O(N__50593),
            .I(N__50570));
    InMux I__10705 (
            .O(N__50592),
            .I(N__50567));
    LocalMux I__10704 (
            .O(N__50589),
            .I(N__50563));
    LocalMux I__10703 (
            .O(N__50586),
            .I(N__50558));
    LocalMux I__10702 (
            .O(N__50583),
            .I(N__50558));
    CascadeMux I__10701 (
            .O(N__50582),
            .I(N__50555));
    InMux I__10700 (
            .O(N__50579),
            .I(N__50545));
    InMux I__10699 (
            .O(N__50576),
            .I(N__50545));
    Span4Mux_h I__10698 (
            .O(N__50573),
            .I(N__50538));
    Span4Mux_h I__10697 (
            .O(N__50570),
            .I(N__50538));
    LocalMux I__10696 (
            .O(N__50567),
            .I(N__50538));
    InMux I__10695 (
            .O(N__50566),
            .I(N__50535));
    Span4Mux_h I__10694 (
            .O(N__50563),
            .I(N__50530));
    Span4Mux_v I__10693 (
            .O(N__50558),
            .I(N__50530));
    InMux I__10692 (
            .O(N__50555),
            .I(N__50525));
    InMux I__10691 (
            .O(N__50554),
            .I(N__50525));
    InMux I__10690 (
            .O(N__50553),
            .I(N__50518));
    InMux I__10689 (
            .O(N__50552),
            .I(N__50518));
    InMux I__10688 (
            .O(N__50551),
            .I(N__50518));
    InMux I__10687 (
            .O(N__50550),
            .I(N__50515));
    LocalMux I__10686 (
            .O(N__50545),
            .I(data_in_frame_0_5));
    Odrv4 I__10685 (
            .O(N__50538),
            .I(data_in_frame_0_5));
    LocalMux I__10684 (
            .O(N__50535),
            .I(data_in_frame_0_5));
    Odrv4 I__10683 (
            .O(N__50530),
            .I(data_in_frame_0_5));
    LocalMux I__10682 (
            .O(N__50525),
            .I(data_in_frame_0_5));
    LocalMux I__10681 (
            .O(N__50518),
            .I(data_in_frame_0_5));
    LocalMux I__10680 (
            .O(N__50515),
            .I(data_in_frame_0_5));
    InMux I__10679 (
            .O(N__50500),
            .I(N__50497));
    LocalMux I__10678 (
            .O(N__50497),
            .I(N__50493));
    InMux I__10677 (
            .O(N__50496),
            .I(N__50490));
    Span4Mux_h I__10676 (
            .O(N__50493),
            .I(N__50487));
    LocalMux I__10675 (
            .O(N__50490),
            .I(N__50482));
    Span4Mux_h I__10674 (
            .O(N__50487),
            .I(N__50479));
    InMux I__10673 (
            .O(N__50486),
            .I(N__50474));
    InMux I__10672 (
            .O(N__50485),
            .I(N__50474));
    Odrv12 I__10671 (
            .O(N__50482),
            .I(\c0.n33_adj_3088 ));
    Odrv4 I__10670 (
            .O(N__50479),
            .I(\c0.n33_adj_3088 ));
    LocalMux I__10669 (
            .O(N__50474),
            .I(\c0.n33_adj_3088 ));
    InMux I__10668 (
            .O(N__50467),
            .I(N__50464));
    LocalMux I__10667 (
            .O(N__50464),
            .I(\c0.n15_adj_3545 ));
    InMux I__10666 (
            .O(N__50461),
            .I(N__50458));
    LocalMux I__10665 (
            .O(N__50458),
            .I(N__50453));
    InMux I__10664 (
            .O(N__50457),
            .I(N__50450));
    CascadeMux I__10663 (
            .O(N__50456),
            .I(N__50447));
    Span4Mux_v I__10662 (
            .O(N__50453),
            .I(N__50442));
    LocalMux I__10661 (
            .O(N__50450),
            .I(N__50442));
    InMux I__10660 (
            .O(N__50447),
            .I(N__50439));
    Odrv4 I__10659 (
            .O(N__50442),
            .I(\c0.n24_adj_3013 ));
    LocalMux I__10658 (
            .O(N__50439),
            .I(\c0.n24_adj_3013 ));
    CascadeMux I__10657 (
            .O(N__50434),
            .I(N__50429));
    CascadeMux I__10656 (
            .O(N__50433),
            .I(N__50426));
    CascadeMux I__10655 (
            .O(N__50432),
            .I(N__50422));
    InMux I__10654 (
            .O(N__50429),
            .I(N__50419));
    InMux I__10653 (
            .O(N__50426),
            .I(N__50412));
    InMux I__10652 (
            .O(N__50425),
            .I(N__50412));
    InMux I__10651 (
            .O(N__50422),
            .I(N__50412));
    LocalMux I__10650 (
            .O(N__50419),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__10649 (
            .O(N__50412),
            .I(\c0.data_in_frame_3_3 ));
    InMux I__10648 (
            .O(N__50407),
            .I(N__50402));
    CascadeMux I__10647 (
            .O(N__50406),
            .I(N__50399));
    InMux I__10646 (
            .O(N__50405),
            .I(N__50396));
    LocalMux I__10645 (
            .O(N__50402),
            .I(N__50390));
    InMux I__10644 (
            .O(N__50399),
            .I(N__50387));
    LocalMux I__10643 (
            .O(N__50396),
            .I(N__50384));
    InMux I__10642 (
            .O(N__50395),
            .I(N__50379));
    InMux I__10641 (
            .O(N__50394),
            .I(N__50379));
    InMux I__10640 (
            .O(N__50393),
            .I(N__50376));
    Span4Mux_v I__10639 (
            .O(N__50390),
            .I(N__50371));
    LocalMux I__10638 (
            .O(N__50387),
            .I(N__50371));
    Odrv4 I__10637 (
            .O(N__50384),
            .I(\c0.data_in_frame_3_2 ));
    LocalMux I__10636 (
            .O(N__50379),
            .I(\c0.data_in_frame_3_2 ));
    LocalMux I__10635 (
            .O(N__50376),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__10634 (
            .O(N__50371),
            .I(\c0.data_in_frame_3_2 ));
    InMux I__10633 (
            .O(N__50362),
            .I(N__50356));
    InMux I__10632 (
            .O(N__50361),
            .I(N__50353));
    InMux I__10631 (
            .O(N__50360),
            .I(N__50350));
    CascadeMux I__10630 (
            .O(N__50359),
            .I(N__50343));
    LocalMux I__10629 (
            .O(N__50356),
            .I(N__50340));
    LocalMux I__10628 (
            .O(N__50353),
            .I(N__50336));
    LocalMux I__10627 (
            .O(N__50350),
            .I(N__50333));
    InMux I__10626 (
            .O(N__50349),
            .I(N__50329));
    InMux I__10625 (
            .O(N__50348),
            .I(N__50326));
    InMux I__10624 (
            .O(N__50347),
            .I(N__50321));
    InMux I__10623 (
            .O(N__50346),
            .I(N__50321));
    InMux I__10622 (
            .O(N__50343),
            .I(N__50318));
    Span12Mux_v I__10621 (
            .O(N__50340),
            .I(N__50314));
    InMux I__10620 (
            .O(N__50339),
            .I(N__50310));
    Span4Mux_h I__10619 (
            .O(N__50336),
            .I(N__50305));
    Span4Mux_v I__10618 (
            .O(N__50333),
            .I(N__50305));
    InMux I__10617 (
            .O(N__50332),
            .I(N__50302));
    LocalMux I__10616 (
            .O(N__50329),
            .I(N__50297));
    LocalMux I__10615 (
            .O(N__50326),
            .I(N__50290));
    LocalMux I__10614 (
            .O(N__50321),
            .I(N__50290));
    LocalMux I__10613 (
            .O(N__50318),
            .I(N__50290));
    InMux I__10612 (
            .O(N__50317),
            .I(N__50287));
    Span12Mux_h I__10611 (
            .O(N__50314),
            .I(N__50282));
    InMux I__10610 (
            .O(N__50313),
            .I(N__50279));
    LocalMux I__10609 (
            .O(N__50310),
            .I(N__50272));
    Span4Mux_h I__10608 (
            .O(N__50305),
            .I(N__50272));
    LocalMux I__10607 (
            .O(N__50302),
            .I(N__50272));
    InMux I__10606 (
            .O(N__50301),
            .I(N__50267));
    InMux I__10605 (
            .O(N__50300),
            .I(N__50267));
    Span4Mux_v I__10604 (
            .O(N__50297),
            .I(N__50260));
    Span4Mux_v I__10603 (
            .O(N__50290),
            .I(N__50260));
    LocalMux I__10602 (
            .O(N__50287),
            .I(N__50260));
    InMux I__10601 (
            .O(N__50286),
            .I(N__50257));
    InMux I__10600 (
            .O(N__50285),
            .I(N__50254));
    Odrv12 I__10599 (
            .O(N__50282),
            .I(data_out_frame_29__3__N_647));
    LocalMux I__10598 (
            .O(N__50279),
            .I(data_out_frame_29__3__N_647));
    Odrv4 I__10597 (
            .O(N__50272),
            .I(data_out_frame_29__3__N_647));
    LocalMux I__10596 (
            .O(N__50267),
            .I(data_out_frame_29__3__N_647));
    Odrv4 I__10595 (
            .O(N__50260),
            .I(data_out_frame_29__3__N_647));
    LocalMux I__10594 (
            .O(N__50257),
            .I(data_out_frame_29__3__N_647));
    LocalMux I__10593 (
            .O(N__50254),
            .I(data_out_frame_29__3__N_647));
    InMux I__10592 (
            .O(N__50239),
            .I(N__50236));
    LocalMux I__10591 (
            .O(N__50236),
            .I(N__50233));
    Odrv12 I__10590 (
            .O(N__50233),
            .I(\c0.n29_adj_3216 ));
    InMux I__10589 (
            .O(N__50230),
            .I(N__50227));
    LocalMux I__10588 (
            .O(N__50227),
            .I(N__50223));
    InMux I__10587 (
            .O(N__50226),
            .I(N__50220));
    Span4Mux_v I__10586 (
            .O(N__50223),
            .I(N__50217));
    LocalMux I__10585 (
            .O(N__50220),
            .I(N__50214));
    Odrv4 I__10584 (
            .O(N__50217),
            .I(\c0.n78 ));
    Odrv12 I__10583 (
            .O(N__50214),
            .I(\c0.n78 ));
    InMux I__10582 (
            .O(N__50209),
            .I(N__50206));
    LocalMux I__10581 (
            .O(N__50206),
            .I(N__50203));
    Span4Mux_v I__10580 (
            .O(N__50203),
            .I(N__50200));
    Sp12to4 I__10579 (
            .O(N__50200),
            .I(N__50197));
    Odrv12 I__10578 (
            .O(N__50197),
            .I(\c0.n37_adj_3215 ));
    CascadeMux I__10577 (
            .O(N__50194),
            .I(\c0.n29_adj_3216_cascade_ ));
    InMux I__10576 (
            .O(N__50191),
            .I(N__50188));
    LocalMux I__10575 (
            .O(N__50188),
            .I(\c0.n44_adj_3217 ));
    CascadeMux I__10574 (
            .O(N__50185),
            .I(\c0.n8_adj_3066_cascade_ ));
    InMux I__10573 (
            .O(N__50182),
            .I(N__50179));
    LocalMux I__10572 (
            .O(N__50179),
            .I(N__50176));
    Span4Mux_v I__10571 (
            .O(N__50176),
            .I(N__50172));
    InMux I__10570 (
            .O(N__50175),
            .I(N__50169));
    Span4Mux_h I__10569 (
            .O(N__50172),
            .I(N__50164));
    LocalMux I__10568 (
            .O(N__50169),
            .I(N__50164));
    Odrv4 I__10567 (
            .O(N__50164),
            .I(\c0.n19170 ));
    CascadeMux I__10566 (
            .O(N__50161),
            .I(\c0.n19170_cascade_ ));
    CascadeMux I__10565 (
            .O(N__50158),
            .I(N__50154));
    InMux I__10564 (
            .O(N__50157),
            .I(N__50151));
    InMux I__10563 (
            .O(N__50154),
            .I(N__50146));
    LocalMux I__10562 (
            .O(N__50151),
            .I(N__50143));
    InMux I__10561 (
            .O(N__50150),
            .I(N__50140));
    CascadeMux I__10560 (
            .O(N__50149),
            .I(N__50137));
    LocalMux I__10559 (
            .O(N__50146),
            .I(N__50134));
    Span4Mux_v I__10558 (
            .O(N__50143),
            .I(N__50129));
    LocalMux I__10557 (
            .O(N__50140),
            .I(N__50129));
    InMux I__10556 (
            .O(N__50137),
            .I(N__50126));
    Span4Mux_v I__10555 (
            .O(N__50134),
            .I(N__50123));
    Span4Mux_h I__10554 (
            .O(N__50129),
            .I(N__50120));
    LocalMux I__10553 (
            .O(N__50126),
            .I(\c0.data_in_frame_8_2 ));
    Odrv4 I__10552 (
            .O(N__50123),
            .I(\c0.data_in_frame_8_2 ));
    Odrv4 I__10551 (
            .O(N__50120),
            .I(\c0.data_in_frame_8_2 ));
    InMux I__10550 (
            .O(N__50113),
            .I(N__50110));
    LocalMux I__10549 (
            .O(N__50110),
            .I(N__50105));
    InMux I__10548 (
            .O(N__50109),
            .I(N__50102));
    InMux I__10547 (
            .O(N__50108),
            .I(N__50099));
    Span4Mux_v I__10546 (
            .O(N__50105),
            .I(N__50092));
    LocalMux I__10545 (
            .O(N__50102),
            .I(N__50092));
    LocalMux I__10544 (
            .O(N__50099),
            .I(N__50092));
    Span4Mux_h I__10543 (
            .O(N__50092),
            .I(N__50089));
    Odrv4 I__10542 (
            .O(N__50089),
            .I(\c0.n21_adj_3053 ));
    CascadeMux I__10541 (
            .O(N__50086),
            .I(N__50083));
    InMux I__10540 (
            .O(N__50083),
            .I(N__50078));
    InMux I__10539 (
            .O(N__50082),
            .I(N__50073));
    CascadeMux I__10538 (
            .O(N__50081),
            .I(N__50070));
    LocalMux I__10537 (
            .O(N__50078),
            .I(N__50067));
    InMux I__10536 (
            .O(N__50077),
            .I(N__50064));
    InMux I__10535 (
            .O(N__50076),
            .I(N__50060));
    LocalMux I__10534 (
            .O(N__50073),
            .I(N__50057));
    InMux I__10533 (
            .O(N__50070),
            .I(N__50054));
    Span4Mux_v I__10532 (
            .O(N__50067),
            .I(N__50049));
    LocalMux I__10531 (
            .O(N__50064),
            .I(N__50049));
    InMux I__10530 (
            .O(N__50063),
            .I(N__50046));
    LocalMux I__10529 (
            .O(N__50060),
            .I(N__50043));
    Span4Mux_h I__10528 (
            .O(N__50057),
            .I(N__50038));
    LocalMux I__10527 (
            .O(N__50054),
            .I(N__50038));
    Span4Mux_v I__10526 (
            .O(N__50049),
            .I(N__50033));
    LocalMux I__10525 (
            .O(N__50046),
            .I(N__50033));
    Span4Mux_h I__10524 (
            .O(N__50043),
            .I(N__50026));
    Span4Mux_v I__10523 (
            .O(N__50038),
            .I(N__50026));
    Span4Mux_h I__10522 (
            .O(N__50033),
            .I(N__50026));
    Odrv4 I__10521 (
            .O(N__50026),
            .I(\c0.n21 ));
    CascadeMux I__10520 (
            .O(N__50023),
            .I(N__50019));
    InMux I__10519 (
            .O(N__50022),
            .I(N__50016));
    InMux I__10518 (
            .O(N__50019),
            .I(N__50013));
    LocalMux I__10517 (
            .O(N__50016),
            .I(N__50010));
    LocalMux I__10516 (
            .O(N__50013),
            .I(\c0.data_in_frame_5_4 ));
    Odrv4 I__10515 (
            .O(N__50010),
            .I(\c0.data_in_frame_5_4 ));
    CascadeMux I__10514 (
            .O(N__50005),
            .I(N__50001));
    InMux I__10513 (
            .O(N__50004),
            .I(N__49998));
    InMux I__10512 (
            .O(N__50001),
            .I(N__49995));
    LocalMux I__10511 (
            .O(N__49998),
            .I(\c0.n25 ));
    LocalMux I__10510 (
            .O(N__49995),
            .I(\c0.n25 ));
    InMux I__10509 (
            .O(N__49990),
            .I(N__49987));
    LocalMux I__10508 (
            .O(N__49987),
            .I(\c0.n89 ));
    CascadeMux I__10507 (
            .O(N__49984),
            .I(N__49981));
    InMux I__10506 (
            .O(N__49981),
            .I(N__49976));
    InMux I__10505 (
            .O(N__49980),
            .I(N__49971));
    InMux I__10504 (
            .O(N__49979),
            .I(N__49968));
    LocalMux I__10503 (
            .O(N__49976),
            .I(N__49965));
    InMux I__10502 (
            .O(N__49975),
            .I(N__49960));
    InMux I__10501 (
            .O(N__49974),
            .I(N__49960));
    LocalMux I__10500 (
            .O(N__49971),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__10499 (
            .O(N__49968),
            .I(\c0.data_in_frame_4_0 ));
    Odrv4 I__10498 (
            .O(N__49965),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__10497 (
            .O(N__49960),
            .I(\c0.data_in_frame_4_0 ));
    InMux I__10496 (
            .O(N__49951),
            .I(N__49948));
    LocalMux I__10495 (
            .O(N__49948),
            .I(N__49945));
    Span4Mux_v I__10494 (
            .O(N__49945),
            .I(N__49942));
    Odrv4 I__10493 (
            .O(N__49942),
            .I(\c0.n17_adj_3113 ));
    InMux I__10492 (
            .O(N__49939),
            .I(N__49936));
    LocalMux I__10491 (
            .O(N__49936),
            .I(\c0.n5_adj_3030 ));
    CascadeMux I__10490 (
            .O(N__49933),
            .I(\c0.n60_cascade_ ));
    InMux I__10489 (
            .O(N__49930),
            .I(N__49927));
    LocalMux I__10488 (
            .O(N__49927),
            .I(N__49924));
    Odrv4 I__10487 (
            .O(N__49924),
            .I(\c0.n93 ));
    InMux I__10486 (
            .O(N__49921),
            .I(N__49918));
    LocalMux I__10485 (
            .O(N__49918),
            .I(N__49913));
    InMux I__10484 (
            .O(N__49917),
            .I(N__49910));
    InMux I__10483 (
            .O(N__49916),
            .I(N__49907));
    Span4Mux_v I__10482 (
            .O(N__49913),
            .I(N__49903));
    LocalMux I__10481 (
            .O(N__49910),
            .I(N__49900));
    LocalMux I__10480 (
            .O(N__49907),
            .I(N__49897));
    InMux I__10479 (
            .O(N__49906),
            .I(N__49894));
    Span4Mux_v I__10478 (
            .O(N__49903),
            .I(N__49891));
    Span4Mux_h I__10477 (
            .O(N__49900),
            .I(N__49886));
    Span4Mux_h I__10476 (
            .O(N__49897),
            .I(N__49886));
    LocalMux I__10475 (
            .O(N__49894),
            .I(\c0.data_in_frame_6_1 ));
    Odrv4 I__10474 (
            .O(N__49891),
            .I(\c0.data_in_frame_6_1 ));
    Odrv4 I__10473 (
            .O(N__49886),
            .I(\c0.data_in_frame_6_1 ));
    InMux I__10472 (
            .O(N__49879),
            .I(N__49876));
    LocalMux I__10471 (
            .O(N__49876),
            .I(N__49872));
    CascadeMux I__10470 (
            .O(N__49875),
            .I(N__49869));
    Span4Mux_v I__10469 (
            .O(N__49872),
            .I(N__49866));
    InMux I__10468 (
            .O(N__49869),
            .I(N__49863));
    Odrv4 I__10467 (
            .O(N__49866),
            .I(\c0.n5_adj_3028 ));
    LocalMux I__10466 (
            .O(N__49863),
            .I(\c0.n5_adj_3028 ));
    InMux I__10465 (
            .O(N__49858),
            .I(N__49855));
    LocalMux I__10464 (
            .O(N__49855),
            .I(N__49852));
    Span4Mux_h I__10463 (
            .O(N__49852),
            .I(N__49848));
    InMux I__10462 (
            .O(N__49851),
            .I(N__49844));
    Span4Mux_v I__10461 (
            .O(N__49848),
            .I(N__49841));
    InMux I__10460 (
            .O(N__49847),
            .I(N__49838));
    LocalMux I__10459 (
            .O(N__49844),
            .I(N__49835));
    Odrv4 I__10458 (
            .O(N__49841),
            .I(\c0.n19443 ));
    LocalMux I__10457 (
            .O(N__49838),
            .I(\c0.n19443 ));
    Odrv4 I__10456 (
            .O(N__49835),
            .I(\c0.n19443 ));
    InMux I__10455 (
            .O(N__49828),
            .I(N__49825));
    LocalMux I__10454 (
            .O(N__49825),
            .I(N__49822));
    Span4Mux_v I__10453 (
            .O(N__49822),
            .I(N__49819));
    Span4Mux_h I__10452 (
            .O(N__49819),
            .I(N__49816));
    Odrv4 I__10451 (
            .O(N__49816),
            .I(\c0.n11687 ));
    InMux I__10450 (
            .O(N__49813),
            .I(N__49810));
    LocalMux I__10449 (
            .O(N__49810),
            .I(N__49806));
    CascadeMux I__10448 (
            .O(N__49809),
            .I(N__49803));
    Span4Mux_v I__10447 (
            .O(N__49806),
            .I(N__49799));
    InMux I__10446 (
            .O(N__49803),
            .I(N__49794));
    InMux I__10445 (
            .O(N__49802),
            .I(N__49794));
    Odrv4 I__10444 (
            .O(N__49799),
            .I(\c0.n20313 ));
    LocalMux I__10443 (
            .O(N__49794),
            .I(\c0.n20313 ));
    InMux I__10442 (
            .O(N__49789),
            .I(N__49786));
    LocalMux I__10441 (
            .O(N__49786),
            .I(N__49782));
    CascadeMux I__10440 (
            .O(N__49785),
            .I(N__49778));
    Span4Mux_h I__10439 (
            .O(N__49782),
            .I(N__49775));
    InMux I__10438 (
            .O(N__49781),
            .I(N__49770));
    InMux I__10437 (
            .O(N__49778),
            .I(N__49770));
    Odrv4 I__10436 (
            .O(N__49775),
            .I(\c0.data_in_frame_26_5 ));
    LocalMux I__10435 (
            .O(N__49770),
            .I(\c0.data_in_frame_26_5 ));
    InMux I__10434 (
            .O(N__49765),
            .I(N__49762));
    LocalMux I__10433 (
            .O(N__49762),
            .I(N__49759));
    Odrv4 I__10432 (
            .O(N__49759),
            .I(\c0.n17840 ));
    InMux I__10431 (
            .O(N__49756),
            .I(N__49751));
    InMux I__10430 (
            .O(N__49755),
            .I(N__49748));
    InMux I__10429 (
            .O(N__49754),
            .I(N__49745));
    LocalMux I__10428 (
            .O(N__49751),
            .I(N__49741));
    LocalMux I__10427 (
            .O(N__49748),
            .I(N__49738));
    LocalMux I__10426 (
            .O(N__49745),
            .I(N__49735));
    CascadeMux I__10425 (
            .O(N__49744),
            .I(N__49731));
    Span4Mux_v I__10424 (
            .O(N__49741),
            .I(N__49723));
    Span4Mux_v I__10423 (
            .O(N__49738),
            .I(N__49723));
    Span4Mux_v I__10422 (
            .O(N__49735),
            .I(N__49723));
    InMux I__10421 (
            .O(N__49734),
            .I(N__49720));
    InMux I__10420 (
            .O(N__49731),
            .I(N__49717));
    InMux I__10419 (
            .O(N__49730),
            .I(N__49714));
    Span4Mux_h I__10418 (
            .O(N__49723),
            .I(N__49711));
    LocalMux I__10417 (
            .O(N__49720),
            .I(N__49706));
    LocalMux I__10416 (
            .O(N__49717),
            .I(N__49706));
    LocalMux I__10415 (
            .O(N__49714),
            .I(data_in_3_0));
    Odrv4 I__10414 (
            .O(N__49711),
            .I(data_in_3_0));
    Odrv12 I__10413 (
            .O(N__49706),
            .I(data_in_3_0));
    InMux I__10412 (
            .O(N__49699),
            .I(N__49696));
    LocalMux I__10411 (
            .O(N__49696),
            .I(N__49693));
    Span4Mux_v I__10410 (
            .O(N__49693),
            .I(N__49688));
    InMux I__10409 (
            .O(N__49692),
            .I(N__49683));
    InMux I__10408 (
            .O(N__49691),
            .I(N__49683));
    Odrv4 I__10407 (
            .O(N__49688),
            .I(\c0.n12_adj_3498 ));
    LocalMux I__10406 (
            .O(N__49683),
            .I(\c0.n12_adj_3498 ));
    CascadeMux I__10405 (
            .O(N__49678),
            .I(N__49673));
    InMux I__10404 (
            .O(N__49677),
            .I(N__49669));
    InMux I__10403 (
            .O(N__49676),
            .I(N__49666));
    InMux I__10402 (
            .O(N__49673),
            .I(N__49662));
    InMux I__10401 (
            .O(N__49672),
            .I(N__49659));
    LocalMux I__10400 (
            .O(N__49669),
            .I(N__49656));
    LocalMux I__10399 (
            .O(N__49666),
            .I(N__49652));
    InMux I__10398 (
            .O(N__49665),
            .I(N__49649));
    LocalMux I__10397 (
            .O(N__49662),
            .I(N__49644));
    LocalMux I__10396 (
            .O(N__49659),
            .I(N__49644));
    Span4Mux_v I__10395 (
            .O(N__49656),
            .I(N__49641));
    InMux I__10394 (
            .O(N__49655),
            .I(N__49638));
    Span4Mux_h I__10393 (
            .O(N__49652),
            .I(N__49633));
    LocalMux I__10392 (
            .O(N__49649),
            .I(N__49633));
    Span4Mux_v I__10391 (
            .O(N__49644),
            .I(N__49630));
    Span4Mux_v I__10390 (
            .O(N__49641),
            .I(N__49627));
    LocalMux I__10389 (
            .O(N__49638),
            .I(N__49624));
    Span4Mux_h I__10388 (
            .O(N__49633),
            .I(N__49619));
    Span4Mux_v I__10387 (
            .O(N__49630),
            .I(N__49619));
    Span4Mux_v I__10386 (
            .O(N__49627),
            .I(N__49615));
    Span4Mux_h I__10385 (
            .O(N__49624),
            .I(N__49612));
    Span4Mux_v I__10384 (
            .O(N__49619),
            .I(N__49609));
    InMux I__10383 (
            .O(N__49618),
            .I(N__49606));
    Odrv4 I__10382 (
            .O(N__49615),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv4 I__10381 (
            .O(N__49612),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv4 I__10380 (
            .O(N__49609),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__10379 (
            .O(N__49606),
            .I(\c0.FRAME_MATCHER_i_5 ));
    SRMux I__10378 (
            .O(N__49597),
            .I(N__49594));
    LocalMux I__10377 (
            .O(N__49594),
            .I(N__49591));
    Sp12to4 I__10376 (
            .O(N__49591),
            .I(N__49588));
    Span12Mux_s7_v I__10375 (
            .O(N__49588),
            .I(N__49585));
    Odrv12 I__10374 (
            .O(N__49585),
            .I(\c0.n6_adj_3149 ));
    CascadeMux I__10373 (
            .O(N__49582),
            .I(N__49578));
    CascadeMux I__10372 (
            .O(N__49581),
            .I(N__49574));
    InMux I__10371 (
            .O(N__49578),
            .I(N__49571));
    InMux I__10370 (
            .O(N__49577),
            .I(N__49566));
    InMux I__10369 (
            .O(N__49574),
            .I(N__49566));
    LocalMux I__10368 (
            .O(N__49571),
            .I(N__49563));
    LocalMux I__10367 (
            .O(N__49566),
            .I(N__49560));
    Span4Mux_h I__10366 (
            .O(N__49563),
            .I(N__49553));
    Span4Mux_v I__10365 (
            .O(N__49560),
            .I(N__49553));
    InMux I__10364 (
            .O(N__49559),
            .I(N__49548));
    InMux I__10363 (
            .O(N__49558),
            .I(N__49548));
    Odrv4 I__10362 (
            .O(N__49553),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__10361 (
            .O(N__49548),
            .I(\c0.data_in_frame_8_6 ));
    InMux I__10360 (
            .O(N__49543),
            .I(N__49540));
    LocalMux I__10359 (
            .O(N__49540),
            .I(N__49537));
    Span4Mux_h I__10358 (
            .O(N__49537),
            .I(N__49532));
    InMux I__10357 (
            .O(N__49536),
            .I(N__49527));
    InMux I__10356 (
            .O(N__49535),
            .I(N__49527));
    Odrv4 I__10355 (
            .O(N__49532),
            .I(\c0.n11936 ));
    LocalMux I__10354 (
            .O(N__49527),
            .I(\c0.n11936 ));
    CascadeMux I__10353 (
            .O(N__49522),
            .I(N__49519));
    InMux I__10352 (
            .O(N__49519),
            .I(N__49516));
    LocalMux I__10351 (
            .O(N__49516),
            .I(N__49513));
    Span4Mux_h I__10350 (
            .O(N__49513),
            .I(N__49510));
    Odrv4 I__10349 (
            .O(N__49510),
            .I(\c0.n12_adj_3141 ));
    InMux I__10348 (
            .O(N__49507),
            .I(N__49502));
    InMux I__10347 (
            .O(N__49506),
            .I(N__49499));
    InMux I__10346 (
            .O(N__49505),
            .I(N__49495));
    LocalMux I__10345 (
            .O(N__49502),
            .I(N__49492));
    LocalMux I__10344 (
            .O(N__49499),
            .I(N__49488));
    InMux I__10343 (
            .O(N__49498),
            .I(N__49484));
    LocalMux I__10342 (
            .O(N__49495),
            .I(N__49479));
    Span4Mux_v I__10341 (
            .O(N__49492),
            .I(N__49479));
    InMux I__10340 (
            .O(N__49491),
            .I(N__49476));
    Span4Mux_v I__10339 (
            .O(N__49488),
            .I(N__49473));
    InMux I__10338 (
            .O(N__49487),
            .I(N__49470));
    LocalMux I__10337 (
            .O(N__49484),
            .I(data_in_frame_24_6));
    Odrv4 I__10336 (
            .O(N__49479),
            .I(data_in_frame_24_6));
    LocalMux I__10335 (
            .O(N__49476),
            .I(data_in_frame_24_6));
    Odrv4 I__10334 (
            .O(N__49473),
            .I(data_in_frame_24_6));
    LocalMux I__10333 (
            .O(N__49470),
            .I(data_in_frame_24_6));
    InMux I__10332 (
            .O(N__49459),
            .I(N__49455));
    InMux I__10331 (
            .O(N__49458),
            .I(N__49451));
    LocalMux I__10330 (
            .O(N__49455),
            .I(N__49448));
    InMux I__10329 (
            .O(N__49454),
            .I(N__49445));
    LocalMux I__10328 (
            .O(N__49451),
            .I(N__49441));
    Span4Mux_v I__10327 (
            .O(N__49448),
            .I(N__49436));
    LocalMux I__10326 (
            .O(N__49445),
            .I(N__49436));
    InMux I__10325 (
            .O(N__49444),
            .I(N__49432));
    Span4Mux_h I__10324 (
            .O(N__49441),
            .I(N__49429));
    Span4Mux_h I__10323 (
            .O(N__49436),
            .I(N__49426));
    InMux I__10322 (
            .O(N__49435),
            .I(N__49423));
    LocalMux I__10321 (
            .O(N__49432),
            .I(data_in_frame_24_4));
    Odrv4 I__10320 (
            .O(N__49429),
            .I(data_in_frame_24_4));
    Odrv4 I__10319 (
            .O(N__49426),
            .I(data_in_frame_24_4));
    LocalMux I__10318 (
            .O(N__49423),
            .I(data_in_frame_24_4));
    CascadeMux I__10317 (
            .O(N__49414),
            .I(\c0.n19465_cascade_ ));
    InMux I__10316 (
            .O(N__49411),
            .I(N__49408));
    LocalMux I__10315 (
            .O(N__49408),
            .I(N__49405));
    Odrv4 I__10314 (
            .O(N__49405),
            .I(\c0.n17 ));
    InMux I__10313 (
            .O(N__49402),
            .I(N__49398));
    InMux I__10312 (
            .O(N__49401),
            .I(N__49393));
    LocalMux I__10311 (
            .O(N__49398),
            .I(N__49390));
    InMux I__10310 (
            .O(N__49397),
            .I(N__49387));
    InMux I__10309 (
            .O(N__49396),
            .I(N__49384));
    LocalMux I__10308 (
            .O(N__49393),
            .I(\c0.n21044 ));
    Odrv4 I__10307 (
            .O(N__49390),
            .I(\c0.n21044 ));
    LocalMux I__10306 (
            .O(N__49387),
            .I(\c0.n21044 ));
    LocalMux I__10305 (
            .O(N__49384),
            .I(\c0.n21044 ));
    InMux I__10304 (
            .O(N__49375),
            .I(N__49372));
    LocalMux I__10303 (
            .O(N__49372),
            .I(N__49368));
    InMux I__10302 (
            .O(N__49371),
            .I(N__49365));
    Span4Mux_h I__10301 (
            .O(N__49368),
            .I(N__49362));
    LocalMux I__10300 (
            .O(N__49365),
            .I(\c0.n19703 ));
    Odrv4 I__10299 (
            .O(N__49362),
            .I(\c0.n19703 ));
    CascadeMux I__10298 (
            .O(N__49357),
            .I(\c0.n19703_cascade_ ));
    InMux I__10297 (
            .O(N__49354),
            .I(N__49351));
    LocalMux I__10296 (
            .O(N__49351),
            .I(\c0.n44_adj_3278 ));
    CascadeMux I__10295 (
            .O(N__49348),
            .I(N__49343));
    InMux I__10294 (
            .O(N__49347),
            .I(N__49340));
    InMux I__10293 (
            .O(N__49346),
            .I(N__49337));
    InMux I__10292 (
            .O(N__49343),
            .I(N__49334));
    LocalMux I__10291 (
            .O(N__49340),
            .I(N__49329));
    LocalMux I__10290 (
            .O(N__49337),
            .I(N__49329));
    LocalMux I__10289 (
            .O(N__49334),
            .I(N__49323));
    Span4Mux_h I__10288 (
            .O(N__49329),
            .I(N__49320));
    InMux I__10287 (
            .O(N__49328),
            .I(N__49317));
    InMux I__10286 (
            .O(N__49327),
            .I(N__49312));
    InMux I__10285 (
            .O(N__49326),
            .I(N__49312));
    Odrv4 I__10284 (
            .O(N__49323),
            .I(\c0.data_in_frame_25_1 ));
    Odrv4 I__10283 (
            .O(N__49320),
            .I(\c0.data_in_frame_25_1 ));
    LocalMux I__10282 (
            .O(N__49317),
            .I(\c0.data_in_frame_25_1 ));
    LocalMux I__10281 (
            .O(N__49312),
            .I(\c0.data_in_frame_25_1 ));
    CascadeMux I__10280 (
            .O(N__49303),
            .I(N__49298));
    InMux I__10279 (
            .O(N__49302),
            .I(N__49295));
    InMux I__10278 (
            .O(N__49301),
            .I(N__49292));
    InMux I__10277 (
            .O(N__49298),
            .I(N__49289));
    LocalMux I__10276 (
            .O(N__49295),
            .I(N__49285));
    LocalMux I__10275 (
            .O(N__49292),
            .I(N__49282));
    LocalMux I__10274 (
            .O(N__49289),
            .I(N__49279));
    InMux I__10273 (
            .O(N__49288),
            .I(N__49276));
    Span4Mux_h I__10272 (
            .O(N__49285),
            .I(N__49269));
    Span4Mux_v I__10271 (
            .O(N__49282),
            .I(N__49269));
    Span4Mux_h I__10270 (
            .O(N__49279),
            .I(N__49269));
    LocalMux I__10269 (
            .O(N__49276),
            .I(N__49266));
    Odrv4 I__10268 (
            .O(N__49269),
            .I(\c0.n18377 ));
    Odrv4 I__10267 (
            .O(N__49266),
            .I(\c0.n18377 ));
    InMux I__10266 (
            .O(N__49261),
            .I(N__49252));
    InMux I__10265 (
            .O(N__49260),
            .I(N__49252));
    InMux I__10264 (
            .O(N__49259),
            .I(N__49249));
    InMux I__10263 (
            .O(N__49258),
            .I(N__49246));
    InMux I__10262 (
            .O(N__49257),
            .I(N__49243));
    LocalMux I__10261 (
            .O(N__49252),
            .I(N__49240));
    LocalMux I__10260 (
            .O(N__49249),
            .I(\c0.data_in_frame_25_2 ));
    LocalMux I__10259 (
            .O(N__49246),
            .I(\c0.data_in_frame_25_2 ));
    LocalMux I__10258 (
            .O(N__49243),
            .I(\c0.data_in_frame_25_2 ));
    Odrv4 I__10257 (
            .O(N__49240),
            .I(\c0.data_in_frame_25_2 ));
    InMux I__10256 (
            .O(N__49231),
            .I(N__49222));
    InMux I__10255 (
            .O(N__49230),
            .I(N__49222));
    InMux I__10254 (
            .O(N__49229),
            .I(N__49219));
    InMux I__10253 (
            .O(N__49228),
            .I(N__49214));
    InMux I__10252 (
            .O(N__49227),
            .I(N__49214));
    LocalMux I__10251 (
            .O(N__49222),
            .I(N__49210));
    LocalMux I__10250 (
            .O(N__49219),
            .I(N__49205));
    LocalMux I__10249 (
            .O(N__49214),
            .I(N__49205));
    CascadeMux I__10248 (
            .O(N__49213),
            .I(N__49202));
    Span4Mux_v I__10247 (
            .O(N__49210),
            .I(N__49199));
    Span4Mux_v I__10246 (
            .O(N__49205),
            .I(N__49196));
    InMux I__10245 (
            .O(N__49202),
            .I(N__49193));
    Span4Mux_h I__10244 (
            .O(N__49199),
            .I(N__49188));
    Span4Mux_v I__10243 (
            .O(N__49196),
            .I(N__49188));
    LocalMux I__10242 (
            .O(N__49193),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__10241 (
            .O(N__49188),
            .I(\c0.data_in_frame_25_3 ));
    CascadeMux I__10240 (
            .O(N__49183),
            .I(N__49179));
    CascadeMux I__10239 (
            .O(N__49182),
            .I(N__49175));
    InMux I__10238 (
            .O(N__49179),
            .I(N__49172));
    InMux I__10237 (
            .O(N__49178),
            .I(N__49169));
    InMux I__10236 (
            .O(N__49175),
            .I(N__49166));
    LocalMux I__10235 (
            .O(N__49172),
            .I(N__49161));
    LocalMux I__10234 (
            .O(N__49169),
            .I(N__49161));
    LocalMux I__10233 (
            .O(N__49166),
            .I(N__49155));
    Span4Mux_h I__10232 (
            .O(N__49161),
            .I(N__49155));
    InMux I__10231 (
            .O(N__49160),
            .I(N__49152));
    Odrv4 I__10230 (
            .O(N__49155),
            .I(\c0.n19400 ));
    LocalMux I__10229 (
            .O(N__49152),
            .I(\c0.n19400 ));
    InMux I__10228 (
            .O(N__49147),
            .I(N__49144));
    LocalMux I__10227 (
            .O(N__49144),
            .I(N__49140));
    InMux I__10226 (
            .O(N__49143),
            .I(N__49137));
    Span4Mux_h I__10225 (
            .O(N__49140),
            .I(N__49133));
    LocalMux I__10224 (
            .O(N__49137),
            .I(N__49130));
    InMux I__10223 (
            .O(N__49136),
            .I(N__49127));
    Span4Mux_v I__10222 (
            .O(N__49133),
            .I(N__49124));
    Span4Mux_h I__10221 (
            .O(N__49130),
            .I(N__49121));
    LocalMux I__10220 (
            .O(N__49127),
            .I(N__49118));
    Odrv4 I__10219 (
            .O(N__49124),
            .I(\c0.n12134 ));
    Odrv4 I__10218 (
            .O(N__49121),
            .I(\c0.n12134 ));
    Odrv12 I__10217 (
            .O(N__49118),
            .I(\c0.n12134 ));
    InMux I__10216 (
            .O(N__49111),
            .I(N__49108));
    LocalMux I__10215 (
            .O(N__49108),
            .I(\c0.n58_adj_3381 ));
    InMux I__10214 (
            .O(N__49105),
            .I(N__49102));
    LocalMux I__10213 (
            .O(N__49102),
            .I(N__49099));
    Span4Mux_v I__10212 (
            .O(N__49099),
            .I(N__49095));
    InMux I__10211 (
            .O(N__49098),
            .I(N__49092));
    Odrv4 I__10210 (
            .O(N__49095),
            .I(\c0.n43_adj_3330 ));
    LocalMux I__10209 (
            .O(N__49092),
            .I(\c0.n43_adj_3330 ));
    InMux I__10208 (
            .O(N__49087),
            .I(N__49084));
    LocalMux I__10207 (
            .O(N__49084),
            .I(\c0.n50_adj_3331 ));
    InMux I__10206 (
            .O(N__49081),
            .I(N__49076));
    InMux I__10205 (
            .O(N__49080),
            .I(N__49073));
    InMux I__10204 (
            .O(N__49079),
            .I(N__49070));
    LocalMux I__10203 (
            .O(N__49076),
            .I(N__49065));
    LocalMux I__10202 (
            .O(N__49073),
            .I(N__49062));
    LocalMux I__10201 (
            .O(N__49070),
            .I(N__49059));
    InMux I__10200 (
            .O(N__49069),
            .I(N__49056));
    InMux I__10199 (
            .O(N__49068),
            .I(N__49053));
    Span4Mux_v I__10198 (
            .O(N__49065),
            .I(N__49050));
    Span4Mux_v I__10197 (
            .O(N__49062),
            .I(N__49045));
    Span4Mux_h I__10196 (
            .O(N__49059),
            .I(N__49045));
    LocalMux I__10195 (
            .O(N__49056),
            .I(N__49040));
    LocalMux I__10194 (
            .O(N__49053),
            .I(N__49040));
    Span4Mux_h I__10193 (
            .O(N__49050),
            .I(N__49037));
    Span4Mux_v I__10192 (
            .O(N__49045),
            .I(N__49034));
    Span4Mux_h I__10191 (
            .O(N__49040),
            .I(N__49031));
    Odrv4 I__10190 (
            .O(N__49037),
            .I(\c0.n35_adj_3266 ));
    Odrv4 I__10189 (
            .O(N__49034),
            .I(\c0.n35_adj_3266 ));
    Odrv4 I__10188 (
            .O(N__49031),
            .I(\c0.n35_adj_3266 ));
    InMux I__10187 (
            .O(N__49024),
            .I(N__49021));
    LocalMux I__10186 (
            .O(N__49021),
            .I(N__49018));
    Span4Mux_v I__10185 (
            .O(N__49018),
            .I(N__49014));
    InMux I__10184 (
            .O(N__49017),
            .I(N__49011));
    Odrv4 I__10183 (
            .O(N__49014),
            .I(\c0.n33_adj_3097 ));
    LocalMux I__10182 (
            .O(N__49011),
            .I(\c0.n33_adj_3097 ));
    CascadeMux I__10181 (
            .O(N__49006),
            .I(N__49003));
    InMux I__10180 (
            .O(N__49003),
            .I(N__49000));
    LocalMux I__10179 (
            .O(N__49000),
            .I(N__48997));
    Span4Mux_v I__10178 (
            .O(N__48997),
            .I(N__48994));
    Odrv4 I__10177 (
            .O(N__48994),
            .I(\c0.n9_adj_3240 ));
    InMux I__10176 (
            .O(N__48991),
            .I(N__48988));
    LocalMux I__10175 (
            .O(N__48988),
            .I(N__48985));
    Span4Mux_v I__10174 (
            .O(N__48985),
            .I(N__48982));
    Odrv4 I__10173 (
            .O(N__48982),
            .I(\c0.n20112 ));
    InMux I__10172 (
            .O(N__48979),
            .I(N__48976));
    LocalMux I__10171 (
            .O(N__48976),
            .I(N__48973));
    Span4Mux_h I__10170 (
            .O(N__48973),
            .I(N__48970));
    Span4Mux_v I__10169 (
            .O(N__48970),
            .I(N__48967));
    Odrv4 I__10168 (
            .O(N__48967),
            .I(\c0.n32_adj_3236 ));
    InMux I__10167 (
            .O(N__48964),
            .I(N__48961));
    LocalMux I__10166 (
            .O(N__48961),
            .I(N__48957));
    InMux I__10165 (
            .O(N__48960),
            .I(N__48954));
    Span4Mux_v I__10164 (
            .O(N__48957),
            .I(N__48949));
    LocalMux I__10163 (
            .O(N__48954),
            .I(N__48949));
    Span4Mux_v I__10162 (
            .O(N__48949),
            .I(N__48946));
    Odrv4 I__10161 (
            .O(N__48946),
            .I(\c0.n28_adj_3245 ));
    CascadeMux I__10160 (
            .O(N__48943),
            .I(\c0.n27_adj_3241_cascade_ ));
    InMux I__10159 (
            .O(N__48940),
            .I(N__48937));
    LocalMux I__10158 (
            .O(N__48937),
            .I(N__48934));
    Span4Mux_v I__10157 (
            .O(N__48934),
            .I(N__48927));
    InMux I__10156 (
            .O(N__48933),
            .I(N__48924));
    InMux I__10155 (
            .O(N__48932),
            .I(N__48921));
    InMux I__10154 (
            .O(N__48931),
            .I(N__48916));
    InMux I__10153 (
            .O(N__48930),
            .I(N__48916));
    Odrv4 I__10152 (
            .O(N__48927),
            .I(\c0.n13_adj_3244 ));
    LocalMux I__10151 (
            .O(N__48924),
            .I(\c0.n13_adj_3244 ));
    LocalMux I__10150 (
            .O(N__48921),
            .I(\c0.n13_adj_3244 ));
    LocalMux I__10149 (
            .O(N__48916),
            .I(\c0.n13_adj_3244 ));
    InMux I__10148 (
            .O(N__48907),
            .I(N__48904));
    LocalMux I__10147 (
            .O(N__48904),
            .I(\c0.n19_adj_3135 ));
    CascadeMux I__10146 (
            .O(N__48901),
            .I(\c0.n19_adj_3135_cascade_ ));
    InMux I__10145 (
            .O(N__48898),
            .I(N__48895));
    LocalMux I__10144 (
            .O(N__48895),
            .I(N__48891));
    InMux I__10143 (
            .O(N__48894),
            .I(N__48888));
    Span4Mux_h I__10142 (
            .O(N__48891),
            .I(N__48885));
    LocalMux I__10141 (
            .O(N__48888),
            .I(\c0.n24_adj_3134 ));
    Odrv4 I__10140 (
            .O(N__48885),
            .I(\c0.n24_adj_3134 ));
    InMux I__10139 (
            .O(N__48880),
            .I(N__48877));
    LocalMux I__10138 (
            .O(N__48877),
            .I(N__48873));
    InMux I__10137 (
            .O(N__48876),
            .I(N__48870));
    Span4Mux_v I__10136 (
            .O(N__48873),
            .I(N__48864));
    LocalMux I__10135 (
            .O(N__48870),
            .I(N__48864));
    InMux I__10134 (
            .O(N__48869),
            .I(N__48861));
    Span4Mux_v I__10133 (
            .O(N__48864),
            .I(N__48855));
    LocalMux I__10132 (
            .O(N__48861),
            .I(N__48855));
    InMux I__10131 (
            .O(N__48860),
            .I(N__48852));
    Span4Mux_h I__10130 (
            .O(N__48855),
            .I(N__48849));
    LocalMux I__10129 (
            .O(N__48852),
            .I(\c0.n86 ));
    Odrv4 I__10128 (
            .O(N__48849),
            .I(\c0.n86 ));
    CascadeMux I__10127 (
            .O(N__48844),
            .I(\c0.n22_adj_3136_cascade_ ));
    CascadeMux I__10126 (
            .O(N__48841),
            .I(\c0.n11936_cascade_ ));
    InMux I__10125 (
            .O(N__48838),
            .I(N__48834));
    InMux I__10124 (
            .O(N__48837),
            .I(N__48831));
    LocalMux I__10123 (
            .O(N__48834),
            .I(N__48826));
    LocalMux I__10122 (
            .O(N__48831),
            .I(N__48823));
    CascadeMux I__10121 (
            .O(N__48830),
            .I(N__48820));
    InMux I__10120 (
            .O(N__48829),
            .I(N__48817));
    Span4Mux_h I__10119 (
            .O(N__48826),
            .I(N__48814));
    Span4Mux_h I__10118 (
            .O(N__48823),
            .I(N__48811));
    InMux I__10117 (
            .O(N__48820),
            .I(N__48808));
    LocalMux I__10116 (
            .O(N__48817),
            .I(N__48805));
    Span4Mux_h I__10115 (
            .O(N__48814),
            .I(N__48802));
    Span4Mux_h I__10114 (
            .O(N__48811),
            .I(N__48799));
    LocalMux I__10113 (
            .O(N__48808),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__10112 (
            .O(N__48805),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__10111 (
            .O(N__48802),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__10110 (
            .O(N__48799),
            .I(\c0.data_in_frame_27_4 ));
    InMux I__10109 (
            .O(N__48790),
            .I(N__48786));
    InMux I__10108 (
            .O(N__48789),
            .I(N__48782));
    LocalMux I__10107 (
            .O(N__48786),
            .I(N__48779));
    CascadeMux I__10106 (
            .O(N__48785),
            .I(N__48775));
    LocalMux I__10105 (
            .O(N__48782),
            .I(N__48772));
    Span4Mux_v I__10104 (
            .O(N__48779),
            .I(N__48769));
    CascadeMux I__10103 (
            .O(N__48778),
            .I(N__48766));
    InMux I__10102 (
            .O(N__48775),
            .I(N__48763));
    Span4Mux_h I__10101 (
            .O(N__48772),
            .I(N__48760));
    Sp12to4 I__10100 (
            .O(N__48769),
            .I(N__48757));
    InMux I__10099 (
            .O(N__48766),
            .I(N__48754));
    LocalMux I__10098 (
            .O(N__48763),
            .I(N__48751));
    Span4Mux_v I__10097 (
            .O(N__48760),
            .I(N__48748));
    Span12Mux_h I__10096 (
            .O(N__48757),
            .I(N__48743));
    LocalMux I__10095 (
            .O(N__48754),
            .I(N__48743));
    Odrv4 I__10094 (
            .O(N__48751),
            .I(\c0.data_in_frame_27_5 ));
    Odrv4 I__10093 (
            .O(N__48748),
            .I(\c0.data_in_frame_27_5 ));
    Odrv12 I__10092 (
            .O(N__48743),
            .I(\c0.data_in_frame_27_5 ));
    InMux I__10091 (
            .O(N__48736),
            .I(N__48733));
    LocalMux I__10090 (
            .O(N__48733),
            .I(N__48730));
    Odrv4 I__10089 (
            .O(N__48730),
            .I(\c0.n17_adj_3318 ));
    CascadeMux I__10088 (
            .O(N__48727),
            .I(\c0.n32_adj_3057_cascade_ ));
    InMux I__10087 (
            .O(N__48724),
            .I(N__48716));
    InMux I__10086 (
            .O(N__48723),
            .I(N__48716));
    InMux I__10085 (
            .O(N__48722),
            .I(N__48711));
    InMux I__10084 (
            .O(N__48721),
            .I(N__48711));
    LocalMux I__10083 (
            .O(N__48716),
            .I(N__48708));
    LocalMux I__10082 (
            .O(N__48711),
            .I(N__48703));
    Span4Mux_v I__10081 (
            .O(N__48708),
            .I(N__48703));
    Span4Mux_v I__10080 (
            .O(N__48703),
            .I(N__48700));
    Odrv4 I__10079 (
            .O(N__48700),
            .I(\c0.n33_adj_3289 ));
    InMux I__10078 (
            .O(N__48697),
            .I(N__48694));
    LocalMux I__10077 (
            .O(N__48694),
            .I(N__48691));
    Odrv4 I__10076 (
            .O(N__48691),
            .I(\c0.n10_adj_3555 ));
    CascadeMux I__10075 (
            .O(N__48688),
            .I(N__48685));
    InMux I__10074 (
            .O(N__48685),
            .I(N__48682));
    LocalMux I__10073 (
            .O(N__48682),
            .I(N__48679));
    Span4Mux_v I__10072 (
            .O(N__48679),
            .I(N__48676));
    Span4Mux_h I__10071 (
            .O(N__48676),
            .I(N__48673));
    Sp12to4 I__10070 (
            .O(N__48673),
            .I(N__48670));
    Odrv12 I__10069 (
            .O(N__48670),
            .I(\c0.n4_adj_3522 ));
    InMux I__10068 (
            .O(N__48667),
            .I(N__48661));
    InMux I__10067 (
            .O(N__48666),
            .I(N__48661));
    LocalMux I__10066 (
            .O(N__48661),
            .I(\c0.n55_adj_3273 ));
    InMux I__10065 (
            .O(N__48658),
            .I(N__48655));
    LocalMux I__10064 (
            .O(N__48655),
            .I(N__48651));
    InMux I__10063 (
            .O(N__48654),
            .I(N__48647));
    Span4Mux_v I__10062 (
            .O(N__48651),
            .I(N__48644));
    InMux I__10061 (
            .O(N__48650),
            .I(N__48641));
    LocalMux I__10060 (
            .O(N__48647),
            .I(\c0.n19514 ));
    Odrv4 I__10059 (
            .O(N__48644),
            .I(\c0.n19514 ));
    LocalMux I__10058 (
            .O(N__48641),
            .I(\c0.n19514 ));
    CascadeMux I__10057 (
            .O(N__48634),
            .I(\c0.n20965_cascade_ ));
    InMux I__10056 (
            .O(N__48631),
            .I(N__48628));
    LocalMux I__10055 (
            .O(N__48628),
            .I(N__48625));
    Span4Mux_h I__10054 (
            .O(N__48625),
            .I(N__48622));
    Odrv4 I__10053 (
            .O(N__48622),
            .I(\c0.n40_adj_3323 ));
    InMux I__10052 (
            .O(N__48619),
            .I(N__48614));
    InMux I__10051 (
            .O(N__48618),
            .I(N__48611));
    CascadeMux I__10050 (
            .O(N__48617),
            .I(N__48608));
    LocalMux I__10049 (
            .O(N__48614),
            .I(N__48605));
    LocalMux I__10048 (
            .O(N__48611),
            .I(N__48602));
    InMux I__10047 (
            .O(N__48608),
            .I(N__48599));
    Span4Mux_v I__10046 (
            .O(N__48605),
            .I(N__48596));
    Span4Mux_v I__10045 (
            .O(N__48602),
            .I(N__48592));
    LocalMux I__10044 (
            .O(N__48599),
            .I(N__48587));
    Span4Mux_v I__10043 (
            .O(N__48596),
            .I(N__48587));
    InMux I__10042 (
            .O(N__48595),
            .I(N__48584));
    Span4Mux_h I__10041 (
            .O(N__48592),
            .I(N__48581));
    Odrv4 I__10040 (
            .O(N__48587),
            .I(\c0.data_in_frame_27_3 ));
    LocalMux I__10039 (
            .O(N__48584),
            .I(\c0.data_in_frame_27_3 ));
    Odrv4 I__10038 (
            .O(N__48581),
            .I(\c0.data_in_frame_27_3 ));
    CascadeMux I__10037 (
            .O(N__48574),
            .I(\c0.n20336_cascade_ ));
    InMux I__10036 (
            .O(N__48571),
            .I(N__48568));
    LocalMux I__10035 (
            .O(N__48568),
            .I(N__48565));
    Span4Mux_v I__10034 (
            .O(N__48565),
            .I(N__48562));
    Odrv4 I__10033 (
            .O(N__48562),
            .I(\c0.n61_adj_3387 ));
    InMux I__10032 (
            .O(N__48559),
            .I(N__48556));
    LocalMux I__10031 (
            .O(N__48556),
            .I(N__48553));
    Odrv4 I__10030 (
            .O(N__48553),
            .I(\c0.n63_adj_3391 ));
    CascadeMux I__10029 (
            .O(N__48550),
            .I(\c0.n21034_cascade_ ));
    CascadeMux I__10028 (
            .O(N__48547),
            .I(\c0.n35_adj_3274_cascade_ ));
    InMux I__10027 (
            .O(N__48544),
            .I(N__48541));
    LocalMux I__10026 (
            .O(N__48541),
            .I(\c0.n59 ));
    InMux I__10025 (
            .O(N__48538),
            .I(N__48535));
    LocalMux I__10024 (
            .O(N__48535),
            .I(N__48531));
    InMux I__10023 (
            .O(N__48534),
            .I(N__48528));
    Span4Mux_h I__10022 (
            .O(N__48531),
            .I(N__48524));
    LocalMux I__10021 (
            .O(N__48528),
            .I(N__48521));
    InMux I__10020 (
            .O(N__48527),
            .I(N__48518));
    Odrv4 I__10019 (
            .O(N__48524),
            .I(\c0.n30_adj_3392 ));
    Odrv12 I__10018 (
            .O(N__48521),
            .I(\c0.n30_adj_3392 ));
    LocalMux I__10017 (
            .O(N__48518),
            .I(\c0.n30_adj_3392 ));
    InMux I__10016 (
            .O(N__48511),
            .I(N__48507));
    InMux I__10015 (
            .O(N__48510),
            .I(N__48504));
    LocalMux I__10014 (
            .O(N__48507),
            .I(N__48501));
    LocalMux I__10013 (
            .O(N__48504),
            .I(N__48496));
    Span4Mux_v I__10012 (
            .O(N__48501),
            .I(N__48496));
    Span4Mux_v I__10011 (
            .O(N__48496),
            .I(N__48493));
    Odrv4 I__10010 (
            .O(N__48493),
            .I(\c0.n21047 ));
    InMux I__10009 (
            .O(N__48490),
            .I(N__48486));
    InMux I__10008 (
            .O(N__48489),
            .I(N__48483));
    LocalMux I__10007 (
            .O(N__48486),
            .I(N__48480));
    LocalMux I__10006 (
            .O(N__48483),
            .I(N__48477));
    Span4Mux_h I__10005 (
            .O(N__48480),
            .I(N__48474));
    Span4Mux_v I__10004 (
            .O(N__48477),
            .I(N__48471));
    Sp12to4 I__10003 (
            .O(N__48474),
            .I(N__48468));
    Span4Mux_v I__10002 (
            .O(N__48471),
            .I(N__48465));
    Odrv12 I__10001 (
            .O(N__48468),
            .I(\c0.n12_adj_3049 ));
    Odrv4 I__10000 (
            .O(N__48465),
            .I(\c0.n12_adj_3049 ));
    InMux I__9999 (
            .O(N__48460),
            .I(N__48457));
    LocalMux I__9998 (
            .O(N__48457),
            .I(N__48454));
    Odrv12 I__9997 (
            .O(N__48454),
            .I(\c0.n91 ));
    CascadeMux I__9996 (
            .O(N__48451),
            .I(N__48447));
    InMux I__9995 (
            .O(N__48450),
            .I(N__48444));
    InMux I__9994 (
            .O(N__48447),
            .I(N__48441));
    LocalMux I__9993 (
            .O(N__48444),
            .I(\c0.n35_adj_3274 ));
    LocalMux I__9992 (
            .O(N__48441),
            .I(\c0.n35_adj_3274 ));
    InMux I__9991 (
            .O(N__48436),
            .I(N__48433));
    LocalMux I__9990 (
            .O(N__48433),
            .I(N__48430));
    Span4Mux_v I__9989 (
            .O(N__48430),
            .I(N__48426));
    InMux I__9988 (
            .O(N__48429),
            .I(N__48423));
    Span4Mux_h I__9987 (
            .O(N__48426),
            .I(N__48420));
    LocalMux I__9986 (
            .O(N__48423),
            .I(N__48417));
    Odrv4 I__9985 (
            .O(N__48420),
            .I(\c0.n17_adj_3451 ));
    Odrv4 I__9984 (
            .O(N__48417),
            .I(\c0.n17_adj_3451 ));
    InMux I__9983 (
            .O(N__48412),
            .I(N__48409));
    LocalMux I__9982 (
            .O(N__48409),
            .I(N__48406));
    Span4Mux_v I__9981 (
            .O(N__48406),
            .I(N__48403));
    Span4Mux_h I__9980 (
            .O(N__48403),
            .I(N__48399));
    InMux I__9979 (
            .O(N__48402),
            .I(N__48396));
    Odrv4 I__9978 (
            .O(N__48399),
            .I(\c0.n20403 ));
    LocalMux I__9977 (
            .O(N__48396),
            .I(\c0.n20403 ));
    InMux I__9976 (
            .O(N__48391),
            .I(N__48388));
    LocalMux I__9975 (
            .O(N__48388),
            .I(\c0.n22_adj_3450 ));
    CascadeMux I__9974 (
            .O(N__48385),
            .I(\c0.n24_adj_3427_cascade_ ));
    InMux I__9973 (
            .O(N__48382),
            .I(N__48378));
    InMux I__9972 (
            .O(N__48381),
            .I(N__48374));
    LocalMux I__9971 (
            .O(N__48378),
            .I(N__48370));
    InMux I__9970 (
            .O(N__48377),
            .I(N__48367));
    LocalMux I__9969 (
            .O(N__48374),
            .I(N__48363));
    InMux I__9968 (
            .O(N__48373),
            .I(N__48360));
    Span4Mux_v I__9967 (
            .O(N__48370),
            .I(N__48355));
    LocalMux I__9966 (
            .O(N__48367),
            .I(N__48355));
    CascadeMux I__9965 (
            .O(N__48366),
            .I(N__48352));
    Span4Mux_v I__9964 (
            .O(N__48363),
            .I(N__48345));
    LocalMux I__9963 (
            .O(N__48360),
            .I(N__48345));
    Span4Mux_h I__9962 (
            .O(N__48355),
            .I(N__48345));
    InMux I__9961 (
            .O(N__48352),
            .I(N__48342));
    Span4Mux_v I__9960 (
            .O(N__48345),
            .I(N__48339));
    LocalMux I__9959 (
            .O(N__48342),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__9958 (
            .O(N__48339),
            .I(\c0.data_in_frame_17_0 ));
    InMux I__9957 (
            .O(N__48334),
            .I(N__48330));
    InMux I__9956 (
            .O(N__48333),
            .I(N__48327));
    LocalMux I__9955 (
            .O(N__48330),
            .I(N__48322));
    LocalMux I__9954 (
            .O(N__48327),
            .I(N__48319));
    InMux I__9953 (
            .O(N__48326),
            .I(N__48314));
    InMux I__9952 (
            .O(N__48325),
            .I(N__48314));
    Span12Mux_v I__9951 (
            .O(N__48322),
            .I(N__48311));
    Odrv4 I__9950 (
            .O(N__48319),
            .I(\c0.data_in_frame_13_1 ));
    LocalMux I__9949 (
            .O(N__48314),
            .I(\c0.data_in_frame_13_1 ));
    Odrv12 I__9948 (
            .O(N__48311),
            .I(\c0.data_in_frame_13_1 ));
    CascadeMux I__9947 (
            .O(N__48304),
            .I(\c0.n18398_cascade_ ));
    CascadeMux I__9946 (
            .O(N__48301),
            .I(\c0.n37_adj_3390_cascade_ ));
    InMux I__9945 (
            .O(N__48298),
            .I(N__48295));
    LocalMux I__9944 (
            .O(N__48295),
            .I(\c0.n37_adj_3390 ));
    CascadeMux I__9943 (
            .O(N__48292),
            .I(\c0.n60_adj_3368_cascade_ ));
    InMux I__9942 (
            .O(N__48289),
            .I(N__48286));
    LocalMux I__9941 (
            .O(N__48286),
            .I(\c0.n51_adj_3376 ));
    InMux I__9940 (
            .O(N__48283),
            .I(N__48280));
    LocalMux I__9939 (
            .O(N__48280),
            .I(N__48276));
    InMux I__9938 (
            .O(N__48279),
            .I(N__48273));
    Span4Mux_v I__9937 (
            .O(N__48276),
            .I(N__48270));
    LocalMux I__9936 (
            .O(N__48273),
            .I(\c0.n19916 ));
    Odrv4 I__9935 (
            .O(N__48270),
            .I(\c0.n19916 ));
    InMux I__9934 (
            .O(N__48265),
            .I(N__48262));
    LocalMux I__9933 (
            .O(N__48262),
            .I(N__48257));
    InMux I__9932 (
            .O(N__48261),
            .I(N__48254));
    InMux I__9931 (
            .O(N__48260),
            .I(N__48251));
    Span4Mux_h I__9930 (
            .O(N__48257),
            .I(N__48248));
    LocalMux I__9929 (
            .O(N__48254),
            .I(N__48243));
    LocalMux I__9928 (
            .O(N__48251),
            .I(N__48243));
    Span4Mux_v I__9927 (
            .O(N__48248),
            .I(N__48240));
    Span4Mux_v I__9926 (
            .O(N__48243),
            .I(N__48237));
    Odrv4 I__9925 (
            .O(N__48240),
            .I(\c0.n18443 ));
    Odrv4 I__9924 (
            .O(N__48237),
            .I(\c0.n18443 ));
    InMux I__9923 (
            .O(N__48232),
            .I(N__48229));
    LocalMux I__9922 (
            .O(N__48229),
            .I(\c0.n39_adj_3334 ));
    InMux I__9921 (
            .O(N__48226),
            .I(N__48220));
    InMux I__9920 (
            .O(N__48225),
            .I(N__48220));
    LocalMux I__9919 (
            .O(N__48220),
            .I(N__48216));
    CascadeMux I__9918 (
            .O(N__48219),
            .I(N__48213));
    Span4Mux_v I__9917 (
            .O(N__48216),
            .I(N__48210));
    InMux I__9916 (
            .O(N__48213),
            .I(N__48207));
    Odrv4 I__9915 (
            .O(N__48210),
            .I(\c0.n19_adj_3336 ));
    LocalMux I__9914 (
            .O(N__48207),
            .I(\c0.n19_adj_3336 ));
    CascadeMux I__9913 (
            .O(N__48202),
            .I(\c0.n39_adj_3334_cascade_ ));
    InMux I__9912 (
            .O(N__48199),
            .I(N__48196));
    LocalMux I__9911 (
            .O(N__48196),
            .I(\c0.n25_adj_3431 ));
    InMux I__9910 (
            .O(N__48193),
            .I(N__48187));
    InMux I__9909 (
            .O(N__48192),
            .I(N__48187));
    LocalMux I__9908 (
            .O(N__48187),
            .I(N__48184));
    Odrv12 I__9907 (
            .O(N__48184),
            .I(\c0.n42_adj_3367 ));
    InMux I__9906 (
            .O(N__48181),
            .I(N__48178));
    LocalMux I__9905 (
            .O(N__48178),
            .I(N__48174));
    InMux I__9904 (
            .O(N__48177),
            .I(N__48171));
    Span4Mux_v I__9903 (
            .O(N__48174),
            .I(N__48168));
    LocalMux I__9902 (
            .O(N__48171),
            .I(\c0.n43_adj_3386 ));
    Odrv4 I__9901 (
            .O(N__48168),
            .I(\c0.n43_adj_3386 ));
    InMux I__9900 (
            .O(N__48163),
            .I(N__48157));
    InMux I__9899 (
            .O(N__48162),
            .I(N__48157));
    LocalMux I__9898 (
            .O(N__48157),
            .I(N__48154));
    Span4Mux_v I__9897 (
            .O(N__48154),
            .I(N__48151));
    Span4Mux_h I__9896 (
            .O(N__48151),
            .I(N__48148));
    Odrv4 I__9895 (
            .O(N__48148),
            .I(\c0.n40_adj_3366 ));
    InMux I__9894 (
            .O(N__48145),
            .I(N__48142));
    LocalMux I__9893 (
            .O(N__48142),
            .I(\c0.n30_adj_3429 ));
    InMux I__9892 (
            .O(N__48139),
            .I(N__48136));
    LocalMux I__9891 (
            .O(N__48136),
            .I(\c0.n46 ));
    InMux I__9890 (
            .O(N__48133),
            .I(N__48127));
    InMux I__9889 (
            .O(N__48132),
            .I(N__48120));
    InMux I__9888 (
            .O(N__48131),
            .I(N__48120));
    InMux I__9887 (
            .O(N__48130),
            .I(N__48120));
    LocalMux I__9886 (
            .O(N__48127),
            .I(N__48117));
    LocalMux I__9885 (
            .O(N__48120),
            .I(N__48114));
    Span4Mux_v I__9884 (
            .O(N__48117),
            .I(N__48111));
    Span4Mux_h I__9883 (
            .O(N__48114),
            .I(N__48108));
    Odrv4 I__9882 (
            .O(N__48111),
            .I(\c0.n8 ));
    Odrv4 I__9881 (
            .O(N__48108),
            .I(\c0.n8 ));
    InMux I__9880 (
            .O(N__48103),
            .I(N__48099));
    CascadeMux I__9879 (
            .O(N__48102),
            .I(N__48096));
    LocalMux I__9878 (
            .O(N__48099),
            .I(N__48093));
    InMux I__9877 (
            .O(N__48096),
            .I(N__48090));
    Odrv12 I__9876 (
            .O(N__48093),
            .I(\c0.n84 ));
    LocalMux I__9875 (
            .O(N__48090),
            .I(\c0.n84 ));
    CascadeMux I__9874 (
            .O(N__48085),
            .I(\c0.n19824_cascade_ ));
    InMux I__9873 (
            .O(N__48082),
            .I(N__48078));
    InMux I__9872 (
            .O(N__48081),
            .I(N__48075));
    LocalMux I__9871 (
            .O(N__48078),
            .I(N__48072));
    LocalMux I__9870 (
            .O(N__48075),
            .I(N__48069));
    Span4Mux_h I__9869 (
            .O(N__48072),
            .I(N__48065));
    Span4Mux_v I__9868 (
            .O(N__48069),
            .I(N__48062));
    InMux I__9867 (
            .O(N__48068),
            .I(N__48059));
    Odrv4 I__9866 (
            .O(N__48065),
            .I(\c0.n29 ));
    Odrv4 I__9865 (
            .O(N__48062),
            .I(\c0.n29 ));
    LocalMux I__9864 (
            .O(N__48059),
            .I(\c0.n29 ));
    CascadeMux I__9863 (
            .O(N__48052),
            .I(\c0.n18_adj_3360_cascade_ ));
    CascadeMux I__9862 (
            .O(N__48049),
            .I(\c0.n32_adj_3362_cascade_ ));
    CascadeMux I__9861 (
            .O(N__48046),
            .I(\c0.n20112_cascade_ ));
    CascadeMux I__9860 (
            .O(N__48043),
            .I(\c0.n12_adj_3249_cascade_ ));
    InMux I__9859 (
            .O(N__48040),
            .I(N__48037));
    LocalMux I__9858 (
            .O(N__48037),
            .I(\c0.n12056 ));
    InMux I__9857 (
            .O(N__48034),
            .I(N__48027));
    InMux I__9856 (
            .O(N__48033),
            .I(N__48027));
    CascadeMux I__9855 (
            .O(N__48032),
            .I(N__48024));
    LocalMux I__9854 (
            .O(N__48027),
            .I(N__48021));
    InMux I__9853 (
            .O(N__48024),
            .I(N__48018));
    Sp12to4 I__9852 (
            .O(N__48021),
            .I(N__48015));
    LocalMux I__9851 (
            .O(N__48018),
            .I(N__48012));
    Odrv12 I__9850 (
            .O(N__48015),
            .I(\c0.n19301 ));
    Odrv12 I__9849 (
            .O(N__48012),
            .I(\c0.n19301 ));
    CascadeMux I__9848 (
            .O(N__48007),
            .I(\c0.n19301_cascade_ ));
    CascadeMux I__9847 (
            .O(N__48004),
            .I(\c0.n31_adj_3126_cascade_ ));
    CascadeMux I__9846 (
            .O(N__48001),
            .I(N__47997));
    CascadeMux I__9845 (
            .O(N__48000),
            .I(N__47994));
    InMux I__9844 (
            .O(N__47997),
            .I(N__47989));
    InMux I__9843 (
            .O(N__47994),
            .I(N__47989));
    LocalMux I__9842 (
            .O(N__47989),
            .I(N__47986));
    Span4Mux_h I__9841 (
            .O(N__47986),
            .I(N__47983));
    Odrv4 I__9840 (
            .O(N__47983),
            .I(\c0.n19427 ));
    InMux I__9839 (
            .O(N__47980),
            .I(N__47977));
    LocalMux I__9838 (
            .O(N__47977),
            .I(N__47972));
    InMux I__9837 (
            .O(N__47976),
            .I(N__47967));
    InMux I__9836 (
            .O(N__47975),
            .I(N__47967));
    Span4Mux_h I__9835 (
            .O(N__47972),
            .I(N__47964));
    LocalMux I__9834 (
            .O(N__47967),
            .I(N__47961));
    Odrv4 I__9833 (
            .O(N__47964),
            .I(\c0.n19551 ));
    Odrv12 I__9832 (
            .O(N__47961),
            .I(\c0.n19551 ));
    InMux I__9831 (
            .O(N__47956),
            .I(N__47953));
    LocalMux I__9830 (
            .O(N__47953),
            .I(N__47950));
    Span4Mux_h I__9829 (
            .O(N__47950),
            .I(N__47947));
    Odrv4 I__9828 (
            .O(N__47947),
            .I(\c0.n27_adj_3455 ));
    CascadeMux I__9827 (
            .O(N__47944),
            .I(\c0.n46_cascade_ ));
    InMux I__9826 (
            .O(N__47941),
            .I(N__47938));
    LocalMux I__9825 (
            .O(N__47938),
            .I(N__47935));
    Span4Mux_h I__9824 (
            .O(N__47935),
            .I(N__47932));
    Span4Mux_v I__9823 (
            .O(N__47932),
            .I(N__47929));
    Odrv4 I__9822 (
            .O(N__47929),
            .I(\c0.n31_adj_3532 ));
    InMux I__9821 (
            .O(N__47926),
            .I(N__47922));
    InMux I__9820 (
            .O(N__47925),
            .I(N__47918));
    LocalMux I__9819 (
            .O(N__47922),
            .I(N__47915));
    InMux I__9818 (
            .O(N__47921),
            .I(N__47912));
    LocalMux I__9817 (
            .O(N__47918),
            .I(N__47908));
    Span4Mux_v I__9816 (
            .O(N__47915),
            .I(N__47903));
    LocalMux I__9815 (
            .O(N__47912),
            .I(N__47903));
    InMux I__9814 (
            .O(N__47911),
            .I(N__47900));
    Span4Mux_v I__9813 (
            .O(N__47908),
            .I(N__47897));
    Span4Mux_h I__9812 (
            .O(N__47903),
            .I(N__47894));
    LocalMux I__9811 (
            .O(N__47900),
            .I(\c0.n11537 ));
    Odrv4 I__9810 (
            .O(N__47897),
            .I(\c0.n11537 ));
    Odrv4 I__9809 (
            .O(N__47894),
            .I(\c0.n11537 ));
    InMux I__9808 (
            .O(N__47887),
            .I(N__47882));
    CascadeMux I__9807 (
            .O(N__47886),
            .I(N__47879));
    InMux I__9806 (
            .O(N__47885),
            .I(N__47876));
    LocalMux I__9805 (
            .O(N__47882),
            .I(N__47873));
    InMux I__9804 (
            .O(N__47879),
            .I(N__47870));
    LocalMux I__9803 (
            .O(N__47876),
            .I(N__47867));
    Span12Mux_h I__9802 (
            .O(N__47873),
            .I(N__47864));
    LocalMux I__9801 (
            .O(N__47870),
            .I(\c0.data_in_frame_15_6 ));
    Odrv4 I__9800 (
            .O(N__47867),
            .I(\c0.data_in_frame_15_6 ));
    Odrv12 I__9799 (
            .O(N__47864),
            .I(\c0.data_in_frame_15_6 ));
    CascadeMux I__9798 (
            .O(N__47857),
            .I(\c0.n16_adj_3481_cascade_ ));
    CascadeMux I__9797 (
            .O(N__47854),
            .I(\c0.n11815_cascade_ ));
    InMux I__9796 (
            .O(N__47851),
            .I(N__47845));
    InMux I__9795 (
            .O(N__47850),
            .I(N__47845));
    LocalMux I__9794 (
            .O(N__47845),
            .I(N__47842));
    Span12Mux_v I__9793 (
            .O(N__47842),
            .I(N__47839));
    Odrv12 I__9792 (
            .O(N__47839),
            .I(\c0.n19291 ));
    CascadeMux I__9791 (
            .O(N__47836),
            .I(N__47831));
    InMux I__9790 (
            .O(N__47835),
            .I(N__47827));
    InMux I__9789 (
            .O(N__47834),
            .I(N__47824));
    InMux I__9788 (
            .O(N__47831),
            .I(N__47821));
    InMux I__9787 (
            .O(N__47830),
            .I(N__47818));
    LocalMux I__9786 (
            .O(N__47827),
            .I(N__47815));
    LocalMux I__9785 (
            .O(N__47824),
            .I(N__47812));
    LocalMux I__9784 (
            .O(N__47821),
            .I(N__47809));
    LocalMux I__9783 (
            .O(N__47818),
            .I(N__47804));
    Span4Mux_h I__9782 (
            .O(N__47815),
            .I(N__47804));
    Span4Mux_v I__9781 (
            .O(N__47812),
            .I(N__47799));
    Span4Mux_v I__9780 (
            .O(N__47809),
            .I(N__47794));
    Span4Mux_v I__9779 (
            .O(N__47804),
            .I(N__47794));
    InMux I__9778 (
            .O(N__47803),
            .I(N__47789));
    InMux I__9777 (
            .O(N__47802),
            .I(N__47789));
    Odrv4 I__9776 (
            .O(N__47799),
            .I(data_in_frame_16_1));
    Odrv4 I__9775 (
            .O(N__47794),
            .I(data_in_frame_16_1));
    LocalMux I__9774 (
            .O(N__47789),
            .I(data_in_frame_16_1));
    CascadeMux I__9773 (
            .O(N__47782),
            .I(\c0.n12056_cascade_ ));
    InMux I__9772 (
            .O(N__47779),
            .I(N__47776));
    LocalMux I__9771 (
            .O(N__47776),
            .I(\c0.n12_adj_3249 ));
    InMux I__9770 (
            .O(N__47773),
            .I(N__47769));
    InMux I__9769 (
            .O(N__47772),
            .I(N__47764));
    LocalMux I__9768 (
            .O(N__47769),
            .I(N__47761));
    InMux I__9767 (
            .O(N__47768),
            .I(N__47758));
    CascadeMux I__9766 (
            .O(N__47767),
            .I(N__47755));
    LocalMux I__9765 (
            .O(N__47764),
            .I(N__47752));
    Span4Mux_v I__9764 (
            .O(N__47761),
            .I(N__47749));
    LocalMux I__9763 (
            .O(N__47758),
            .I(N__47746));
    InMux I__9762 (
            .O(N__47755),
            .I(N__47742));
    Span4Mux_v I__9761 (
            .O(N__47752),
            .I(N__47739));
    Span4Mux_h I__9760 (
            .O(N__47749),
            .I(N__47734));
    Span4Mux_v I__9759 (
            .O(N__47746),
            .I(N__47734));
    InMux I__9758 (
            .O(N__47745),
            .I(N__47731));
    LocalMux I__9757 (
            .O(N__47742),
            .I(\c0.data_in_frame_12_2 ));
    Odrv4 I__9756 (
            .O(N__47739),
            .I(\c0.data_in_frame_12_2 ));
    Odrv4 I__9755 (
            .O(N__47734),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__9754 (
            .O(N__47731),
            .I(\c0.data_in_frame_12_2 ));
    InMux I__9753 (
            .O(N__47722),
            .I(N__47719));
    LocalMux I__9752 (
            .O(N__47719),
            .I(N__47716));
    Span4Mux_v I__9751 (
            .O(N__47716),
            .I(N__47712));
    InMux I__9750 (
            .O(N__47715),
            .I(N__47709));
    Odrv4 I__9749 (
            .O(N__47712),
            .I(\c0.n7_adj_3491 ));
    LocalMux I__9748 (
            .O(N__47709),
            .I(\c0.n7_adj_3491 ));
    InMux I__9747 (
            .O(N__47704),
            .I(N__47701));
    LocalMux I__9746 (
            .O(N__47701),
            .I(N__47698));
    Span4Mux_v I__9745 (
            .O(N__47698),
            .I(N__47695));
    Odrv4 I__9744 (
            .O(N__47695),
            .I(\c0.n30_adj_3531 ));
    InMux I__9743 (
            .O(N__47692),
            .I(N__47689));
    LocalMux I__9742 (
            .O(N__47689),
            .I(N__47685));
    InMux I__9741 (
            .O(N__47688),
            .I(N__47681));
    Span4Mux_v I__9740 (
            .O(N__47685),
            .I(N__47678));
    InMux I__9739 (
            .O(N__47684),
            .I(N__47675));
    LocalMux I__9738 (
            .O(N__47681),
            .I(N__47670));
    Span4Mux_h I__9737 (
            .O(N__47678),
            .I(N__47670));
    LocalMux I__9736 (
            .O(N__47675),
            .I(N__47667));
    Span4Mux_v I__9735 (
            .O(N__47670),
            .I(N__47664));
    Span4Mux_v I__9734 (
            .O(N__47667),
            .I(N__47661));
    Odrv4 I__9733 (
            .O(N__47664),
            .I(\c0.n12_adj_3034 ));
    Odrv4 I__9732 (
            .O(N__47661),
            .I(\c0.n12_adj_3034 ));
    CascadeMux I__9731 (
            .O(N__47656),
            .I(\c0.n32_adj_3077_cascade_ ));
    CascadeMux I__9730 (
            .O(N__47653),
            .I(N__47650));
    InMux I__9729 (
            .O(N__47650),
            .I(N__47647));
    LocalMux I__9728 (
            .O(N__47647),
            .I(N__47643));
    InMux I__9727 (
            .O(N__47646),
            .I(N__47640));
    Span4Mux_h I__9726 (
            .O(N__47643),
            .I(N__47635));
    LocalMux I__9725 (
            .O(N__47640),
            .I(N__47635));
    Odrv4 I__9724 (
            .O(N__47635),
            .I(\c0.n19372 ));
    CascadeMux I__9723 (
            .O(N__47632),
            .I(\c0.n21047_cascade_ ));
    InMux I__9722 (
            .O(N__47629),
            .I(N__47626));
    LocalMux I__9721 (
            .O(N__47626),
            .I(N__47623));
    Odrv4 I__9720 (
            .O(N__47623),
            .I(\c0.n42_adj_3111 ));
    InMux I__9719 (
            .O(N__47620),
            .I(N__47616));
    CascadeMux I__9718 (
            .O(N__47619),
            .I(N__47611));
    LocalMux I__9717 (
            .O(N__47616),
            .I(N__47608));
    InMux I__9716 (
            .O(N__47615),
            .I(N__47605));
    InMux I__9715 (
            .O(N__47614),
            .I(N__47602));
    InMux I__9714 (
            .O(N__47611),
            .I(N__47599));
    Span4Mux_v I__9713 (
            .O(N__47608),
            .I(N__47593));
    LocalMux I__9712 (
            .O(N__47605),
            .I(N__47588));
    LocalMux I__9711 (
            .O(N__47602),
            .I(N__47588));
    LocalMux I__9710 (
            .O(N__47599),
            .I(N__47585));
    InMux I__9709 (
            .O(N__47598),
            .I(N__47582));
    InMux I__9708 (
            .O(N__47597),
            .I(N__47577));
    InMux I__9707 (
            .O(N__47596),
            .I(N__47577));
    Span4Mux_h I__9706 (
            .O(N__47593),
            .I(N__47572));
    Span4Mux_v I__9705 (
            .O(N__47588),
            .I(N__47572));
    Span4Mux_v I__9704 (
            .O(N__47585),
            .I(N__47569));
    LocalMux I__9703 (
            .O(N__47582),
            .I(\c0.data_in_frame_3_0 ));
    LocalMux I__9702 (
            .O(N__47577),
            .I(\c0.data_in_frame_3_0 ));
    Odrv4 I__9701 (
            .O(N__47572),
            .I(\c0.data_in_frame_3_0 ));
    Odrv4 I__9700 (
            .O(N__47569),
            .I(\c0.data_in_frame_3_0 ));
    InMux I__9699 (
            .O(N__47560),
            .I(N__47556));
    CascadeMux I__9698 (
            .O(N__47559),
            .I(N__47552));
    LocalMux I__9697 (
            .O(N__47556),
            .I(N__47549));
    InMux I__9696 (
            .O(N__47555),
            .I(N__47542));
    InMux I__9695 (
            .O(N__47552),
            .I(N__47539));
    Span4Mux_h I__9694 (
            .O(N__47549),
            .I(N__47536));
    InMux I__9693 (
            .O(N__47548),
            .I(N__47531));
    InMux I__9692 (
            .O(N__47547),
            .I(N__47531));
    InMux I__9691 (
            .O(N__47546),
            .I(N__47526));
    InMux I__9690 (
            .O(N__47545),
            .I(N__47526));
    LocalMux I__9689 (
            .O(N__47542),
            .I(N__47521));
    LocalMux I__9688 (
            .O(N__47539),
            .I(N__47521));
    Odrv4 I__9687 (
            .O(N__47536),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__9686 (
            .O(N__47531),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__9685 (
            .O(N__47526),
            .I(\c0.data_in_frame_2_6 ));
    Odrv12 I__9684 (
            .O(N__47521),
            .I(\c0.data_in_frame_2_6 ));
    CascadeMux I__9683 (
            .O(N__47512),
            .I(\c0.n10_adj_3014_cascade_ ));
    InMux I__9682 (
            .O(N__47509),
            .I(N__47505));
    CascadeMux I__9681 (
            .O(N__47508),
            .I(N__47502));
    LocalMux I__9680 (
            .O(N__47505),
            .I(N__47499));
    InMux I__9679 (
            .O(N__47502),
            .I(N__47496));
    Span4Mux_h I__9678 (
            .O(N__47499),
            .I(N__47491));
    LocalMux I__9677 (
            .O(N__47496),
            .I(N__47491));
    Span4Mux_v I__9676 (
            .O(N__47491),
            .I(N__47487));
    InMux I__9675 (
            .O(N__47490),
            .I(N__47484));
    Odrv4 I__9674 (
            .O(N__47487),
            .I(\c0.n40 ));
    LocalMux I__9673 (
            .O(N__47484),
            .I(\c0.n40 ));
    CascadeMux I__9672 (
            .O(N__47479),
            .I(\c0.n16_adj_3218_cascade_ ));
    InMux I__9671 (
            .O(N__47476),
            .I(N__47473));
    LocalMux I__9670 (
            .O(N__47473),
            .I(\c0.n10_adj_3538 ));
    InMux I__9669 (
            .O(N__47470),
            .I(N__47467));
    LocalMux I__9668 (
            .O(N__47467),
            .I(N__47464));
    Odrv12 I__9667 (
            .O(N__47464),
            .I(\c0.n85 ));
    InMux I__9666 (
            .O(N__47461),
            .I(N__47458));
    LocalMux I__9665 (
            .O(N__47458),
            .I(N__47455));
    Span4Mux_h I__9664 (
            .O(N__47455),
            .I(N__47451));
    InMux I__9663 (
            .O(N__47454),
            .I(N__47448));
    Odrv4 I__9662 (
            .O(N__47451),
            .I(\c0.n37 ));
    LocalMux I__9661 (
            .O(N__47448),
            .I(\c0.n37 ));
    CascadeMux I__9660 (
            .O(N__47443),
            .I(\c0.n67_cascade_ ));
    InMux I__9659 (
            .O(N__47440),
            .I(N__47437));
    LocalMux I__9658 (
            .O(N__47437),
            .I(\c0.n96 ));
    InMux I__9657 (
            .O(N__47434),
            .I(N__47431));
    LocalMux I__9656 (
            .O(N__47431),
            .I(\c0.n83 ));
    InMux I__9655 (
            .O(N__47428),
            .I(N__47425));
    LocalMux I__9654 (
            .O(N__47425),
            .I(N__47421));
    InMux I__9653 (
            .O(N__47424),
            .I(N__47418));
    Span4Mux_v I__9652 (
            .O(N__47421),
            .I(N__47413));
    LocalMux I__9651 (
            .O(N__47418),
            .I(N__47413));
    Span4Mux_h I__9650 (
            .O(N__47413),
            .I(N__47410));
    Odrv4 I__9649 (
            .O(N__47410),
            .I(\c0.n40_adj_3032 ));
    CascadeMux I__9648 (
            .O(N__47407),
            .I(\c0.n100_cascade_ ));
    CascadeMux I__9647 (
            .O(N__47404),
            .I(N__47401));
    InMux I__9646 (
            .O(N__47401),
            .I(N__47398));
    LocalMux I__9645 (
            .O(N__47398),
            .I(\c0.n102 ));
    InMux I__9644 (
            .O(N__47395),
            .I(N__47392));
    LocalMux I__9643 (
            .O(N__47392),
            .I(N__47388));
    InMux I__9642 (
            .O(N__47391),
            .I(N__47385));
    Span4Mux_h I__9641 (
            .O(N__47388),
            .I(N__47382));
    LocalMux I__9640 (
            .O(N__47385),
            .I(N__47379));
    Odrv4 I__9639 (
            .O(N__47382),
            .I(\c0.n4_adj_3009 ));
    Odrv12 I__9638 (
            .O(N__47379),
            .I(\c0.n4_adj_3009 ));
    InMux I__9637 (
            .O(N__47374),
            .I(N__47371));
    LocalMux I__9636 (
            .O(N__47371),
            .I(N__47366));
    InMux I__9635 (
            .O(N__47370),
            .I(N__47361));
    InMux I__9634 (
            .O(N__47369),
            .I(N__47361));
    Odrv4 I__9633 (
            .O(N__47366),
            .I(\c0.n21_adj_3010 ));
    LocalMux I__9632 (
            .O(N__47361),
            .I(\c0.n21_adj_3010 ));
    InMux I__9631 (
            .O(N__47356),
            .I(N__47353));
    LocalMux I__9630 (
            .O(N__47353),
            .I(\c0.n28_adj_3023 ));
    InMux I__9629 (
            .O(N__47350),
            .I(N__47347));
    LocalMux I__9628 (
            .O(N__47347),
            .I(\c0.n17_adj_3508 ));
    CascadeMux I__9627 (
            .O(N__47344),
            .I(N__47341));
    InMux I__9626 (
            .O(N__47341),
            .I(N__47337));
    InMux I__9625 (
            .O(N__47340),
            .I(N__47333));
    LocalMux I__9624 (
            .O(N__47337),
            .I(N__47330));
    InMux I__9623 (
            .O(N__47336),
            .I(N__47327));
    LocalMux I__9622 (
            .O(N__47333),
            .I(N__47322));
    Span4Mux_h I__9621 (
            .O(N__47330),
            .I(N__47322));
    LocalMux I__9620 (
            .O(N__47327),
            .I(\c0.n19966 ));
    Odrv4 I__9619 (
            .O(N__47322),
            .I(\c0.n19966 ));
    InMux I__9618 (
            .O(N__47317),
            .I(N__47314));
    LocalMux I__9617 (
            .O(N__47314),
            .I(\c0.n30_adj_3075 ));
    InMux I__9616 (
            .O(N__47311),
            .I(N__47308));
    LocalMux I__9615 (
            .O(N__47308),
            .I(N__47305));
    Span4Mux_v I__9614 (
            .O(N__47305),
            .I(N__47302));
    Odrv4 I__9613 (
            .O(N__47302),
            .I(\c0.n21277 ));
    InMux I__9612 (
            .O(N__47299),
            .I(N__47289));
    InMux I__9611 (
            .O(N__47298),
            .I(N__47289));
    InMux I__9610 (
            .O(N__47297),
            .I(N__47289));
    InMux I__9609 (
            .O(N__47296),
            .I(N__47286));
    LocalMux I__9608 (
            .O(N__47289),
            .I(\c0.n4_adj_3406 ));
    LocalMux I__9607 (
            .O(N__47286),
            .I(\c0.n4_adj_3406 ));
    CascadeMux I__9606 (
            .O(N__47281),
            .I(\c0.n14_adj_3476_cascade_ ));
    CascadeMux I__9605 (
            .O(N__47278),
            .I(N__47275));
    InMux I__9604 (
            .O(N__47275),
            .I(N__47271));
    InMux I__9603 (
            .O(N__47274),
            .I(N__47266));
    LocalMux I__9602 (
            .O(N__47271),
            .I(N__47263));
    InMux I__9601 (
            .O(N__47270),
            .I(N__47260));
    CascadeMux I__9600 (
            .O(N__47269),
            .I(N__47256));
    LocalMux I__9599 (
            .O(N__47266),
            .I(N__47252));
    Span4Mux_v I__9598 (
            .O(N__47263),
            .I(N__47247));
    LocalMux I__9597 (
            .O(N__47260),
            .I(N__47247));
    InMux I__9596 (
            .O(N__47259),
            .I(N__47244));
    InMux I__9595 (
            .O(N__47256),
            .I(N__47239));
    InMux I__9594 (
            .O(N__47255),
            .I(N__47239));
    Span4Mux_v I__9593 (
            .O(N__47252),
            .I(N__47236));
    Odrv4 I__9592 (
            .O(N__47247),
            .I(\c0.data_in_frame_7_3 ));
    LocalMux I__9591 (
            .O(N__47244),
            .I(\c0.data_in_frame_7_3 ));
    LocalMux I__9590 (
            .O(N__47239),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__9589 (
            .O(N__47236),
            .I(\c0.data_in_frame_7_3 ));
    InMux I__9588 (
            .O(N__47227),
            .I(N__47224));
    LocalMux I__9587 (
            .O(N__47224),
            .I(\c0.n19508 ));
    InMux I__9586 (
            .O(N__47221),
            .I(N__47218));
    LocalMux I__9585 (
            .O(N__47218),
            .I(N__47213));
    InMux I__9584 (
            .O(N__47217),
            .I(N__47210));
    CascadeMux I__9583 (
            .O(N__47216),
            .I(N__47207));
    Span4Mux_h I__9582 (
            .O(N__47213),
            .I(N__47200));
    LocalMux I__9581 (
            .O(N__47210),
            .I(N__47200));
    InMux I__9580 (
            .O(N__47207),
            .I(N__47197));
    InMux I__9579 (
            .O(N__47206),
            .I(N__47192));
    InMux I__9578 (
            .O(N__47205),
            .I(N__47192));
    Span4Mux_v I__9577 (
            .O(N__47200),
            .I(N__47189));
    LocalMux I__9576 (
            .O(N__47197),
            .I(\c0.data_in_frame_2_0 ));
    LocalMux I__9575 (
            .O(N__47192),
            .I(\c0.data_in_frame_2_0 ));
    Odrv4 I__9574 (
            .O(N__47189),
            .I(\c0.data_in_frame_2_0 ));
    CascadeMux I__9573 (
            .O(N__47182),
            .I(N__47179));
    InMux I__9572 (
            .O(N__47179),
            .I(N__47176));
    LocalMux I__9571 (
            .O(N__47176),
            .I(\c0.n8_adj_3397 ));
    CascadeMux I__9570 (
            .O(N__47173),
            .I(\c0.n11833_cascade_ ));
    CascadeMux I__9569 (
            .O(N__47170),
            .I(\c0.n92_cascade_ ));
    InMux I__9568 (
            .O(N__47167),
            .I(N__47164));
    LocalMux I__9567 (
            .O(N__47164),
            .I(\c0.n80 ));
    InMux I__9566 (
            .O(N__47161),
            .I(N__47158));
    LocalMux I__9565 (
            .O(N__47158),
            .I(\c0.n19196 ));
    CascadeMux I__9564 (
            .O(N__47155),
            .I(N__47149));
    CascadeMux I__9563 (
            .O(N__47154),
            .I(N__47146));
    CascadeMux I__9562 (
            .O(N__47153),
            .I(N__47142));
    CascadeMux I__9561 (
            .O(N__47152),
            .I(N__47139));
    InMux I__9560 (
            .O(N__47149),
            .I(N__47136));
    InMux I__9559 (
            .O(N__47146),
            .I(N__47131));
    InMux I__9558 (
            .O(N__47145),
            .I(N__47131));
    InMux I__9557 (
            .O(N__47142),
            .I(N__47128));
    InMux I__9556 (
            .O(N__47139),
            .I(N__47125));
    LocalMux I__9555 (
            .O(N__47136),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__9554 (
            .O(N__47131),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__9553 (
            .O(N__47128),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__9552 (
            .O(N__47125),
            .I(\c0.data_in_frame_4_5 ));
    InMux I__9551 (
            .O(N__47116),
            .I(N__47113));
    LocalMux I__9550 (
            .O(N__47113),
            .I(\c0.n54 ));
    InMux I__9549 (
            .O(N__47110),
            .I(N__47107));
    LocalMux I__9548 (
            .O(N__47107),
            .I(\c0.n90 ));
    InMux I__9547 (
            .O(N__47104),
            .I(N__47101));
    LocalMux I__9546 (
            .O(N__47101),
            .I(\c0.n98 ));
    InMux I__9545 (
            .O(N__47098),
            .I(N__47095));
    LocalMux I__9544 (
            .O(N__47095),
            .I(N__47092));
    Span4Mux_v I__9543 (
            .O(N__47092),
            .I(N__47089));
    Odrv4 I__9542 (
            .O(N__47089),
            .I(\c0.n12085 ));
    InMux I__9541 (
            .O(N__47086),
            .I(N__47083));
    LocalMux I__9540 (
            .O(N__47083),
            .I(N__47079));
    InMux I__9539 (
            .O(N__47082),
            .I(N__47076));
    Odrv4 I__9538 (
            .O(N__47079),
            .I(\c0.n11865 ));
    LocalMux I__9537 (
            .O(N__47076),
            .I(\c0.n11865 ));
    CascadeMux I__9536 (
            .O(N__47071),
            .I(\c0.n12085_cascade_ ));
    CascadeMux I__9535 (
            .O(N__47068),
            .I(N__47065));
    InMux I__9534 (
            .O(N__47065),
            .I(N__47062));
    LocalMux I__9533 (
            .O(N__47062),
            .I(N__47059));
    Span4Mux_h I__9532 (
            .O(N__47059),
            .I(N__47056));
    Span4Mux_v I__9531 (
            .O(N__47056),
            .I(N__47053));
    Span4Mux_h I__9530 (
            .O(N__47053),
            .I(N__47049));
    InMux I__9529 (
            .O(N__47052),
            .I(N__47046));
    Odrv4 I__9528 (
            .O(N__47049),
            .I(\c0.n6495 ));
    LocalMux I__9527 (
            .O(N__47046),
            .I(\c0.n6495 ));
    InMux I__9526 (
            .O(N__47041),
            .I(N__47038));
    LocalMux I__9525 (
            .O(N__47038),
            .I(N__47035));
    Span4Mux_h I__9524 (
            .O(N__47035),
            .I(N__47029));
    InMux I__9523 (
            .O(N__47034),
            .I(N__47026));
    InMux I__9522 (
            .O(N__47033),
            .I(N__47021));
    InMux I__9521 (
            .O(N__47032),
            .I(N__47021));
    Odrv4 I__9520 (
            .O(N__47029),
            .I(data_in_2_4));
    LocalMux I__9519 (
            .O(N__47026),
            .I(data_in_2_4));
    LocalMux I__9518 (
            .O(N__47021),
            .I(data_in_2_4));
    CascadeMux I__9517 (
            .O(N__47014),
            .I(N__47010));
    CascadeMux I__9516 (
            .O(N__47013),
            .I(N__47007));
    InMux I__9515 (
            .O(N__47010),
            .I(N__47003));
    InMux I__9514 (
            .O(N__47007),
            .I(N__47000));
    InMux I__9513 (
            .O(N__47006),
            .I(N__46997));
    LocalMux I__9512 (
            .O(N__47003),
            .I(N__46994));
    LocalMux I__9511 (
            .O(N__47000),
            .I(N__46987));
    LocalMux I__9510 (
            .O(N__46997),
            .I(N__46987));
    Span4Mux_h I__9509 (
            .O(N__46994),
            .I(N__46984));
    InMux I__9508 (
            .O(N__46993),
            .I(N__46981));
    InMux I__9507 (
            .O(N__46992),
            .I(N__46978));
    Span4Mux_h I__9506 (
            .O(N__46987),
            .I(N__46975));
    Span4Mux_v I__9505 (
            .O(N__46984),
            .I(N__46972));
    LocalMux I__9504 (
            .O(N__46981),
            .I(data_in_1_4));
    LocalMux I__9503 (
            .O(N__46978),
            .I(data_in_1_4));
    Odrv4 I__9502 (
            .O(N__46975),
            .I(data_in_1_4));
    Odrv4 I__9501 (
            .O(N__46972),
            .I(data_in_1_4));
    InMux I__9500 (
            .O(N__46963),
            .I(N__46960));
    LocalMux I__9499 (
            .O(N__46960),
            .I(N__46957));
    Span4Mux_v I__9498 (
            .O(N__46957),
            .I(N__46954));
    Odrv4 I__9497 (
            .O(N__46954),
            .I(\c0.n6_adj_3343 ));
    InMux I__9496 (
            .O(N__46951),
            .I(N__46948));
    LocalMux I__9495 (
            .O(N__46948),
            .I(N__46945));
    Span12Mux_v I__9494 (
            .O(N__46945),
            .I(N__46942));
    Odrv12 I__9493 (
            .O(N__46942),
            .I(\c0.data_out_frame_28_7 ));
    InMux I__9492 (
            .O(N__46939),
            .I(N__46924));
    InMux I__9491 (
            .O(N__46938),
            .I(N__46924));
    SRMux I__9490 (
            .O(N__46937),
            .I(N__46911));
    CEMux I__9489 (
            .O(N__46936),
            .I(N__46908));
    InMux I__9488 (
            .O(N__46935),
            .I(N__46890));
    InMux I__9487 (
            .O(N__46934),
            .I(N__46890));
    InMux I__9486 (
            .O(N__46933),
            .I(N__46890));
    InMux I__9485 (
            .O(N__46932),
            .I(N__46890));
    InMux I__9484 (
            .O(N__46931),
            .I(N__46890));
    InMux I__9483 (
            .O(N__46930),
            .I(N__46881));
    InMux I__9482 (
            .O(N__46929),
            .I(N__46881));
    LocalMux I__9481 (
            .O(N__46924),
            .I(N__46878));
    InMux I__9480 (
            .O(N__46923),
            .I(N__46867));
    InMux I__9479 (
            .O(N__46922),
            .I(N__46867));
    InMux I__9478 (
            .O(N__46921),
            .I(N__46867));
    InMux I__9477 (
            .O(N__46920),
            .I(N__46867));
    InMux I__9476 (
            .O(N__46919),
            .I(N__46867));
    InMux I__9475 (
            .O(N__46918),
            .I(N__46861));
    CascadeMux I__9474 (
            .O(N__46917),
            .I(N__46852));
    CascadeMux I__9473 (
            .O(N__46916),
            .I(N__46849));
    InMux I__9472 (
            .O(N__46915),
            .I(N__46843));
    InMux I__9471 (
            .O(N__46914),
            .I(N__46843));
    LocalMux I__9470 (
            .O(N__46911),
            .I(N__46840));
    LocalMux I__9469 (
            .O(N__46908),
            .I(N__46837));
    InMux I__9468 (
            .O(N__46907),
            .I(N__46830));
    InMux I__9467 (
            .O(N__46906),
            .I(N__46830));
    InMux I__9466 (
            .O(N__46905),
            .I(N__46830));
    CascadeMux I__9465 (
            .O(N__46904),
            .I(N__46827));
    InMux I__9464 (
            .O(N__46903),
            .I(N__46821));
    InMux I__9463 (
            .O(N__46902),
            .I(N__46816));
    InMux I__9462 (
            .O(N__46901),
            .I(N__46816));
    LocalMux I__9461 (
            .O(N__46890),
            .I(N__46813));
    InMux I__9460 (
            .O(N__46889),
            .I(N__46810));
    InMux I__9459 (
            .O(N__46888),
            .I(N__46807));
    InMux I__9458 (
            .O(N__46887),
            .I(N__46804));
    InMux I__9457 (
            .O(N__46886),
            .I(N__46800));
    LocalMux I__9456 (
            .O(N__46881),
            .I(N__46788));
    Span4Mux_v I__9455 (
            .O(N__46878),
            .I(N__46788));
    LocalMux I__9454 (
            .O(N__46867),
            .I(N__46788));
    InMux I__9453 (
            .O(N__46866),
            .I(N__46781));
    InMux I__9452 (
            .O(N__46865),
            .I(N__46781));
    InMux I__9451 (
            .O(N__46864),
            .I(N__46781));
    LocalMux I__9450 (
            .O(N__46861),
            .I(N__46776));
    InMux I__9449 (
            .O(N__46860),
            .I(N__46773));
    InMux I__9448 (
            .O(N__46859),
            .I(N__46770));
    CEMux I__9447 (
            .O(N__46858),
            .I(N__46767));
    CascadeMux I__9446 (
            .O(N__46857),
            .I(N__46761));
    InMux I__9445 (
            .O(N__46856),
            .I(N__46756));
    InMux I__9444 (
            .O(N__46855),
            .I(N__46756));
    InMux I__9443 (
            .O(N__46852),
            .I(N__46749));
    InMux I__9442 (
            .O(N__46849),
            .I(N__46749));
    InMux I__9441 (
            .O(N__46848),
            .I(N__46749));
    LocalMux I__9440 (
            .O(N__46843),
            .I(N__46744));
    Span4Mux_v I__9439 (
            .O(N__46840),
            .I(N__46744));
    Span4Mux_v I__9438 (
            .O(N__46837),
            .I(N__46739));
    LocalMux I__9437 (
            .O(N__46830),
            .I(N__46739));
    InMux I__9436 (
            .O(N__46827),
            .I(N__46714));
    InMux I__9435 (
            .O(N__46826),
            .I(N__46714));
    InMux I__9434 (
            .O(N__46825),
            .I(N__46714));
    InMux I__9433 (
            .O(N__46824),
            .I(N__46714));
    LocalMux I__9432 (
            .O(N__46821),
            .I(N__46709));
    LocalMux I__9431 (
            .O(N__46816),
            .I(N__46709));
    Span4Mux_h I__9430 (
            .O(N__46813),
            .I(N__46704));
    LocalMux I__9429 (
            .O(N__46810),
            .I(N__46704));
    LocalMux I__9428 (
            .O(N__46807),
            .I(N__46699));
    LocalMux I__9427 (
            .O(N__46804),
            .I(N__46699));
    SRMux I__9426 (
            .O(N__46803),
            .I(N__46696));
    LocalMux I__9425 (
            .O(N__46800),
            .I(N__46693));
    InMux I__9424 (
            .O(N__46799),
            .I(N__46688));
    InMux I__9423 (
            .O(N__46798),
            .I(N__46683));
    InMux I__9422 (
            .O(N__46797),
            .I(N__46683));
    InMux I__9421 (
            .O(N__46796),
            .I(N__46678));
    InMux I__9420 (
            .O(N__46795),
            .I(N__46678));
    Span4Mux_h I__9419 (
            .O(N__46788),
            .I(N__46673));
    LocalMux I__9418 (
            .O(N__46781),
            .I(N__46673));
    InMux I__9417 (
            .O(N__46780),
            .I(N__46668));
    InMux I__9416 (
            .O(N__46779),
            .I(N__46668));
    Span4Mux_h I__9415 (
            .O(N__46776),
            .I(N__46665));
    LocalMux I__9414 (
            .O(N__46773),
            .I(N__46658));
    LocalMux I__9413 (
            .O(N__46770),
            .I(N__46658));
    LocalMux I__9412 (
            .O(N__46767),
            .I(N__46658));
    CascadeMux I__9411 (
            .O(N__46766),
            .I(N__46655));
    CascadeMux I__9410 (
            .O(N__46765),
            .I(N__46652));
    InMux I__9409 (
            .O(N__46764),
            .I(N__46639));
    InMux I__9408 (
            .O(N__46761),
            .I(N__46636));
    LocalMux I__9407 (
            .O(N__46756),
            .I(N__46627));
    LocalMux I__9406 (
            .O(N__46749),
            .I(N__46627));
    Span4Mux_h I__9405 (
            .O(N__46744),
            .I(N__46627));
    Span4Mux_h I__9404 (
            .O(N__46739),
            .I(N__46627));
    SRMux I__9403 (
            .O(N__46738),
            .I(N__46624));
    InMux I__9402 (
            .O(N__46737),
            .I(N__46619));
    InMux I__9401 (
            .O(N__46736),
            .I(N__46610));
    InMux I__9400 (
            .O(N__46735),
            .I(N__46610));
    InMux I__9399 (
            .O(N__46734),
            .I(N__46610));
    InMux I__9398 (
            .O(N__46733),
            .I(N__46610));
    InMux I__9397 (
            .O(N__46732),
            .I(N__46603));
    InMux I__9396 (
            .O(N__46731),
            .I(N__46603));
    InMux I__9395 (
            .O(N__46730),
            .I(N__46603));
    SRMux I__9394 (
            .O(N__46729),
            .I(N__46600));
    InMux I__9393 (
            .O(N__46728),
            .I(N__46593));
    InMux I__9392 (
            .O(N__46727),
            .I(N__46593));
    InMux I__9391 (
            .O(N__46726),
            .I(N__46593));
    InMux I__9390 (
            .O(N__46725),
            .I(N__46588));
    InMux I__9389 (
            .O(N__46724),
            .I(N__46588));
    InMux I__9388 (
            .O(N__46723),
            .I(N__46585));
    LocalMux I__9387 (
            .O(N__46714),
            .I(N__46582));
    Span4Mux_v I__9386 (
            .O(N__46709),
            .I(N__46577));
    Span4Mux_v I__9385 (
            .O(N__46704),
            .I(N__46577));
    Span4Mux_v I__9384 (
            .O(N__46699),
            .I(N__46572));
    LocalMux I__9383 (
            .O(N__46696),
            .I(N__46572));
    Span4Mux_v I__9382 (
            .O(N__46693),
            .I(N__46569));
    InMux I__9381 (
            .O(N__46692),
            .I(N__46564));
    InMux I__9380 (
            .O(N__46691),
            .I(N__46564));
    LocalMux I__9379 (
            .O(N__46688),
            .I(N__46549));
    LocalMux I__9378 (
            .O(N__46683),
            .I(N__46549));
    LocalMux I__9377 (
            .O(N__46678),
            .I(N__46549));
    Span4Mux_h I__9376 (
            .O(N__46673),
            .I(N__46549));
    LocalMux I__9375 (
            .O(N__46668),
            .I(N__46549));
    Span4Mux_h I__9374 (
            .O(N__46665),
            .I(N__46549));
    Span4Mux_h I__9373 (
            .O(N__46658),
            .I(N__46549));
    InMux I__9372 (
            .O(N__46655),
            .I(N__46542));
    InMux I__9371 (
            .O(N__46652),
            .I(N__46542));
    InMux I__9370 (
            .O(N__46651),
            .I(N__46542));
    InMux I__9369 (
            .O(N__46650),
            .I(N__46531));
    InMux I__9368 (
            .O(N__46649),
            .I(N__46531));
    InMux I__9367 (
            .O(N__46648),
            .I(N__46531));
    InMux I__9366 (
            .O(N__46647),
            .I(N__46531));
    InMux I__9365 (
            .O(N__46646),
            .I(N__46531));
    InMux I__9364 (
            .O(N__46645),
            .I(N__46526));
    InMux I__9363 (
            .O(N__46644),
            .I(N__46526));
    InMux I__9362 (
            .O(N__46643),
            .I(N__46523));
    InMux I__9361 (
            .O(N__46642),
            .I(N__46520));
    LocalMux I__9360 (
            .O(N__46639),
            .I(N__46513));
    LocalMux I__9359 (
            .O(N__46636),
            .I(N__46513));
    Span4Mux_v I__9358 (
            .O(N__46627),
            .I(N__46513));
    LocalMux I__9357 (
            .O(N__46624),
            .I(N__46510));
    InMux I__9356 (
            .O(N__46623),
            .I(N__46505));
    InMux I__9355 (
            .O(N__46622),
            .I(N__46505));
    LocalMux I__9354 (
            .O(N__46619),
            .I(N__46498));
    LocalMux I__9353 (
            .O(N__46610),
            .I(N__46498));
    LocalMux I__9352 (
            .O(N__46603),
            .I(N__46498));
    LocalMux I__9351 (
            .O(N__46600),
            .I(N__46495));
    LocalMux I__9350 (
            .O(N__46593),
            .I(N__46490));
    LocalMux I__9349 (
            .O(N__46588),
            .I(N__46490));
    LocalMux I__9348 (
            .O(N__46585),
            .I(N__46485));
    Span4Mux_v I__9347 (
            .O(N__46582),
            .I(N__46485));
    Span4Mux_v I__9346 (
            .O(N__46577),
            .I(N__46478));
    Span4Mux_v I__9345 (
            .O(N__46572),
            .I(N__46478));
    Span4Mux_h I__9344 (
            .O(N__46569),
            .I(N__46478));
    LocalMux I__9343 (
            .O(N__46564),
            .I(N__46473));
    Sp12to4 I__9342 (
            .O(N__46549),
            .I(N__46473));
    LocalMux I__9341 (
            .O(N__46542),
            .I(N__46468));
    LocalMux I__9340 (
            .O(N__46531),
            .I(N__46468));
    LocalMux I__9339 (
            .O(N__46526),
            .I(N__46463));
    LocalMux I__9338 (
            .O(N__46523),
            .I(N__46463));
    LocalMux I__9337 (
            .O(N__46520),
            .I(N__46458));
    Span4Mux_v I__9336 (
            .O(N__46513),
            .I(N__46458));
    Span4Mux_v I__9335 (
            .O(N__46510),
            .I(N__46455));
    LocalMux I__9334 (
            .O(N__46505),
            .I(N__46450));
    Span4Mux_v I__9333 (
            .O(N__46498),
            .I(N__46450));
    Span4Mux_h I__9332 (
            .O(N__46495),
            .I(N__46443));
    Span4Mux_v I__9331 (
            .O(N__46490),
            .I(N__46443));
    Span4Mux_h I__9330 (
            .O(N__46485),
            .I(N__46443));
    Sp12to4 I__9329 (
            .O(N__46478),
            .I(N__46438));
    Span12Mux_v I__9328 (
            .O(N__46473),
            .I(N__46438));
    Span4Mux_v I__9327 (
            .O(N__46468),
            .I(N__46431));
    Span4Mux_h I__9326 (
            .O(N__46463),
            .I(N__46431));
    Span4Mux_h I__9325 (
            .O(N__46458),
            .I(N__46431));
    Odrv4 I__9324 (
            .O(N__46455),
            .I(n8112));
    Odrv4 I__9323 (
            .O(N__46450),
            .I(n8112));
    Odrv4 I__9322 (
            .O(N__46443),
            .I(n8112));
    Odrv12 I__9321 (
            .O(N__46438),
            .I(n8112));
    Odrv4 I__9320 (
            .O(N__46431),
            .I(n8112));
    CascadeMux I__9319 (
            .O(N__46420),
            .I(N__46417));
    InMux I__9318 (
            .O(N__46417),
            .I(N__46411));
    InMux I__9317 (
            .O(N__46416),
            .I(N__46408));
    InMux I__9316 (
            .O(N__46415),
            .I(N__46405));
    InMux I__9315 (
            .O(N__46414),
            .I(N__46402));
    LocalMux I__9314 (
            .O(N__46411),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__9313 (
            .O(N__46408),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__9312 (
            .O(N__46405),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__9311 (
            .O(N__46402),
            .I(\c0.data_in_frame_4_3 ));
    InMux I__9310 (
            .O(N__46393),
            .I(N__46387));
    InMux I__9309 (
            .O(N__46392),
            .I(N__46384));
    InMux I__9308 (
            .O(N__46391),
            .I(N__46381));
    InMux I__9307 (
            .O(N__46390),
            .I(N__46378));
    LocalMux I__9306 (
            .O(N__46387),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__9305 (
            .O(N__46384),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__9304 (
            .O(N__46381),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__9303 (
            .O(N__46378),
            .I(\c0.data_in_frame_4_2 ));
    CascadeMux I__9302 (
            .O(N__46369),
            .I(N__46365));
    CascadeMux I__9301 (
            .O(N__46368),
            .I(N__46362));
    InMux I__9300 (
            .O(N__46365),
            .I(N__46359));
    InMux I__9299 (
            .O(N__46362),
            .I(N__46356));
    LocalMux I__9298 (
            .O(N__46359),
            .I(N__46351));
    LocalMux I__9297 (
            .O(N__46356),
            .I(N__46351));
    Odrv12 I__9296 (
            .O(N__46351),
            .I(\c0.data_in_frame_6_4 ));
    CascadeMux I__9295 (
            .O(N__46348),
            .I(\c0.n13_adj_3496_cascade_ ));
    CascadeMux I__9294 (
            .O(N__46345),
            .I(N__46342));
    InMux I__9293 (
            .O(N__46342),
            .I(N__46338));
    InMux I__9292 (
            .O(N__46341),
            .I(N__46335));
    LocalMux I__9291 (
            .O(N__46338),
            .I(N__46330));
    LocalMux I__9290 (
            .O(N__46335),
            .I(N__46327));
    InMux I__9289 (
            .O(N__46334),
            .I(N__46324));
    InMux I__9288 (
            .O(N__46333),
            .I(N__46321));
    Span4Mux_h I__9287 (
            .O(N__46330),
            .I(N__46318));
    Span4Mux_h I__9286 (
            .O(N__46327),
            .I(N__46315));
    LocalMux I__9285 (
            .O(N__46324),
            .I(N__46312));
    LocalMux I__9284 (
            .O(N__46321),
            .I(\c0.data_in_frame_2_2 ));
    Odrv4 I__9283 (
            .O(N__46318),
            .I(\c0.data_in_frame_2_2 ));
    Odrv4 I__9282 (
            .O(N__46315),
            .I(\c0.data_in_frame_2_2 ));
    Odrv12 I__9281 (
            .O(N__46312),
            .I(\c0.data_in_frame_2_2 ));
    InMux I__9280 (
            .O(N__46303),
            .I(N__46297));
    InMux I__9279 (
            .O(N__46302),
            .I(N__46294));
    InMux I__9278 (
            .O(N__46301),
            .I(N__46289));
    CascadeMux I__9277 (
            .O(N__46300),
            .I(N__46284));
    LocalMux I__9276 (
            .O(N__46297),
            .I(N__46280));
    LocalMux I__9275 (
            .O(N__46294),
            .I(N__46277));
    CascadeMux I__9274 (
            .O(N__46293),
            .I(N__46274));
    CascadeMux I__9273 (
            .O(N__46292),
            .I(N__46270));
    LocalMux I__9272 (
            .O(N__46289),
            .I(N__46266));
    CascadeMux I__9271 (
            .O(N__46288),
            .I(N__46262));
    InMux I__9270 (
            .O(N__46287),
            .I(N__46257));
    InMux I__9269 (
            .O(N__46284),
            .I(N__46257));
    InMux I__9268 (
            .O(N__46283),
            .I(N__46254));
    Span4Mux_v I__9267 (
            .O(N__46280),
            .I(N__46251));
    Span4Mux_h I__9266 (
            .O(N__46277),
            .I(N__46248));
    InMux I__9265 (
            .O(N__46274),
            .I(N__46241));
    InMux I__9264 (
            .O(N__46273),
            .I(N__46241));
    InMux I__9263 (
            .O(N__46270),
            .I(N__46241));
    InMux I__9262 (
            .O(N__46269),
            .I(N__46238));
    Span4Mux_h I__9261 (
            .O(N__46266),
            .I(N__46235));
    InMux I__9260 (
            .O(N__46265),
            .I(N__46230));
    InMux I__9259 (
            .O(N__46262),
            .I(N__46230));
    LocalMux I__9258 (
            .O(N__46257),
            .I(data_in_frame_0_0));
    LocalMux I__9257 (
            .O(N__46254),
            .I(data_in_frame_0_0));
    Odrv4 I__9256 (
            .O(N__46251),
            .I(data_in_frame_0_0));
    Odrv4 I__9255 (
            .O(N__46248),
            .I(data_in_frame_0_0));
    LocalMux I__9254 (
            .O(N__46241),
            .I(data_in_frame_0_0));
    LocalMux I__9253 (
            .O(N__46238),
            .I(data_in_frame_0_0));
    Odrv4 I__9252 (
            .O(N__46235),
            .I(data_in_frame_0_0));
    LocalMux I__9251 (
            .O(N__46230),
            .I(data_in_frame_0_0));
    InMux I__9250 (
            .O(N__46213),
            .I(N__46210));
    LocalMux I__9249 (
            .O(N__46210),
            .I(\c0.n19277 ));
    InMux I__9248 (
            .O(N__46207),
            .I(N__46203));
    CascadeMux I__9247 (
            .O(N__46206),
            .I(N__46200));
    LocalMux I__9246 (
            .O(N__46203),
            .I(N__46197));
    InMux I__9245 (
            .O(N__46200),
            .I(N__46194));
    Odrv4 I__9244 (
            .O(N__46197),
            .I(\c0.n7_adj_3078 ));
    LocalMux I__9243 (
            .O(N__46194),
            .I(\c0.n7_adj_3078 ));
    InMux I__9242 (
            .O(N__46189),
            .I(N__46186));
    LocalMux I__9241 (
            .O(N__46186),
            .I(N__46183));
    Span4Mux_v I__9240 (
            .O(N__46183),
            .I(N__46180));
    Odrv4 I__9239 (
            .O(N__46180),
            .I(\c0.n17880 ));
    InMux I__9238 (
            .O(N__46177),
            .I(N__46174));
    LocalMux I__9237 (
            .O(N__46174),
            .I(N__46171));
    Odrv4 I__9236 (
            .O(N__46171),
            .I(\c0.n26_adj_3523 ));
    CascadeMux I__9235 (
            .O(N__46168),
            .I(N__46164));
    InMux I__9234 (
            .O(N__46167),
            .I(N__46161));
    InMux I__9233 (
            .O(N__46164),
            .I(N__46158));
    LocalMux I__9232 (
            .O(N__46161),
            .I(data_in_0_4));
    LocalMux I__9231 (
            .O(N__46158),
            .I(data_in_0_4));
    InMux I__9230 (
            .O(N__46153),
            .I(N__46149));
    InMux I__9229 (
            .O(N__46152),
            .I(N__46146));
    LocalMux I__9228 (
            .O(N__46149),
            .I(N__46143));
    LocalMux I__9227 (
            .O(N__46146),
            .I(N__46140));
    Span4Mux_h I__9226 (
            .O(N__46143),
            .I(N__46131));
    Span4Mux_v I__9225 (
            .O(N__46140),
            .I(N__46128));
    InMux I__9224 (
            .O(N__46139),
            .I(N__46125));
    InMux I__9223 (
            .O(N__46138),
            .I(N__46116));
    InMux I__9222 (
            .O(N__46137),
            .I(N__46116));
    InMux I__9221 (
            .O(N__46136),
            .I(N__46116));
    InMux I__9220 (
            .O(N__46135),
            .I(N__46116));
    InMux I__9219 (
            .O(N__46134),
            .I(N__46113));
    Odrv4 I__9218 (
            .O(N__46131),
            .I(n20896));
    Odrv4 I__9217 (
            .O(N__46128),
            .I(n20896));
    LocalMux I__9216 (
            .O(N__46125),
            .I(n20896));
    LocalMux I__9215 (
            .O(N__46116),
            .I(n20896));
    LocalMux I__9214 (
            .O(N__46113),
            .I(n20896));
    InMux I__9213 (
            .O(N__46102),
            .I(N__46099));
    LocalMux I__9212 (
            .O(N__46099),
            .I(\c0.n18457 ));
    InMux I__9211 (
            .O(N__46096),
            .I(N__46090));
    InMux I__9210 (
            .O(N__46095),
            .I(N__46087));
    InMux I__9209 (
            .O(N__46094),
            .I(N__46084));
    InMux I__9208 (
            .O(N__46093),
            .I(N__46081));
    LocalMux I__9207 (
            .O(N__46090),
            .I(N__46078));
    LocalMux I__9206 (
            .O(N__46087),
            .I(N__46075));
    LocalMux I__9205 (
            .O(N__46084),
            .I(\c0.n21076 ));
    LocalMux I__9204 (
            .O(N__46081),
            .I(\c0.n21076 ));
    Odrv4 I__9203 (
            .O(N__46078),
            .I(\c0.n21076 ));
    Odrv4 I__9202 (
            .O(N__46075),
            .I(\c0.n21076 ));
    InMux I__9201 (
            .O(N__46066),
            .I(N__46063));
    LocalMux I__9200 (
            .O(N__46063),
            .I(N__46060));
    Odrv12 I__9199 (
            .O(N__46060),
            .I(\c0.n33_adj_3308 ));
    CascadeMux I__9198 (
            .O(N__46057),
            .I(N__46054));
    InMux I__9197 (
            .O(N__46054),
            .I(N__46048));
    InMux I__9196 (
            .O(N__46053),
            .I(N__46048));
    LocalMux I__9195 (
            .O(N__46048),
            .I(\c0.n18417 ));
    CascadeMux I__9194 (
            .O(N__46045),
            .I(\c0.n18417_cascade_ ));
    InMux I__9193 (
            .O(N__46042),
            .I(N__46039));
    LocalMux I__9192 (
            .O(N__46039),
            .I(\c0.n19_adj_3292 ));
    InMux I__9191 (
            .O(N__46036),
            .I(N__46030));
    InMux I__9190 (
            .O(N__46035),
            .I(N__46030));
    LocalMux I__9189 (
            .O(N__46030),
            .I(\c0.data_in_frame_29_4 ));
    InMux I__9188 (
            .O(N__46027),
            .I(N__46024));
    LocalMux I__9187 (
            .O(N__46024),
            .I(N__46020));
    CascadeMux I__9186 (
            .O(N__46023),
            .I(N__46017));
    Span4Mux_h I__9185 (
            .O(N__46020),
            .I(N__46014));
    InMux I__9184 (
            .O(N__46017),
            .I(N__46011));
    Span4Mux_v I__9183 (
            .O(N__46014),
            .I(N__46008));
    LocalMux I__9182 (
            .O(N__46011),
            .I(\c0.data_in_frame_29_2 ));
    Odrv4 I__9181 (
            .O(N__46008),
            .I(\c0.data_in_frame_29_2 ));
    InMux I__9180 (
            .O(N__46003),
            .I(N__46000));
    LocalMux I__9179 (
            .O(N__46000),
            .I(N__45996));
    InMux I__9178 (
            .O(N__45999),
            .I(N__45993));
    Span4Mux_h I__9177 (
            .O(N__45996),
            .I(N__45990));
    LocalMux I__9176 (
            .O(N__45993),
            .I(\c0.data_in_frame_29_1 ));
    Odrv4 I__9175 (
            .O(N__45990),
            .I(\c0.data_in_frame_29_1 ));
    CascadeMux I__9174 (
            .O(N__45985),
            .I(N__45982));
    InMux I__9173 (
            .O(N__45982),
            .I(N__45979));
    LocalMux I__9172 (
            .O(N__45979),
            .I(N__45976));
    Span4Mux_v I__9171 (
            .O(N__45976),
            .I(N__45972));
    InMux I__9170 (
            .O(N__45975),
            .I(N__45969));
    Span4Mux_v I__9169 (
            .O(N__45972),
            .I(N__45966));
    LocalMux I__9168 (
            .O(N__45969),
            .I(N__45963));
    Span4Mux_h I__9167 (
            .O(N__45966),
            .I(N__45960));
    Odrv4 I__9166 (
            .O(N__45963),
            .I(\c0.data_in_frame_28_1 ));
    Odrv4 I__9165 (
            .O(N__45960),
            .I(\c0.data_in_frame_28_1 ));
    CascadeMux I__9164 (
            .O(N__45955),
            .I(N__45951));
    CascadeMux I__9163 (
            .O(N__45954),
            .I(N__45948));
    InMux I__9162 (
            .O(N__45951),
            .I(N__45945));
    InMux I__9161 (
            .O(N__45948),
            .I(N__45942));
    LocalMux I__9160 (
            .O(N__45945),
            .I(\c0.data_in_frame_28_0 ));
    LocalMux I__9159 (
            .O(N__45942),
            .I(\c0.data_in_frame_28_0 ));
    InMux I__9158 (
            .O(N__45937),
            .I(N__45932));
    InMux I__9157 (
            .O(N__45936),
            .I(N__45926));
    InMux I__9156 (
            .O(N__45935),
            .I(N__45923));
    LocalMux I__9155 (
            .O(N__45932),
            .I(N__45920));
    CascadeMux I__9154 (
            .O(N__45931),
            .I(N__45917));
    InMux I__9153 (
            .O(N__45930),
            .I(N__45912));
    InMux I__9152 (
            .O(N__45929),
            .I(N__45912));
    LocalMux I__9151 (
            .O(N__45926),
            .I(N__45909));
    LocalMux I__9150 (
            .O(N__45923),
            .I(N__45906));
    Span4Mux_h I__9149 (
            .O(N__45920),
            .I(N__45903));
    InMux I__9148 (
            .O(N__45917),
            .I(N__45900));
    LocalMux I__9147 (
            .O(N__45912),
            .I(\c0.n20324 ));
    Odrv4 I__9146 (
            .O(N__45909),
            .I(\c0.n20324 ));
    Odrv12 I__9145 (
            .O(N__45906),
            .I(\c0.n20324 ));
    Odrv4 I__9144 (
            .O(N__45903),
            .I(\c0.n20324 ));
    LocalMux I__9143 (
            .O(N__45900),
            .I(\c0.n20324 ));
    InMux I__9142 (
            .O(N__45889),
            .I(N__45886));
    LocalMux I__9141 (
            .O(N__45886),
            .I(N__45883));
    Odrv4 I__9140 (
            .O(N__45883),
            .I(\c0.n14_adj_3349 ));
    CascadeMux I__9139 (
            .O(N__45880),
            .I(\c0.n21044_cascade_ ));
    InMux I__9138 (
            .O(N__45877),
            .I(N__45871));
    InMux I__9137 (
            .O(N__45876),
            .I(N__45871));
    LocalMux I__9136 (
            .O(N__45871),
            .I(N__45865));
    CascadeMux I__9135 (
            .O(N__45870),
            .I(N__45862));
    InMux I__9134 (
            .O(N__45869),
            .I(N__45859));
    CascadeMux I__9133 (
            .O(N__45868),
            .I(N__45856));
    Span4Mux_v I__9132 (
            .O(N__45865),
            .I(N__45853));
    InMux I__9131 (
            .O(N__45862),
            .I(N__45850));
    LocalMux I__9130 (
            .O(N__45859),
            .I(N__45847));
    InMux I__9129 (
            .O(N__45856),
            .I(N__45844));
    Span4Mux_h I__9128 (
            .O(N__45853),
            .I(N__45841));
    LocalMux I__9127 (
            .O(N__45850),
            .I(N__45836));
    Span4Mux_h I__9126 (
            .O(N__45847),
            .I(N__45836));
    LocalMux I__9125 (
            .O(N__45844),
            .I(\c0.data_in_frame_26_7 ));
    Odrv4 I__9124 (
            .O(N__45841),
            .I(\c0.data_in_frame_26_7 ));
    Odrv4 I__9123 (
            .O(N__45836),
            .I(\c0.data_in_frame_26_7 ));
    CascadeMux I__9122 (
            .O(N__45829),
            .I(\c0.n16_adj_3109_cascade_ ));
    InMux I__9121 (
            .O(N__45826),
            .I(N__45822));
    InMux I__9120 (
            .O(N__45825),
            .I(N__45819));
    LocalMux I__9119 (
            .O(N__45822),
            .I(\c0.n21071 ));
    LocalMux I__9118 (
            .O(N__45819),
            .I(\c0.n21071 ));
    CascadeMux I__9117 (
            .O(N__45814),
            .I(N__45811));
    InMux I__9116 (
            .O(N__45811),
            .I(N__45805));
    InMux I__9115 (
            .O(N__45810),
            .I(N__45805));
    LocalMux I__9114 (
            .O(N__45805),
            .I(N__45801));
    InMux I__9113 (
            .O(N__45804),
            .I(N__45798));
    Span4Mux_v I__9112 (
            .O(N__45801),
            .I(N__45793));
    LocalMux I__9111 (
            .O(N__45798),
            .I(N__45793));
    Odrv4 I__9110 (
            .O(N__45793),
            .I(\c0.n20479 ));
    InMux I__9109 (
            .O(N__45790),
            .I(N__45787));
    LocalMux I__9108 (
            .O(N__45787),
            .I(\c0.n77 ));
    InMux I__9107 (
            .O(N__45784),
            .I(N__45781));
    LocalMux I__9106 (
            .O(N__45781),
            .I(N__45777));
    InMux I__9105 (
            .O(N__45780),
            .I(N__45774));
    Span4Mux_h I__9104 (
            .O(N__45777),
            .I(N__45771));
    LocalMux I__9103 (
            .O(N__45774),
            .I(\c0.n34_adj_3096 ));
    Odrv4 I__9102 (
            .O(N__45771),
            .I(\c0.n34_adj_3096 ));
    InMux I__9101 (
            .O(N__45766),
            .I(N__45762));
    InMux I__9100 (
            .O(N__45765),
            .I(N__45759));
    LocalMux I__9099 (
            .O(N__45762),
            .I(N__45756));
    LocalMux I__9098 (
            .O(N__45759),
            .I(N__45753));
    Odrv12 I__9097 (
            .O(N__45756),
            .I(\c0.n32_adj_3095 ));
    Odrv4 I__9096 (
            .O(N__45753),
            .I(\c0.n32_adj_3095 ));
    CascadeMux I__9095 (
            .O(N__45748),
            .I(\c0.n18457_cascade_ ));
    InMux I__9094 (
            .O(N__45745),
            .I(N__45741));
    InMux I__9093 (
            .O(N__45744),
            .I(N__45738));
    LocalMux I__9092 (
            .O(N__45741),
            .I(\c0.n23_adj_3222 ));
    LocalMux I__9091 (
            .O(N__45738),
            .I(\c0.n23_adj_3222 ));
    CascadeMux I__9090 (
            .O(N__45733),
            .I(\c0.n43_adj_3280_cascade_ ));
    InMux I__9089 (
            .O(N__45730),
            .I(N__45727));
    LocalMux I__9088 (
            .O(N__45727),
            .I(\c0.n41_adj_3281 ));
    InMux I__9087 (
            .O(N__45724),
            .I(N__45721));
    LocalMux I__9086 (
            .O(N__45721),
            .I(\c0.n50_adj_3283 ));
    CascadeMux I__9085 (
            .O(N__45718),
            .I(\c0.n19511_cascade_ ));
    InMux I__9084 (
            .O(N__45715),
            .I(N__45710));
    InMux I__9083 (
            .O(N__45714),
            .I(N__45705));
    InMux I__9082 (
            .O(N__45713),
            .I(N__45705));
    LocalMux I__9081 (
            .O(N__45710),
            .I(N__45699));
    LocalMux I__9080 (
            .O(N__45705),
            .I(N__45696));
    InMux I__9079 (
            .O(N__45704),
            .I(N__45691));
    InMux I__9078 (
            .O(N__45703),
            .I(N__45691));
    InMux I__9077 (
            .O(N__45702),
            .I(N__45688));
    Span4Mux_v I__9076 (
            .O(N__45699),
            .I(N__45685));
    Sp12to4 I__9075 (
            .O(N__45696),
            .I(N__45680));
    LocalMux I__9074 (
            .O(N__45691),
            .I(N__45680));
    LocalMux I__9073 (
            .O(N__45688),
            .I(\c0.n21110 ));
    Odrv4 I__9072 (
            .O(N__45685),
            .I(\c0.n21110 ));
    Odrv12 I__9071 (
            .O(N__45680),
            .I(\c0.n21110 ));
    InMux I__9070 (
            .O(N__45673),
            .I(N__45670));
    LocalMux I__9069 (
            .O(N__45670),
            .I(N__45667));
    Span12Mux_v I__9068 (
            .O(N__45667),
            .I(N__45664));
    Odrv12 I__9067 (
            .O(N__45664),
            .I(\c0.n20_adj_3448 ));
    InMux I__9066 (
            .O(N__45661),
            .I(N__45657));
    InMux I__9065 (
            .O(N__45660),
            .I(N__45654));
    LocalMux I__9064 (
            .O(N__45657),
            .I(\c0.n20431 ));
    LocalMux I__9063 (
            .O(N__45654),
            .I(\c0.n20431 ));
    InMux I__9062 (
            .O(N__45649),
            .I(N__45646));
    LocalMux I__9061 (
            .O(N__45646),
            .I(N__45643));
    Odrv12 I__9060 (
            .O(N__45643),
            .I(\c0.n64_adj_3512 ));
    InMux I__9059 (
            .O(N__45640),
            .I(N__45634));
    CascadeMux I__9058 (
            .O(N__45639),
            .I(N__45630));
    InMux I__9057 (
            .O(N__45638),
            .I(N__45626));
    InMux I__9056 (
            .O(N__45637),
            .I(N__45623));
    LocalMux I__9055 (
            .O(N__45634),
            .I(N__45620));
    InMux I__9054 (
            .O(N__45633),
            .I(N__45613));
    InMux I__9053 (
            .O(N__45630),
            .I(N__45613));
    InMux I__9052 (
            .O(N__45629),
            .I(N__45613));
    LocalMux I__9051 (
            .O(N__45626),
            .I(N__45609));
    LocalMux I__9050 (
            .O(N__45623),
            .I(N__45606));
    Span4Mux_v I__9049 (
            .O(N__45620),
            .I(N__45603));
    LocalMux I__9048 (
            .O(N__45613),
            .I(N__45600));
    InMux I__9047 (
            .O(N__45612),
            .I(N__45597));
    Span4Mux_h I__9046 (
            .O(N__45609),
            .I(N__45594));
    Span12Mux_h I__9045 (
            .O(N__45606),
            .I(N__45591));
    Span4Mux_v I__9044 (
            .O(N__45603),
            .I(N__45586));
    Span4Mux_h I__9043 (
            .O(N__45600),
            .I(N__45586));
    LocalMux I__9042 (
            .O(N__45597),
            .I(data_in_frame_16_4));
    Odrv4 I__9041 (
            .O(N__45594),
            .I(data_in_frame_16_4));
    Odrv12 I__9040 (
            .O(N__45591),
            .I(data_in_frame_16_4));
    Odrv4 I__9039 (
            .O(N__45586),
            .I(data_in_frame_16_4));
    InMux I__9038 (
            .O(N__45577),
            .I(N__45574));
    LocalMux I__9037 (
            .O(N__45574),
            .I(N__45571));
    Span4Mux_v I__9036 (
            .O(N__45571),
            .I(N__45568));
    Odrv4 I__9035 (
            .O(N__45568),
            .I(\c0.n7_adj_3440 ));
    InMux I__9034 (
            .O(N__45565),
            .I(N__45561));
    InMux I__9033 (
            .O(N__45564),
            .I(N__45557));
    LocalMux I__9032 (
            .O(N__45561),
            .I(N__45554));
    InMux I__9031 (
            .O(N__45560),
            .I(N__45551));
    LocalMux I__9030 (
            .O(N__45557),
            .I(N__45546));
    Span4Mux_v I__9029 (
            .O(N__45554),
            .I(N__45546));
    LocalMux I__9028 (
            .O(N__45551),
            .I(\c0.data_in_frame_13_0 ));
    Odrv4 I__9027 (
            .O(N__45546),
            .I(\c0.data_in_frame_13_0 ));
    CascadeMux I__9026 (
            .O(N__45541),
            .I(N__45538));
    InMux I__9025 (
            .O(N__45538),
            .I(N__45535));
    LocalMux I__9024 (
            .O(N__45535),
            .I(N__45532));
    Span4Mux_h I__9023 (
            .O(N__45532),
            .I(N__45529));
    Span4Mux_v I__9022 (
            .O(N__45529),
            .I(N__45526));
    Odrv4 I__9021 (
            .O(N__45526),
            .I(\c0.n11_adj_3219 ));
    InMux I__9020 (
            .O(N__45523),
            .I(N__45520));
    LocalMux I__9019 (
            .O(N__45520),
            .I(N__45517));
    Odrv12 I__9018 (
            .O(N__45517),
            .I(\c0.n13_adj_3221 ));
    InMux I__9017 (
            .O(N__45514),
            .I(N__45511));
    LocalMux I__9016 (
            .O(N__45511),
            .I(N__45506));
    InMux I__9015 (
            .O(N__45510),
            .I(N__45501));
    InMux I__9014 (
            .O(N__45509),
            .I(N__45501));
    Odrv4 I__9013 (
            .O(N__45506),
            .I(data_in_frame_23_3));
    LocalMux I__9012 (
            .O(N__45501),
            .I(data_in_frame_23_3));
    InMux I__9011 (
            .O(N__45496),
            .I(N__45493));
    LocalMux I__9010 (
            .O(N__45493),
            .I(\c0.n25_adj_3524 ));
    InMux I__9009 (
            .O(N__45490),
            .I(N__45487));
    LocalMux I__9008 (
            .O(N__45487),
            .I(\c0.n19384 ));
    InMux I__9007 (
            .O(N__45484),
            .I(N__45481));
    LocalMux I__9006 (
            .O(N__45481),
            .I(N__45478));
    Odrv4 I__9005 (
            .O(N__45478),
            .I(\c0.n13_adj_3463 ));
    InMux I__9004 (
            .O(N__45475),
            .I(N__45472));
    LocalMux I__9003 (
            .O(N__45472),
            .I(N__45469));
    Span4Mux_v I__9002 (
            .O(N__45469),
            .I(N__45466));
    Odrv4 I__9001 (
            .O(N__45466),
            .I(\c0.n10 ));
    CascadeMux I__9000 (
            .O(N__45463),
            .I(\c0.n19384_cascade_ ));
    InMux I__8999 (
            .O(N__45460),
            .I(N__45453));
    InMux I__8998 (
            .O(N__45459),
            .I(N__45453));
    CascadeMux I__8997 (
            .O(N__45458),
            .I(N__45449));
    LocalMux I__8996 (
            .O(N__45453),
            .I(N__45446));
    CascadeMux I__8995 (
            .O(N__45452),
            .I(N__45443));
    InMux I__8994 (
            .O(N__45449),
            .I(N__45440));
    Span4Mux_v I__8993 (
            .O(N__45446),
            .I(N__45437));
    InMux I__8992 (
            .O(N__45443),
            .I(N__45434));
    LocalMux I__8991 (
            .O(N__45440),
            .I(N__45430));
    Span4Mux_v I__8990 (
            .O(N__45437),
            .I(N__45425));
    LocalMux I__8989 (
            .O(N__45434),
            .I(N__45425));
    InMux I__8988 (
            .O(N__45433),
            .I(N__45422));
    Span4Mux_h I__8987 (
            .O(N__45430),
            .I(N__45417));
    Span4Mux_h I__8986 (
            .O(N__45425),
            .I(N__45417));
    LocalMux I__8985 (
            .O(N__45422),
            .I(data_in_frame_16_5));
    Odrv4 I__8984 (
            .O(N__45417),
            .I(data_in_frame_16_5));
    InMux I__8983 (
            .O(N__45412),
            .I(N__45409));
    LocalMux I__8982 (
            .O(N__45409),
            .I(N__45405));
    InMux I__8981 (
            .O(N__45408),
            .I(N__45402));
    Span4Mux_v I__8980 (
            .O(N__45405),
            .I(N__45399));
    LocalMux I__8979 (
            .O(N__45402),
            .I(data_in_frame_19_0));
    Odrv4 I__8978 (
            .O(N__45399),
            .I(data_in_frame_19_0));
    CascadeMux I__8977 (
            .O(N__45394),
            .I(\c0.n9_adj_3430_cascade_ ));
    InMux I__8976 (
            .O(N__45391),
            .I(N__45385));
    InMux I__8975 (
            .O(N__45390),
            .I(N__45385));
    LocalMux I__8974 (
            .O(N__45385),
            .I(N__45382));
    Span4Mux_v I__8973 (
            .O(N__45382),
            .I(N__45379));
    Odrv4 I__8972 (
            .O(N__45379),
            .I(\c0.n10_adj_3445 ));
    InMux I__8971 (
            .O(N__45376),
            .I(N__45373));
    LocalMux I__8970 (
            .O(N__45373),
            .I(\c0.n9_adj_3430 ));
    CascadeMux I__8969 (
            .O(N__45370),
            .I(N__45367));
    InMux I__8968 (
            .O(N__45367),
            .I(N__45361));
    InMux I__8967 (
            .O(N__45366),
            .I(N__45361));
    LocalMux I__8966 (
            .O(N__45361),
            .I(\c0.n14_adj_3421 ));
    CascadeMux I__8965 (
            .O(N__45358),
            .I(\c0.n18433_cascade_ ));
    InMux I__8964 (
            .O(N__45355),
            .I(N__45352));
    LocalMux I__8963 (
            .O(N__45352),
            .I(N__45349));
    Odrv4 I__8962 (
            .O(N__45349),
            .I(\c0.n19511 ));
    InMux I__8961 (
            .O(N__45346),
            .I(N__45340));
    InMux I__8960 (
            .O(N__45345),
            .I(N__45340));
    LocalMux I__8959 (
            .O(N__45340),
            .I(N__45335));
    InMux I__8958 (
            .O(N__45339),
            .I(N__45329));
    InMux I__8957 (
            .O(N__45338),
            .I(N__45329));
    Span4Mux_h I__8956 (
            .O(N__45335),
            .I(N__45326));
    InMux I__8955 (
            .O(N__45334),
            .I(N__45323));
    LocalMux I__8954 (
            .O(N__45329),
            .I(\c0.n49 ));
    Odrv4 I__8953 (
            .O(N__45326),
            .I(\c0.n49 ));
    LocalMux I__8952 (
            .O(N__45323),
            .I(\c0.n49 ));
    InMux I__8951 (
            .O(N__45316),
            .I(N__45310));
    InMux I__8950 (
            .O(N__45315),
            .I(N__45310));
    LocalMux I__8949 (
            .O(N__45310),
            .I(N__45307));
    Span4Mux_h I__8948 (
            .O(N__45307),
            .I(N__45303));
    InMux I__8947 (
            .O(N__45306),
            .I(N__45300));
    Span4Mux_h I__8946 (
            .O(N__45303),
            .I(N__45297));
    LocalMux I__8945 (
            .O(N__45300),
            .I(N__45294));
    Span4Mux_h I__8944 (
            .O(N__45297),
            .I(N__45291));
    Span4Mux_h I__8943 (
            .O(N__45294),
            .I(N__45287));
    Sp12to4 I__8942 (
            .O(N__45291),
            .I(N__45284));
    InMux I__8941 (
            .O(N__45290),
            .I(N__45281));
    Odrv4 I__8940 (
            .O(N__45287),
            .I(\c0.n48_adj_3409 ));
    Odrv12 I__8939 (
            .O(N__45284),
            .I(\c0.n48_adj_3409 ));
    LocalMux I__8938 (
            .O(N__45281),
            .I(\c0.n48_adj_3409 ));
    CascadeMux I__8937 (
            .O(N__45274),
            .I(\c0.n22_adj_3287_cascade_ ));
    InMux I__8936 (
            .O(N__45271),
            .I(N__45267));
    InMux I__8935 (
            .O(N__45270),
            .I(N__45264));
    LocalMux I__8934 (
            .O(N__45267),
            .I(N__45259));
    LocalMux I__8933 (
            .O(N__45264),
            .I(N__45259));
    Span4Mux_v I__8932 (
            .O(N__45259),
            .I(N__45256));
    Odrv4 I__8931 (
            .O(N__45256),
            .I(\c0.n39_adj_3050 ));
    CascadeMux I__8930 (
            .O(N__45253),
            .I(\c0.n20451_cascade_ ));
    InMux I__8929 (
            .O(N__45250),
            .I(N__45247));
    LocalMux I__8928 (
            .O(N__45247),
            .I(N__45244));
    Span4Mux_h I__8927 (
            .O(N__45244),
            .I(N__45241));
    Odrv4 I__8926 (
            .O(N__45241),
            .I(\c0.n5_adj_3220 ));
    InMux I__8925 (
            .O(N__45238),
            .I(N__45235));
    LocalMux I__8924 (
            .O(N__45235),
            .I(N__45231));
    InMux I__8923 (
            .O(N__45234),
            .I(N__45228));
    Span4Mux_v I__8922 (
            .O(N__45231),
            .I(N__45225));
    LocalMux I__8921 (
            .O(N__45228),
            .I(data_in_frame_18_1));
    Odrv4 I__8920 (
            .O(N__45225),
            .I(data_in_frame_18_1));
    CascadeMux I__8919 (
            .O(N__45220),
            .I(\c0.n27_adj_3529_cascade_ ));
    CascadeMux I__8918 (
            .O(N__45217),
            .I(\c0.n32_adj_3530_cascade_ ));
    CascadeMux I__8917 (
            .O(N__45214),
            .I(\c0.n19244_cascade_ ));
    InMux I__8916 (
            .O(N__45211),
            .I(N__45208));
    LocalMux I__8915 (
            .O(N__45208),
            .I(N__45205));
    Span4Mux_h I__8914 (
            .O(N__45205),
            .I(N__45202));
    Odrv4 I__8913 (
            .O(N__45202),
            .I(\c0.n85_adj_3074 ));
    CascadeMux I__8912 (
            .O(N__45199),
            .I(\c0.n85_adj_3074_cascade_ ));
    InMux I__8911 (
            .O(N__45196),
            .I(N__45193));
    LocalMux I__8910 (
            .O(N__45193),
            .I(\c0.n10_adj_3474 ));
    InMux I__8909 (
            .O(N__45190),
            .I(N__45183));
    InMux I__8908 (
            .O(N__45189),
            .I(N__45183));
    InMux I__8907 (
            .O(N__45188),
            .I(N__45176));
    LocalMux I__8906 (
            .O(N__45183),
            .I(N__45173));
    InMux I__8905 (
            .O(N__45182),
            .I(N__45170));
    InMux I__8904 (
            .O(N__45181),
            .I(N__45163));
    InMux I__8903 (
            .O(N__45180),
            .I(N__45163));
    InMux I__8902 (
            .O(N__45179),
            .I(N__45163));
    LocalMux I__8901 (
            .O(N__45176),
            .I(\c0.n20801 ));
    Odrv4 I__8900 (
            .O(N__45173),
            .I(\c0.n20801 ));
    LocalMux I__8899 (
            .O(N__45170),
            .I(\c0.n20801 ));
    LocalMux I__8898 (
            .O(N__45163),
            .I(\c0.n20801 ));
    InMux I__8897 (
            .O(N__45154),
            .I(N__45151));
    LocalMux I__8896 (
            .O(N__45151),
            .I(N__45148));
    Span4Mux_v I__8895 (
            .O(N__45148),
            .I(N__45145));
    Odrv4 I__8894 (
            .O(N__45145),
            .I(\c0.n12_adj_3477 ));
    InMux I__8893 (
            .O(N__45142),
            .I(N__45138));
    InMux I__8892 (
            .O(N__45141),
            .I(N__45134));
    LocalMux I__8891 (
            .O(N__45138),
            .I(N__45131));
    InMux I__8890 (
            .O(N__45137),
            .I(N__45128));
    LocalMux I__8889 (
            .O(N__45134),
            .I(N__45124));
    Span4Mux_v I__8888 (
            .O(N__45131),
            .I(N__45121));
    LocalMux I__8887 (
            .O(N__45128),
            .I(N__45118));
    InMux I__8886 (
            .O(N__45127),
            .I(N__45115));
    Span12Mux_v I__8885 (
            .O(N__45124),
            .I(N__45112));
    Span4Mux_h I__8884 (
            .O(N__45121),
            .I(N__45107));
    Span4Mux_v I__8883 (
            .O(N__45118),
            .I(N__45107));
    LocalMux I__8882 (
            .O(N__45115),
            .I(\c0.data_in_frame_14_4 ));
    Odrv12 I__8881 (
            .O(N__45112),
            .I(\c0.data_in_frame_14_4 ));
    Odrv4 I__8880 (
            .O(N__45107),
            .I(\c0.data_in_frame_14_4 ));
    CascadeMux I__8879 (
            .O(N__45100),
            .I(\c0.n21110_cascade_ ));
    InMux I__8878 (
            .O(N__45097),
            .I(N__45094));
    LocalMux I__8877 (
            .O(N__45094),
            .I(N__45090));
    InMux I__8876 (
            .O(N__45093),
            .I(N__45087));
    Span4Mux_v I__8875 (
            .O(N__45090),
            .I(N__45084));
    LocalMux I__8874 (
            .O(N__45087),
            .I(N__45081));
    Span4Mux_v I__8873 (
            .O(N__45084),
            .I(N__45078));
    Span4Mux_v I__8872 (
            .O(N__45081),
            .I(N__45075));
    Odrv4 I__8871 (
            .O(N__45078),
            .I(\c0.n20246 ));
    Odrv4 I__8870 (
            .O(N__45075),
            .I(\c0.n20246 ));
    CascadeMux I__8869 (
            .O(N__45070),
            .I(N__45066));
    CascadeMux I__8868 (
            .O(N__45069),
            .I(N__45063));
    InMux I__8867 (
            .O(N__45066),
            .I(N__45060));
    InMux I__8866 (
            .O(N__45063),
            .I(N__45057));
    LocalMux I__8865 (
            .O(N__45060),
            .I(\c0.data_in_frame_14_3 ));
    LocalMux I__8864 (
            .O(N__45057),
            .I(\c0.data_in_frame_14_3 ));
    InMux I__8863 (
            .O(N__45052),
            .I(N__45048));
    CascadeMux I__8862 (
            .O(N__45051),
            .I(N__45045));
    LocalMux I__8861 (
            .O(N__45048),
            .I(N__45042));
    InMux I__8860 (
            .O(N__45045),
            .I(N__45039));
    Span4Mux_h I__8859 (
            .O(N__45042),
            .I(N__45035));
    LocalMux I__8858 (
            .O(N__45039),
            .I(N__45032));
    InMux I__8857 (
            .O(N__45038),
            .I(N__45029));
    Odrv4 I__8856 (
            .O(N__45035),
            .I(\c0.n67_adj_3063 ));
    Odrv12 I__8855 (
            .O(N__45032),
            .I(\c0.n67_adj_3063 ));
    LocalMux I__8854 (
            .O(N__45029),
            .I(\c0.n67_adj_3063 ));
    CascadeMux I__8853 (
            .O(N__45022),
            .I(N__45017));
    InMux I__8852 (
            .O(N__45021),
            .I(N__45009));
    InMux I__8851 (
            .O(N__45020),
            .I(N__45009));
    InMux I__8850 (
            .O(N__45017),
            .I(N__45006));
    InMux I__8849 (
            .O(N__45016),
            .I(N__44999));
    InMux I__8848 (
            .O(N__45015),
            .I(N__44999));
    InMux I__8847 (
            .O(N__45014),
            .I(N__44999));
    LocalMux I__8846 (
            .O(N__45009),
            .I(N__44996));
    LocalMux I__8845 (
            .O(N__45006),
            .I(N__44991));
    LocalMux I__8844 (
            .O(N__44999),
            .I(N__44991));
    Odrv12 I__8843 (
            .O(N__44996),
            .I(\c0.n20490 ));
    Odrv4 I__8842 (
            .O(N__44991),
            .I(\c0.n20490 ));
    InMux I__8841 (
            .O(N__44986),
            .I(N__44980));
    InMux I__8840 (
            .O(N__44985),
            .I(N__44980));
    LocalMux I__8839 (
            .O(N__44980),
            .I(N__44976));
    InMux I__8838 (
            .O(N__44979),
            .I(N__44973));
    Span4Mux_v I__8837 (
            .O(N__44976),
            .I(N__44964));
    LocalMux I__8836 (
            .O(N__44973),
            .I(N__44964));
    InMux I__8835 (
            .O(N__44972),
            .I(N__44957));
    InMux I__8834 (
            .O(N__44971),
            .I(N__44957));
    InMux I__8833 (
            .O(N__44970),
            .I(N__44957));
    InMux I__8832 (
            .O(N__44969),
            .I(N__44954));
    Odrv4 I__8831 (
            .O(N__44964),
            .I(\c0.n19433 ));
    LocalMux I__8830 (
            .O(N__44957),
            .I(\c0.n19433 ));
    LocalMux I__8829 (
            .O(N__44954),
            .I(\c0.n19433 ));
    CascadeMux I__8828 (
            .O(N__44947),
            .I(N__44941));
    InMux I__8827 (
            .O(N__44946),
            .I(N__44938));
    InMux I__8826 (
            .O(N__44945),
            .I(N__44935));
    InMux I__8825 (
            .O(N__44944),
            .I(N__44932));
    InMux I__8824 (
            .O(N__44941),
            .I(N__44929));
    LocalMux I__8823 (
            .O(N__44938),
            .I(\c0.n42_adj_3064 ));
    LocalMux I__8822 (
            .O(N__44935),
            .I(\c0.n42_adj_3064 ));
    LocalMux I__8821 (
            .O(N__44932),
            .I(\c0.n42_adj_3064 ));
    LocalMux I__8820 (
            .O(N__44929),
            .I(\c0.n42_adj_3064 ));
    InMux I__8819 (
            .O(N__44920),
            .I(N__44917));
    LocalMux I__8818 (
            .O(N__44917),
            .I(N__44914));
    Span4Mux_v I__8817 (
            .O(N__44914),
            .I(N__44911));
    Odrv4 I__8816 (
            .O(N__44911),
            .I(\c0.n12_adj_3518 ));
    CascadeMux I__8815 (
            .O(N__44908),
            .I(\c0.n12_adj_3517_cascade_ ));
    CascadeMux I__8814 (
            .O(N__44905),
            .I(N__44901));
    CascadeMux I__8813 (
            .O(N__44904),
            .I(N__44898));
    InMux I__8812 (
            .O(N__44901),
            .I(N__44894));
    InMux I__8811 (
            .O(N__44898),
            .I(N__44889));
    InMux I__8810 (
            .O(N__44897),
            .I(N__44886));
    LocalMux I__8809 (
            .O(N__44894),
            .I(N__44883));
    InMux I__8808 (
            .O(N__44893),
            .I(N__44880));
    InMux I__8807 (
            .O(N__44892),
            .I(N__44877));
    LocalMux I__8806 (
            .O(N__44889),
            .I(N__44874));
    LocalMux I__8805 (
            .O(N__44886),
            .I(N__44871));
    Span4Mux_v I__8804 (
            .O(N__44883),
            .I(N__44868));
    LocalMux I__8803 (
            .O(N__44880),
            .I(N__44865));
    LocalMux I__8802 (
            .O(N__44877),
            .I(N__44860));
    Span4Mux_v I__8801 (
            .O(N__44874),
            .I(N__44860));
    Span4Mux_v I__8800 (
            .O(N__44871),
            .I(N__44855));
    Span4Mux_h I__8799 (
            .O(N__44868),
            .I(N__44855));
    Odrv4 I__8798 (
            .O(N__44865),
            .I(data_in_frame_18_5));
    Odrv4 I__8797 (
            .O(N__44860),
            .I(data_in_frame_18_5));
    Odrv4 I__8796 (
            .O(N__44855),
            .I(data_in_frame_18_5));
    InMux I__8795 (
            .O(N__44848),
            .I(N__44845));
    LocalMux I__8794 (
            .O(N__44845),
            .I(N__44842));
    Odrv4 I__8793 (
            .O(N__44842),
            .I(\c0.n21_adj_3337 ));
    CascadeMux I__8792 (
            .O(N__44839),
            .I(N__44836));
    InMux I__8791 (
            .O(N__44836),
            .I(N__44833));
    LocalMux I__8790 (
            .O(N__44833),
            .I(N__44830));
    Odrv12 I__8789 (
            .O(N__44830),
            .I(\c0.n20_adj_3487 ));
    InMux I__8788 (
            .O(N__44827),
            .I(N__44824));
    LocalMux I__8787 (
            .O(N__44824),
            .I(N__44821));
    Odrv4 I__8786 (
            .O(N__44821),
            .I(\c0.n18_adj_3369 ));
    CascadeMux I__8785 (
            .O(N__44818),
            .I(\c0.n19477_cascade_ ));
    CascadeMux I__8784 (
            .O(N__44815),
            .I(\c0.n12_adj_3348_cascade_ ));
    CascadeMux I__8783 (
            .O(N__44812),
            .I(\c0.n21045_cascade_ ));
    InMux I__8782 (
            .O(N__44809),
            .I(N__44806));
    LocalMux I__8781 (
            .O(N__44806),
            .I(N__44801));
    InMux I__8780 (
            .O(N__44805),
            .I(N__44798));
    InMux I__8779 (
            .O(N__44804),
            .I(N__44795));
    Odrv4 I__8778 (
            .O(N__44801),
            .I(\c0.n27_adj_3118 ));
    LocalMux I__8777 (
            .O(N__44798),
            .I(\c0.n27_adj_3118 ));
    LocalMux I__8776 (
            .O(N__44795),
            .I(\c0.n27_adj_3118 ));
    InMux I__8775 (
            .O(N__44788),
            .I(N__44785));
    LocalMux I__8774 (
            .O(N__44785),
            .I(N__44782));
    Span4Mux_v I__8773 (
            .O(N__44782),
            .I(N__44779));
    Span4Mux_h I__8772 (
            .O(N__44779),
            .I(N__44776));
    Span4Mux_v I__8771 (
            .O(N__44776),
            .I(N__44772));
    InMux I__8770 (
            .O(N__44775),
            .I(N__44769));
    Odrv4 I__8769 (
            .O(N__44772),
            .I(\c0.n19_adj_3303 ));
    LocalMux I__8768 (
            .O(N__44769),
            .I(\c0.n19_adj_3303 ));
    InMux I__8767 (
            .O(N__44764),
            .I(N__44761));
    LocalMux I__8766 (
            .O(N__44761),
            .I(N__44758));
    Span12Mux_v I__8765 (
            .O(N__44758),
            .I(N__44755));
    Odrv12 I__8764 (
            .O(N__44755),
            .I(\c0.n12 ));
    InMux I__8763 (
            .O(N__44752),
            .I(N__44749));
    LocalMux I__8762 (
            .O(N__44749),
            .I(N__44746));
    Odrv4 I__8761 (
            .O(N__44746),
            .I(\c0.n44_adj_3117 ));
    InMux I__8760 (
            .O(N__44743),
            .I(N__44740));
    LocalMux I__8759 (
            .O(N__44740),
            .I(\c0.n43_adj_3116 ));
    CascadeMux I__8758 (
            .O(N__44737),
            .I(\c0.n27_adj_3118_cascade_ ));
    InMux I__8757 (
            .O(N__44734),
            .I(N__44731));
    LocalMux I__8756 (
            .O(N__44731),
            .I(N__44727));
    InMux I__8755 (
            .O(N__44730),
            .I(N__44724));
    Odrv4 I__8754 (
            .O(N__44727),
            .I(\c0.n20052 ));
    LocalMux I__8753 (
            .O(N__44724),
            .I(\c0.n20052 ));
    InMux I__8752 (
            .O(N__44719),
            .I(N__44713));
    InMux I__8751 (
            .O(N__44718),
            .I(N__44707));
    InMux I__8750 (
            .O(N__44717),
            .I(N__44707));
    InMux I__8749 (
            .O(N__44716),
            .I(N__44704));
    LocalMux I__8748 (
            .O(N__44713),
            .I(N__44701));
    CascadeMux I__8747 (
            .O(N__44712),
            .I(N__44698));
    LocalMux I__8746 (
            .O(N__44707),
            .I(N__44693));
    LocalMux I__8745 (
            .O(N__44704),
            .I(N__44693));
    Span4Mux_v I__8744 (
            .O(N__44701),
            .I(N__44690));
    InMux I__8743 (
            .O(N__44698),
            .I(N__44687));
    Span4Mux_v I__8742 (
            .O(N__44693),
            .I(N__44684));
    Span4Mux_v I__8741 (
            .O(N__44690),
            .I(N__44681));
    LocalMux I__8740 (
            .O(N__44687),
            .I(N__44676));
    Span4Mux_v I__8739 (
            .O(N__44684),
            .I(N__44676));
    Odrv4 I__8738 (
            .O(N__44681),
            .I(\c0.data_in_frame_14_5 ));
    Odrv4 I__8737 (
            .O(N__44676),
            .I(\c0.data_in_frame_14_5 ));
    InMux I__8736 (
            .O(N__44671),
            .I(N__44668));
    LocalMux I__8735 (
            .O(N__44668),
            .I(N__44665));
    Odrv12 I__8734 (
            .O(N__44665),
            .I(\c0.n11_adj_3340 ));
    CascadeMux I__8733 (
            .O(N__44662),
            .I(\c0.n19916_cascade_ ));
    CascadeMux I__8732 (
            .O(N__44659),
            .I(N__44655));
    InMux I__8731 (
            .O(N__44658),
            .I(N__44651));
    InMux I__8730 (
            .O(N__44655),
            .I(N__44646));
    InMux I__8729 (
            .O(N__44654),
            .I(N__44646));
    LocalMux I__8728 (
            .O(N__44651),
            .I(\c0.n22_adj_3356 ));
    LocalMux I__8727 (
            .O(N__44646),
            .I(\c0.n22_adj_3356 ));
    InMux I__8726 (
            .O(N__44641),
            .I(N__44638));
    LocalMux I__8725 (
            .O(N__44638),
            .I(\c0.n22_adj_3022 ));
    CascadeMux I__8724 (
            .O(N__44635),
            .I(N__44628));
    CascadeMux I__8723 (
            .O(N__44634),
            .I(N__44625));
    InMux I__8722 (
            .O(N__44633),
            .I(N__44619));
    InMux I__8721 (
            .O(N__44632),
            .I(N__44619));
    InMux I__8720 (
            .O(N__44631),
            .I(N__44616));
    InMux I__8719 (
            .O(N__44628),
            .I(N__44613));
    InMux I__8718 (
            .O(N__44625),
            .I(N__44610));
    CascadeMux I__8717 (
            .O(N__44624),
            .I(N__44607));
    LocalMux I__8716 (
            .O(N__44619),
            .I(N__44602));
    LocalMux I__8715 (
            .O(N__44616),
            .I(N__44602));
    LocalMux I__8714 (
            .O(N__44613),
            .I(N__44597));
    LocalMux I__8713 (
            .O(N__44610),
            .I(N__44597));
    InMux I__8712 (
            .O(N__44607),
            .I(N__44594));
    Span4Mux_v I__8711 (
            .O(N__44602),
            .I(N__44589));
    Span4Mux_h I__8710 (
            .O(N__44597),
            .I(N__44589));
    LocalMux I__8709 (
            .O(N__44594),
            .I(\c0.data_in_frame_12_4 ));
    Odrv4 I__8708 (
            .O(N__44589),
            .I(\c0.data_in_frame_12_4 ));
    InMux I__8707 (
            .O(N__44584),
            .I(N__44581));
    LocalMux I__8706 (
            .O(N__44581),
            .I(N__44578));
    Span4Mux_v I__8705 (
            .O(N__44578),
            .I(N__44575));
    Odrv4 I__8704 (
            .O(N__44575),
            .I(\c0.n18_adj_3372 ));
    InMux I__8703 (
            .O(N__44572),
            .I(N__44568));
    CascadeMux I__8702 (
            .O(N__44571),
            .I(N__44565));
    LocalMux I__8701 (
            .O(N__44568),
            .I(N__44562));
    InMux I__8700 (
            .O(N__44565),
            .I(N__44559));
    Odrv4 I__8699 (
            .O(N__44562),
            .I(\c0.n88 ));
    LocalMux I__8698 (
            .O(N__44559),
            .I(\c0.n88 ));
    CascadeMux I__8697 (
            .O(N__44554),
            .I(N__44551));
    InMux I__8696 (
            .O(N__44551),
            .I(N__44548));
    LocalMux I__8695 (
            .O(N__44548),
            .I(\c0.n33 ));
    InMux I__8694 (
            .O(N__44545),
            .I(N__44542));
    LocalMux I__8693 (
            .O(N__44542),
            .I(N__44539));
    Span4Mux_h I__8692 (
            .O(N__44539),
            .I(N__44535));
    InMux I__8691 (
            .O(N__44538),
            .I(N__44532));
    Odrv4 I__8690 (
            .O(N__44535),
            .I(\c0.n20029 ));
    LocalMux I__8689 (
            .O(N__44532),
            .I(\c0.n20029 ));
    InMux I__8688 (
            .O(N__44527),
            .I(N__44524));
    LocalMux I__8687 (
            .O(N__44524),
            .I(\c0.n26_adj_3114 ));
    CascadeMux I__8686 (
            .O(N__44521),
            .I(N__44518));
    InMux I__8685 (
            .O(N__44518),
            .I(N__44514));
    InMux I__8684 (
            .O(N__44517),
            .I(N__44511));
    LocalMux I__8683 (
            .O(N__44514),
            .I(\c0.n30 ));
    LocalMux I__8682 (
            .O(N__44511),
            .I(\c0.n30 ));
    InMux I__8681 (
            .O(N__44506),
            .I(N__44503));
    LocalMux I__8680 (
            .O(N__44503),
            .I(N__44500));
    Span4Mux_h I__8679 (
            .O(N__44500),
            .I(N__44496));
    InMux I__8678 (
            .O(N__44499),
            .I(N__44493));
    Odrv4 I__8677 (
            .O(N__44496),
            .I(\c0.n18422 ));
    LocalMux I__8676 (
            .O(N__44493),
            .I(\c0.n18422 ));
    CascadeMux I__8675 (
            .O(N__44488),
            .I(\c0.n18422_cascade_ ));
    CascadeMux I__8674 (
            .O(N__44485),
            .I(\c0.n19433_cascade_ ));
    CascadeMux I__8673 (
            .O(N__44482),
            .I(N__44476));
    CascadeMux I__8672 (
            .O(N__44481),
            .I(N__44473));
    CascadeMux I__8671 (
            .O(N__44480),
            .I(N__44469));
    InMux I__8670 (
            .O(N__44479),
            .I(N__44466));
    InMux I__8669 (
            .O(N__44476),
            .I(N__44462));
    InMux I__8668 (
            .O(N__44473),
            .I(N__44459));
    InMux I__8667 (
            .O(N__44472),
            .I(N__44454));
    InMux I__8666 (
            .O(N__44469),
            .I(N__44454));
    LocalMux I__8665 (
            .O(N__44466),
            .I(N__44451));
    InMux I__8664 (
            .O(N__44465),
            .I(N__44448));
    LocalMux I__8663 (
            .O(N__44462),
            .I(N__44445));
    LocalMux I__8662 (
            .O(N__44459),
            .I(\c0.data_in_frame_10_3 ));
    LocalMux I__8661 (
            .O(N__44454),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__8660 (
            .O(N__44451),
            .I(\c0.data_in_frame_10_3 ));
    LocalMux I__8659 (
            .O(N__44448),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__8658 (
            .O(N__44445),
            .I(\c0.data_in_frame_10_3 ));
    CascadeMux I__8657 (
            .O(N__44434),
            .I(\c0.n11891_cascade_ ));
    InMux I__8656 (
            .O(N__44431),
            .I(N__44428));
    LocalMux I__8655 (
            .O(N__44428),
            .I(\c0.n14_adj_3371 ));
    InMux I__8654 (
            .O(N__44425),
            .I(N__44420));
    CascadeMux I__8653 (
            .O(N__44424),
            .I(N__44417));
    CascadeMux I__8652 (
            .O(N__44423),
            .I(N__44414));
    LocalMux I__8651 (
            .O(N__44420),
            .I(N__44410));
    InMux I__8650 (
            .O(N__44417),
            .I(N__44403));
    InMux I__8649 (
            .O(N__44414),
            .I(N__44403));
    InMux I__8648 (
            .O(N__44413),
            .I(N__44403));
    Odrv4 I__8647 (
            .O(N__44410),
            .I(\c0.data_in_frame_3_6 ));
    LocalMux I__8646 (
            .O(N__44403),
            .I(\c0.data_in_frame_3_6 ));
    CascadeMux I__8645 (
            .O(N__44398),
            .I(\c0.n10_adj_3538_cascade_ ));
    CascadeMux I__8644 (
            .O(N__44395),
            .I(N__44390));
    InMux I__8643 (
            .O(N__44394),
            .I(N__44387));
    CascadeMux I__8642 (
            .O(N__44393),
            .I(N__44384));
    InMux I__8641 (
            .O(N__44390),
            .I(N__44379));
    LocalMux I__8640 (
            .O(N__44387),
            .I(N__44376));
    InMux I__8639 (
            .O(N__44384),
            .I(N__44373));
    InMux I__8638 (
            .O(N__44383),
            .I(N__44368));
    InMux I__8637 (
            .O(N__44382),
            .I(N__44368));
    LocalMux I__8636 (
            .O(N__44379),
            .I(\c0.data_in_frame_2_5 ));
    Odrv12 I__8635 (
            .O(N__44376),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__8634 (
            .O(N__44373),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__8633 (
            .O(N__44368),
            .I(\c0.data_in_frame_2_5 ));
    CascadeMux I__8632 (
            .O(N__44359),
            .I(\c0.n22_adj_3356_cascade_ ));
    InMux I__8631 (
            .O(N__44356),
            .I(N__44352));
    InMux I__8630 (
            .O(N__44355),
            .I(N__44349));
    LocalMux I__8629 (
            .O(N__44352),
            .I(\c0.n13_adj_3513 ));
    LocalMux I__8628 (
            .O(N__44349),
            .I(\c0.n13_adj_3513 ));
    CascadeMux I__8627 (
            .O(N__44344),
            .I(N__44341));
    InMux I__8626 (
            .O(N__44341),
            .I(N__44338));
    LocalMux I__8625 (
            .O(N__44338),
            .I(\c0.n23_adj_3021 ));
    CascadeMux I__8624 (
            .O(N__44335),
            .I(\c0.n23_adj_3021_cascade_ ));
    CascadeMux I__8623 (
            .O(N__44332),
            .I(\c0.n26_adj_3114_cascade_ ));
    InMux I__8622 (
            .O(N__44329),
            .I(N__44323));
    InMux I__8621 (
            .O(N__44328),
            .I(N__44323));
    LocalMux I__8620 (
            .O(N__44323),
            .I(\c0.n24_adj_3011 ));
    InMux I__8619 (
            .O(N__44320),
            .I(N__44317));
    LocalMux I__8618 (
            .O(N__44317),
            .I(N__44314));
    Odrv4 I__8617 (
            .O(N__44314),
            .I(\c0.n22 ));
    InMux I__8616 (
            .O(N__44311),
            .I(N__44305));
    InMux I__8615 (
            .O(N__44310),
            .I(N__44305));
    LocalMux I__8614 (
            .O(N__44305),
            .I(N__44301));
    InMux I__8613 (
            .O(N__44304),
            .I(N__44298));
    Odrv12 I__8612 (
            .O(N__44301),
            .I(\c0.n12131 ));
    LocalMux I__8611 (
            .O(N__44298),
            .I(\c0.n12131 ));
    InMux I__8610 (
            .O(N__44293),
            .I(N__44287));
    InMux I__8609 (
            .O(N__44292),
            .I(N__44287));
    LocalMux I__8608 (
            .O(N__44287),
            .I(\c0.n19415 ));
    CascadeMux I__8607 (
            .O(N__44284),
            .I(\c0.n19415_cascade_ ));
    InMux I__8606 (
            .O(N__44281),
            .I(N__44275));
    InMux I__8605 (
            .O(N__44280),
            .I(N__44275));
    LocalMux I__8604 (
            .O(N__44275),
            .I(\c0.n54_adj_3502 ));
    InMux I__8603 (
            .O(N__44272),
            .I(N__44268));
    InMux I__8602 (
            .O(N__44271),
            .I(N__44265));
    LocalMux I__8601 (
            .O(N__44268),
            .I(\c0.n39_adj_3398 ));
    LocalMux I__8600 (
            .O(N__44265),
            .I(\c0.n39_adj_3398 ));
    InMux I__8599 (
            .O(N__44260),
            .I(N__44257));
    LocalMux I__8598 (
            .O(N__44257),
            .I(N__44254));
    Span4Mux_h I__8597 (
            .O(N__44254),
            .I(N__44249));
    CascadeMux I__8596 (
            .O(N__44253),
            .I(N__44244));
    InMux I__8595 (
            .O(N__44252),
            .I(N__44241));
    Span4Mux_v I__8594 (
            .O(N__44249),
            .I(N__44237));
    InMux I__8593 (
            .O(N__44248),
            .I(N__44234));
    InMux I__8592 (
            .O(N__44247),
            .I(N__44230));
    InMux I__8591 (
            .O(N__44244),
            .I(N__44227));
    LocalMux I__8590 (
            .O(N__44241),
            .I(N__44224));
    InMux I__8589 (
            .O(N__44240),
            .I(N__44221));
    Span4Mux_v I__8588 (
            .O(N__44237),
            .I(N__44217));
    LocalMux I__8587 (
            .O(N__44234),
            .I(N__44212));
    InMux I__8586 (
            .O(N__44233),
            .I(N__44209));
    LocalMux I__8585 (
            .O(N__44230),
            .I(N__44206));
    LocalMux I__8584 (
            .O(N__44227),
            .I(N__44199));
    Span4Mux_h I__8583 (
            .O(N__44224),
            .I(N__44199));
    LocalMux I__8582 (
            .O(N__44221),
            .I(N__44199));
    InMux I__8581 (
            .O(N__44220),
            .I(N__44196));
    Span4Mux_v I__8580 (
            .O(N__44217),
            .I(N__44193));
    InMux I__8579 (
            .O(N__44216),
            .I(N__44188));
    InMux I__8578 (
            .O(N__44215),
            .I(N__44188));
    Span12Mux_h I__8577 (
            .O(N__44212),
            .I(N__44185));
    LocalMux I__8576 (
            .O(N__44209),
            .I(N__44180));
    Span4Mux_v I__8575 (
            .O(N__44206),
            .I(N__44180));
    Span4Mux_v I__8574 (
            .O(N__44199),
            .I(N__44177));
    LocalMux I__8573 (
            .O(N__44196),
            .I(N__44174));
    Span4Mux_h I__8572 (
            .O(N__44193),
            .I(N__44171));
    LocalMux I__8571 (
            .O(N__44188),
            .I(\c0.n9_adj_3025 ));
    Odrv12 I__8570 (
            .O(N__44185),
            .I(\c0.n9_adj_3025 ));
    Odrv4 I__8569 (
            .O(N__44180),
            .I(\c0.n9_adj_3025 ));
    Odrv4 I__8568 (
            .O(N__44177),
            .I(\c0.n9_adj_3025 ));
    Odrv12 I__8567 (
            .O(N__44174),
            .I(\c0.n9_adj_3025 ));
    Odrv4 I__8566 (
            .O(N__44171),
            .I(\c0.n9_adj_3025 ));
    InMux I__8565 (
            .O(N__44158),
            .I(N__44152));
    InMux I__8564 (
            .O(N__44157),
            .I(N__44148));
    InMux I__8563 (
            .O(N__44156),
            .I(N__44143));
    InMux I__8562 (
            .O(N__44155),
            .I(N__44143));
    LocalMux I__8561 (
            .O(N__44152),
            .I(N__44140));
    InMux I__8560 (
            .O(N__44151),
            .I(N__44137));
    LocalMux I__8559 (
            .O(N__44148),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__8558 (
            .O(N__44143),
            .I(\c0.data_in_frame_2_7 ));
    Odrv12 I__8557 (
            .O(N__44140),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__8556 (
            .O(N__44137),
            .I(\c0.data_in_frame_2_7 ));
    CascadeMux I__8555 (
            .O(N__44128),
            .I(N__44121));
    InMux I__8554 (
            .O(N__44127),
            .I(N__44114));
    InMux I__8553 (
            .O(N__44126),
            .I(N__44109));
    InMux I__8552 (
            .O(N__44125),
            .I(N__44109));
    InMux I__8551 (
            .O(N__44124),
            .I(N__44102));
    InMux I__8550 (
            .O(N__44121),
            .I(N__44102));
    InMux I__8549 (
            .O(N__44120),
            .I(N__44102));
    InMux I__8548 (
            .O(N__44119),
            .I(N__44099));
    InMux I__8547 (
            .O(N__44118),
            .I(N__44094));
    InMux I__8546 (
            .O(N__44117),
            .I(N__44094));
    LocalMux I__8545 (
            .O(N__44114),
            .I(N__44091));
    LocalMux I__8544 (
            .O(N__44109),
            .I(N__44088));
    LocalMux I__8543 (
            .O(N__44102),
            .I(N__44083));
    LocalMux I__8542 (
            .O(N__44099),
            .I(N__44083));
    LocalMux I__8541 (
            .O(N__44094),
            .I(N__44080));
    Span4Mux_v I__8540 (
            .O(N__44091),
            .I(N__44077));
    Span4Mux_v I__8539 (
            .O(N__44088),
            .I(N__44072));
    Span4Mux_v I__8538 (
            .O(N__44083),
            .I(N__44072));
    Span4Mux_h I__8537 (
            .O(N__44080),
            .I(N__44069));
    Span4Mux_h I__8536 (
            .O(N__44077),
            .I(N__44066));
    Span4Mux_h I__8535 (
            .O(N__44072),
            .I(N__44063));
    Span4Mux_h I__8534 (
            .O(N__44069),
            .I(N__44058));
    Span4Mux_v I__8533 (
            .O(N__44066),
            .I(N__44058));
    Odrv4 I__8532 (
            .O(N__44063),
            .I(\c0.n9_adj_3351 ));
    Odrv4 I__8531 (
            .O(N__44058),
            .I(\c0.n9_adj_3351 ));
    CascadeMux I__8530 (
            .O(N__44053),
            .I(N__44050));
    InMux I__8529 (
            .O(N__44050),
            .I(N__44042));
    InMux I__8528 (
            .O(N__44049),
            .I(N__44042));
    InMux I__8527 (
            .O(N__44048),
            .I(N__44039));
    CascadeMux I__8526 (
            .O(N__44047),
            .I(N__44036));
    LocalMux I__8525 (
            .O(N__44042),
            .I(N__44031));
    LocalMux I__8524 (
            .O(N__44039),
            .I(N__44031));
    InMux I__8523 (
            .O(N__44036),
            .I(N__44025));
    Span4Mux_h I__8522 (
            .O(N__44031),
            .I(N__44022));
    InMux I__8521 (
            .O(N__44030),
            .I(N__44019));
    InMux I__8520 (
            .O(N__44029),
            .I(N__44014));
    InMux I__8519 (
            .O(N__44028),
            .I(N__44014));
    LocalMux I__8518 (
            .O(N__44025),
            .I(\c0.data_in_frame_4_6 ));
    Odrv4 I__8517 (
            .O(N__44022),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__8516 (
            .O(N__44019),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__8515 (
            .O(N__44014),
            .I(\c0.data_in_frame_4_6 ));
    InMux I__8514 (
            .O(N__44005),
            .I(N__44002));
    LocalMux I__8513 (
            .O(N__44002),
            .I(N__43999));
    Span4Mux_h I__8512 (
            .O(N__43999),
            .I(N__43996));
    Odrv4 I__8511 (
            .O(N__43996),
            .I(\c0.n11_adj_3507 ));
    CascadeMux I__8510 (
            .O(N__43993),
            .I(N__43990));
    InMux I__8509 (
            .O(N__43990),
            .I(N__43987));
    LocalMux I__8508 (
            .O(N__43987),
            .I(\c0.n13_adj_3504 ));
    CascadeMux I__8507 (
            .O(N__43984),
            .I(\c0.n12131_cascade_ ));
    InMux I__8506 (
            .O(N__43981),
            .I(N__43978));
    LocalMux I__8505 (
            .O(N__43978),
            .I(N__43975));
    Span4Mux_h I__8504 (
            .O(N__43975),
            .I(N__43969));
    InMux I__8503 (
            .O(N__43974),
            .I(N__43966));
    InMux I__8502 (
            .O(N__43973),
            .I(N__43961));
    InMux I__8501 (
            .O(N__43972),
            .I(N__43961));
    Odrv4 I__8500 (
            .O(N__43969),
            .I(data_in_3_4));
    LocalMux I__8499 (
            .O(N__43966),
            .I(data_in_3_4));
    LocalMux I__8498 (
            .O(N__43961),
            .I(data_in_3_4));
    InMux I__8497 (
            .O(N__43954),
            .I(N__43950));
    InMux I__8496 (
            .O(N__43953),
            .I(N__43947));
    LocalMux I__8495 (
            .O(N__43950),
            .I(data_in_0_0));
    LocalMux I__8494 (
            .O(N__43947),
            .I(data_in_0_0));
    InMux I__8493 (
            .O(N__43942),
            .I(N__43937));
    InMux I__8492 (
            .O(N__43941),
            .I(N__43934));
    InMux I__8491 (
            .O(N__43940),
            .I(N__43931));
    LocalMux I__8490 (
            .O(N__43937),
            .I(data_in_1_7));
    LocalMux I__8489 (
            .O(N__43934),
            .I(data_in_1_7));
    LocalMux I__8488 (
            .O(N__43931),
            .I(data_in_1_7));
    InMux I__8487 (
            .O(N__43924),
            .I(N__43918));
    InMux I__8486 (
            .O(N__43923),
            .I(N__43918));
    LocalMux I__8485 (
            .O(N__43918),
            .I(\c0.n10_adj_3231 ));
    InMux I__8484 (
            .O(N__43915),
            .I(N__43912));
    LocalMux I__8483 (
            .O(N__43912),
            .I(N__43909));
    Span4Mux_v I__8482 (
            .O(N__43909),
            .I(N__43903));
    InMux I__8481 (
            .O(N__43908),
            .I(N__43898));
    InMux I__8480 (
            .O(N__43907),
            .I(N__43898));
    InMux I__8479 (
            .O(N__43906),
            .I(N__43895));
    Odrv4 I__8478 (
            .O(N__43903),
            .I(data_in_2_1));
    LocalMux I__8477 (
            .O(N__43898),
            .I(data_in_2_1));
    LocalMux I__8476 (
            .O(N__43895),
            .I(data_in_2_1));
    InMux I__8475 (
            .O(N__43888),
            .I(N__43883));
    InMux I__8474 (
            .O(N__43887),
            .I(N__43880));
    InMux I__8473 (
            .O(N__43886),
            .I(N__43877));
    LocalMux I__8472 (
            .O(N__43883),
            .I(data_in_1_1));
    LocalMux I__8471 (
            .O(N__43880),
            .I(data_in_1_1));
    LocalMux I__8470 (
            .O(N__43877),
            .I(data_in_1_1));
    InMux I__8469 (
            .O(N__43870),
            .I(N__43866));
    InMux I__8468 (
            .O(N__43869),
            .I(N__43863));
    LocalMux I__8467 (
            .O(N__43866),
            .I(N__43860));
    LocalMux I__8466 (
            .O(N__43863),
            .I(N__43856));
    Span4Mux_v I__8465 (
            .O(N__43860),
            .I(N__43853));
    InMux I__8464 (
            .O(N__43859),
            .I(N__43850));
    Span4Mux_h I__8463 (
            .O(N__43856),
            .I(N__43846));
    Sp12to4 I__8462 (
            .O(N__43853),
            .I(N__43841));
    LocalMux I__8461 (
            .O(N__43850),
            .I(N__43841));
    InMux I__8460 (
            .O(N__43849),
            .I(N__43836));
    Sp12to4 I__8459 (
            .O(N__43846),
            .I(N__43831));
    Span12Mux_h I__8458 (
            .O(N__43841),
            .I(N__43831));
    InMux I__8457 (
            .O(N__43840),
            .I(N__43826));
    InMux I__8456 (
            .O(N__43839),
            .I(N__43826));
    LocalMux I__8455 (
            .O(N__43836),
            .I(r_Bit_Index_2));
    Odrv12 I__8454 (
            .O(N__43831),
            .I(r_Bit_Index_2));
    LocalMux I__8453 (
            .O(N__43826),
            .I(r_Bit_Index_2));
    InMux I__8452 (
            .O(N__43819),
            .I(N__43814));
    InMux I__8451 (
            .O(N__43818),
            .I(N__43811));
    InMux I__8450 (
            .O(N__43817),
            .I(N__43808));
    LocalMux I__8449 (
            .O(N__43814),
            .I(N__43805));
    LocalMux I__8448 (
            .O(N__43811),
            .I(N__43802));
    LocalMux I__8447 (
            .O(N__43808),
            .I(N__43794));
    Span4Mux_h I__8446 (
            .O(N__43805),
            .I(N__43794));
    Sp12to4 I__8445 (
            .O(N__43802),
            .I(N__43791));
    InMux I__8444 (
            .O(N__43801),
            .I(N__43783));
    InMux I__8443 (
            .O(N__43800),
            .I(N__43783));
    InMux I__8442 (
            .O(N__43799),
            .I(N__43783));
    Sp12to4 I__8441 (
            .O(N__43794),
            .I(N__43778));
    Span12Mux_s7_v I__8440 (
            .O(N__43791),
            .I(N__43778));
    InMux I__8439 (
            .O(N__43790),
            .I(N__43775));
    LocalMux I__8438 (
            .O(N__43783),
            .I(N__43772));
    Span12Mux_v I__8437 (
            .O(N__43778),
            .I(N__43769));
    LocalMux I__8436 (
            .O(N__43775),
            .I(r_Bit_Index_1));
    Odrv12 I__8435 (
            .O(N__43772),
            .I(r_Bit_Index_1));
    Odrv12 I__8434 (
            .O(N__43769),
            .I(r_Bit_Index_1));
    InMux I__8433 (
            .O(N__43762),
            .I(N__43759));
    LocalMux I__8432 (
            .O(N__43759),
            .I(N__43756));
    Span4Mux_h I__8431 (
            .O(N__43756),
            .I(N__43752));
    InMux I__8430 (
            .O(N__43755),
            .I(N__43749));
    Odrv4 I__8429 (
            .O(N__43752),
            .I(n4));
    LocalMux I__8428 (
            .O(N__43749),
            .I(n4));
    InMux I__8427 (
            .O(N__43744),
            .I(N__43738));
    InMux I__8426 (
            .O(N__43743),
            .I(N__43738));
    LocalMux I__8425 (
            .O(N__43738),
            .I(N__43735));
    Span4Mux_h I__8424 (
            .O(N__43735),
            .I(N__43732));
    Odrv4 I__8423 (
            .O(N__43732),
            .I(n4_adj_3579));
    CascadeMux I__8422 (
            .O(N__43729),
            .I(\c0.n15_adj_3297_cascade_ ));
    InMux I__8421 (
            .O(N__43726),
            .I(N__43723));
    LocalMux I__8420 (
            .O(N__43723),
            .I(\c0.n21003 ));
    CascadeMux I__8419 (
            .O(N__43720),
            .I(\c0.n21_adj_3300_cascade_ ));
    InMux I__8418 (
            .O(N__43717),
            .I(N__43714));
    LocalMux I__8417 (
            .O(N__43714),
            .I(\c0.n23_adj_3304 ));
    CascadeMux I__8416 (
            .O(N__43711),
            .I(\c0.n21247_cascade_ ));
    InMux I__8415 (
            .O(N__43708),
            .I(N__43705));
    LocalMux I__8414 (
            .O(N__43705),
            .I(\c0.n24_adj_3298 ));
    InMux I__8413 (
            .O(N__43702),
            .I(N__43699));
    LocalMux I__8412 (
            .O(N__43699),
            .I(\c0.n14_adj_3354 ));
    InMux I__8411 (
            .O(N__43696),
            .I(N__43690));
    InMux I__8410 (
            .O(N__43695),
            .I(N__43690));
    LocalMux I__8409 (
            .O(N__43690),
            .I(\c0.n34 ));
    CascadeMux I__8408 (
            .O(N__43687),
            .I(N__43684));
    InMux I__8407 (
            .O(N__43684),
            .I(N__43681));
    LocalMux I__8406 (
            .O(N__43681),
            .I(\c0.n19403 ));
    CascadeMux I__8405 (
            .O(N__43678),
            .I(N__43674));
    InMux I__8404 (
            .O(N__43677),
            .I(N__43669));
    InMux I__8403 (
            .O(N__43674),
            .I(N__43669));
    LocalMux I__8402 (
            .O(N__43669),
            .I(N__43665));
    InMux I__8401 (
            .O(N__43668),
            .I(N__43662));
    Span4Mux_v I__8400 (
            .O(N__43665),
            .I(N__43659));
    LocalMux I__8399 (
            .O(N__43662),
            .I(\c0.data_in_frame_26_6 ));
    Odrv4 I__8398 (
            .O(N__43659),
            .I(\c0.data_in_frame_26_6 ));
    CascadeMux I__8397 (
            .O(N__43654),
            .I(N__43651));
    InMux I__8396 (
            .O(N__43651),
            .I(N__43648));
    LocalMux I__8395 (
            .O(N__43648),
            .I(\c0.n38_adj_3051 ));
    CascadeMux I__8394 (
            .O(N__43645),
            .I(\c0.n38_adj_3051_cascade_ ));
    InMux I__8393 (
            .O(N__43642),
            .I(N__43638));
    InMux I__8392 (
            .O(N__43641),
            .I(N__43635));
    LocalMux I__8391 (
            .O(N__43638),
            .I(N__43632));
    LocalMux I__8390 (
            .O(N__43635),
            .I(\c0.n19496 ));
    Odrv4 I__8389 (
            .O(N__43632),
            .I(\c0.n19496 ));
    InMux I__8388 (
            .O(N__43627),
            .I(N__43624));
    LocalMux I__8387 (
            .O(N__43624),
            .I(N__43621));
    Odrv4 I__8386 (
            .O(N__43621),
            .I(\c0.n17947 ));
    InMux I__8385 (
            .O(N__43618),
            .I(N__43614));
    InMux I__8384 (
            .O(N__43617),
            .I(N__43611));
    LocalMux I__8383 (
            .O(N__43614),
            .I(N__43606));
    LocalMux I__8382 (
            .O(N__43611),
            .I(N__43606));
    Span4Mux_v I__8381 (
            .O(N__43606),
            .I(N__43603));
    Odrv4 I__8380 (
            .O(N__43603),
            .I(\c0.n60_adj_3065 ));
    InMux I__8379 (
            .O(N__43600),
            .I(N__43597));
    LocalMux I__8378 (
            .O(N__43597),
            .I(N__43594));
    Span4Mux_v I__8377 (
            .O(N__43594),
            .I(N__43591));
    Odrv4 I__8376 (
            .O(N__43591),
            .I(\c0.n64 ));
    CascadeMux I__8375 (
            .O(N__43588),
            .I(\c0.n51_cascade_ ));
    InMux I__8374 (
            .O(N__43585),
            .I(N__43579));
    InMux I__8373 (
            .O(N__43584),
            .I(N__43579));
    LocalMux I__8372 (
            .O(N__43579),
            .I(\c0.n32_adj_3052 ));
    InMux I__8371 (
            .O(N__43576),
            .I(N__43573));
    LocalMux I__8370 (
            .O(N__43573),
            .I(\c0.n45_adj_3284 ));
    CascadeMux I__8369 (
            .O(N__43570),
            .I(N__43567));
    InMux I__8368 (
            .O(N__43567),
            .I(N__43564));
    LocalMux I__8367 (
            .O(N__43564),
            .I(\c0.n40_adj_3282 ));
    InMux I__8366 (
            .O(N__43561),
            .I(N__43558));
    LocalMux I__8365 (
            .O(N__43558),
            .I(\c0.n20930 ));
    InMux I__8364 (
            .O(N__43555),
            .I(N__43551));
    InMux I__8363 (
            .O(N__43554),
            .I(N__43548));
    LocalMux I__8362 (
            .O(N__43551),
            .I(N__43544));
    LocalMux I__8361 (
            .O(N__43548),
            .I(N__43541));
    InMux I__8360 (
            .O(N__43547),
            .I(N__43538));
    Odrv4 I__8359 (
            .O(N__43544),
            .I(\c0.n19342 ));
    Odrv12 I__8358 (
            .O(N__43541),
            .I(\c0.n19342 ));
    LocalMux I__8357 (
            .O(N__43538),
            .I(\c0.n19342 ));
    CascadeMux I__8356 (
            .O(N__43531),
            .I(\c0.n36_adj_3307_cascade_ ));
    InMux I__8355 (
            .O(N__43528),
            .I(N__43525));
    LocalMux I__8354 (
            .O(N__43525),
            .I(\c0.n39_adj_3312 ));
    InMux I__8353 (
            .O(N__43522),
            .I(N__43517));
    InMux I__8352 (
            .O(N__43521),
            .I(N__43514));
    InMux I__8351 (
            .O(N__43520),
            .I(N__43511));
    LocalMux I__8350 (
            .O(N__43517),
            .I(N__43506));
    LocalMux I__8349 (
            .O(N__43514),
            .I(N__43506));
    LocalMux I__8348 (
            .O(N__43511),
            .I(N__43503));
    Span4Mux_v I__8347 (
            .O(N__43506),
            .I(N__43498));
    Span4Mux_v I__8346 (
            .O(N__43503),
            .I(N__43498));
    Odrv4 I__8345 (
            .O(N__43498),
            .I(\c0.n29_adj_3148 ));
    InMux I__8344 (
            .O(N__43495),
            .I(N__43492));
    LocalMux I__8343 (
            .O(N__43492),
            .I(\c0.n78_adj_3357 ));
    CascadeMux I__8342 (
            .O(N__43489),
            .I(\c0.n75_cascade_ ));
    CascadeMux I__8341 (
            .O(N__43486),
            .I(\c0.n93_adj_3373_cascade_ ));
    InMux I__8340 (
            .O(N__43483),
            .I(N__43480));
    LocalMux I__8339 (
            .O(N__43480),
            .I(N__43477));
    Odrv4 I__8338 (
            .O(N__43477),
            .I(\c0.n96_adj_3419 ));
    CascadeMux I__8337 (
            .O(N__43474),
            .I(\c0.n23_adj_3222_cascade_ ));
    InMux I__8336 (
            .O(N__43471),
            .I(N__43468));
    LocalMux I__8335 (
            .O(N__43468),
            .I(\c0.n76 ));
    CascadeMux I__8334 (
            .O(N__43465),
            .I(N__43462));
    InMux I__8333 (
            .O(N__43462),
            .I(N__43459));
    LocalMux I__8332 (
            .O(N__43459),
            .I(N__43456));
    Span12Mux_v I__8331 (
            .O(N__43456),
            .I(N__43451));
    InMux I__8330 (
            .O(N__43455),
            .I(N__43446));
    InMux I__8329 (
            .O(N__43454),
            .I(N__43446));
    Odrv12 I__8328 (
            .O(N__43451),
            .I(encoder0_position_31));
    LocalMux I__8327 (
            .O(N__43446),
            .I(encoder0_position_31));
    InMux I__8326 (
            .O(N__43441),
            .I(N__43438));
    LocalMux I__8325 (
            .O(N__43438),
            .I(N__43435));
    Span4Mux_h I__8324 (
            .O(N__43435),
            .I(N__43431));
    InMux I__8323 (
            .O(N__43434),
            .I(N__43428));
    Span4Mux_v I__8322 (
            .O(N__43431),
            .I(N__43425));
    LocalMux I__8321 (
            .O(N__43428),
            .I(data_out_frame_6_7));
    Odrv4 I__8320 (
            .O(N__43425),
            .I(data_out_frame_6_7));
    CascadeMux I__8319 (
            .O(N__43420),
            .I(N__43416));
    InMux I__8318 (
            .O(N__43419),
            .I(N__43411));
    InMux I__8317 (
            .O(N__43416),
            .I(N__43411));
    LocalMux I__8316 (
            .O(N__43411),
            .I(N__43407));
    InMux I__8315 (
            .O(N__43410),
            .I(N__43404));
    Span4Mux_v I__8314 (
            .O(N__43407),
            .I(N__43401));
    LocalMux I__8313 (
            .O(N__43404),
            .I(data_in_frame_23_2));
    Odrv4 I__8312 (
            .O(N__43401),
            .I(data_in_frame_23_2));
    CascadeMux I__8311 (
            .O(N__43396),
            .I(\c0.n13_adj_3405_cascade_ ));
    CascadeMux I__8310 (
            .O(N__43393),
            .I(N__43390));
    InMux I__8309 (
            .O(N__43390),
            .I(N__43386));
    InMux I__8308 (
            .O(N__43389),
            .I(N__43382));
    LocalMux I__8307 (
            .O(N__43386),
            .I(N__43379));
    InMux I__8306 (
            .O(N__43385),
            .I(N__43376));
    LocalMux I__8305 (
            .O(N__43382),
            .I(N__43373));
    Span4Mux_v I__8304 (
            .O(N__43379),
            .I(N__43370));
    LocalMux I__8303 (
            .O(N__43376),
            .I(\c0.data_in_frame_27_0 ));
    Odrv4 I__8302 (
            .O(N__43373),
            .I(\c0.data_in_frame_27_0 ));
    Odrv4 I__8301 (
            .O(N__43370),
            .I(\c0.data_in_frame_27_0 ));
    CascadeMux I__8300 (
            .O(N__43363),
            .I(\c0.n17880_cascade_ ));
    CascadeMux I__8299 (
            .O(N__43360),
            .I(\c0.n19342_cascade_ ));
    InMux I__8298 (
            .O(N__43357),
            .I(N__43354));
    LocalMux I__8297 (
            .O(N__43354),
            .I(\c0.n12035 ));
    CascadeMux I__8296 (
            .O(N__43351),
            .I(\c0.n19496_cascade_ ));
    InMux I__8295 (
            .O(N__43348),
            .I(N__43345));
    LocalMux I__8294 (
            .O(N__43345),
            .I(N__43342));
    Span4Mux_h I__8293 (
            .O(N__43342),
            .I(N__43339));
    Odrv4 I__8292 (
            .O(N__43339),
            .I(\c0.n15_adj_3395 ));
    CascadeMux I__8291 (
            .O(N__43336),
            .I(\c0.n15489_cascade_ ));
    InMux I__8290 (
            .O(N__43333),
            .I(N__43329));
    InMux I__8289 (
            .O(N__43332),
            .I(N__43326));
    LocalMux I__8288 (
            .O(N__43329),
            .I(\c0.data_in_frame_15_2 ));
    LocalMux I__8287 (
            .O(N__43326),
            .I(\c0.data_in_frame_15_2 ));
    CascadeMux I__8286 (
            .O(N__43321),
            .I(\c0.n20801_cascade_ ));
    CascadeMux I__8285 (
            .O(N__43318),
            .I(\c0.n96_adj_3401_cascade_ ));
    InMux I__8284 (
            .O(N__43315),
            .I(N__43312));
    LocalMux I__8283 (
            .O(N__43312),
            .I(N__43309));
    Span4Mux_v I__8282 (
            .O(N__43309),
            .I(N__43306));
    Odrv4 I__8281 (
            .O(N__43306),
            .I(\c0.n99 ));
    InMux I__8280 (
            .O(N__43303),
            .I(N__43300));
    LocalMux I__8279 (
            .O(N__43300),
            .I(N__43296));
    InMux I__8278 (
            .O(N__43299),
            .I(N__43293));
    Span4Mux_v I__8277 (
            .O(N__43296),
            .I(N__43290));
    LocalMux I__8276 (
            .O(N__43293),
            .I(N__43287));
    Odrv4 I__8275 (
            .O(N__43290),
            .I(\c0.n47_adj_3408 ));
    Odrv4 I__8274 (
            .O(N__43287),
            .I(\c0.n47_adj_3408 ));
    InMux I__8273 (
            .O(N__43282),
            .I(N__43279));
    LocalMux I__8272 (
            .O(N__43279),
            .I(N__43270));
    InMux I__8271 (
            .O(N__43278),
            .I(N__43267));
    InMux I__8270 (
            .O(N__43277),
            .I(N__43262));
    InMux I__8269 (
            .O(N__43276),
            .I(N__43262));
    InMux I__8268 (
            .O(N__43275),
            .I(N__43257));
    InMux I__8267 (
            .O(N__43274),
            .I(N__43257));
    InMux I__8266 (
            .O(N__43273),
            .I(N__43254));
    Span4Mux_v I__8265 (
            .O(N__43270),
            .I(N__43247));
    LocalMux I__8264 (
            .O(N__43267),
            .I(N__43247));
    LocalMux I__8263 (
            .O(N__43262),
            .I(N__43247));
    LocalMux I__8262 (
            .O(N__43257),
            .I(\c0.n18435 ));
    LocalMux I__8261 (
            .O(N__43254),
            .I(\c0.n18435 ));
    Odrv4 I__8260 (
            .O(N__43247),
            .I(\c0.n18435 ));
    CascadeMux I__8259 (
            .O(N__43240),
            .I(\c0.n42_adj_3064_cascade_ ));
    InMux I__8258 (
            .O(N__43237),
            .I(N__43234));
    LocalMux I__8257 (
            .O(N__43234),
            .I(N__43231));
    Span4Mux_v I__8256 (
            .O(N__43231),
            .I(N__43227));
    InMux I__8255 (
            .O(N__43230),
            .I(N__43224));
    Span4Mux_v I__8254 (
            .O(N__43227),
            .I(N__43221));
    LocalMux I__8253 (
            .O(N__43224),
            .I(N__43218));
    Odrv4 I__8252 (
            .O(N__43221),
            .I(\c0.n5_adj_3040 ));
    Odrv4 I__8251 (
            .O(N__43218),
            .I(\c0.n5_adj_3040 ));
    InMux I__8250 (
            .O(N__43213),
            .I(N__43210));
    LocalMux I__8249 (
            .O(N__43210),
            .I(N__43207));
    Span4Mux_v I__8248 (
            .O(N__43207),
            .I(N__43204));
    Span4Mux_v I__8247 (
            .O(N__43204),
            .I(N__43201));
    Odrv4 I__8246 (
            .O(N__43201),
            .I(\c0.n42_adj_3560 ));
    CascadeMux I__8245 (
            .O(N__43198),
            .I(\c0.n35_adj_3342_cascade_ ));
    InMux I__8244 (
            .O(N__43195),
            .I(N__43192));
    LocalMux I__8243 (
            .O(N__43192),
            .I(N__43189));
    Span4Mux_h I__8242 (
            .O(N__43189),
            .I(N__43186));
    Span4Mux_v I__8241 (
            .O(N__43186),
            .I(N__43183));
    Odrv4 I__8240 (
            .O(N__43183),
            .I(\c0.n39_adj_3339 ));
    InMux I__8239 (
            .O(N__43180),
            .I(N__43176));
    CascadeMux I__8238 (
            .O(N__43179),
            .I(N__43173));
    LocalMux I__8237 (
            .O(N__43176),
            .I(N__43170));
    InMux I__8236 (
            .O(N__43173),
            .I(N__43167));
    Span4Mux_v I__8235 (
            .O(N__43170),
            .I(N__43164));
    LocalMux I__8234 (
            .O(N__43167),
            .I(N__43161));
    Odrv4 I__8233 (
            .O(N__43164),
            .I(\c0.n12_adj_3015 ));
    Odrv4 I__8232 (
            .O(N__43161),
            .I(\c0.n12_adj_3015 ));
    CascadeMux I__8231 (
            .O(N__43156),
            .I(\c0.n44_adj_3561_cascade_ ));
    InMux I__8230 (
            .O(N__43153),
            .I(N__43150));
    LocalMux I__8229 (
            .O(N__43150),
            .I(N__43146));
    InMux I__8228 (
            .O(N__43149),
            .I(N__43143));
    Span4Mux_h I__8227 (
            .O(N__43146),
            .I(N__43140));
    LocalMux I__8226 (
            .O(N__43143),
            .I(N__43137));
    Span4Mux_v I__8225 (
            .O(N__43140),
            .I(N__43132));
    Span4Mux_h I__8224 (
            .O(N__43137),
            .I(N__43132));
    Span4Mux_h I__8223 (
            .O(N__43132),
            .I(N__43129));
    Odrv4 I__8222 (
            .O(N__43129),
            .I(\c0.n13_adj_3017 ));
    InMux I__8221 (
            .O(N__43126),
            .I(N__43123));
    LocalMux I__8220 (
            .O(N__43123),
            .I(\c0.n21118 ));
    InMux I__8219 (
            .O(N__43120),
            .I(N__43117));
    LocalMux I__8218 (
            .O(N__43117),
            .I(N__43113));
    InMux I__8217 (
            .O(N__43116),
            .I(N__43110));
    Span4Mux_h I__8216 (
            .O(N__43113),
            .I(N__43107));
    LocalMux I__8215 (
            .O(N__43110),
            .I(data_in_frame_18_2));
    Odrv4 I__8214 (
            .O(N__43107),
            .I(data_in_frame_18_2));
    CascadeMux I__8213 (
            .O(N__43102),
            .I(\c0.n21118_cascade_ ));
    InMux I__8212 (
            .O(N__43099),
            .I(N__43096));
    LocalMux I__8211 (
            .O(N__43096),
            .I(\c0.n13_adj_3139 ));
    InMux I__8210 (
            .O(N__43093),
            .I(N__43090));
    LocalMux I__8209 (
            .O(N__43090),
            .I(N__43084));
    InMux I__8208 (
            .O(N__43089),
            .I(N__43081));
    InMux I__8207 (
            .O(N__43088),
            .I(N__43078));
    InMux I__8206 (
            .O(N__43087),
            .I(N__43075));
    Sp12to4 I__8205 (
            .O(N__43084),
            .I(N__43070));
    LocalMux I__8204 (
            .O(N__43081),
            .I(N__43070));
    LocalMux I__8203 (
            .O(N__43078),
            .I(\c0.n36_adj_3267 ));
    LocalMux I__8202 (
            .O(N__43075),
            .I(\c0.n36_adj_3267 ));
    Odrv12 I__8201 (
            .O(N__43070),
            .I(\c0.n36_adj_3267 ));
    CascadeMux I__8200 (
            .O(N__43063),
            .I(\c0.n96_adj_3418_cascade_ ));
    InMux I__8199 (
            .O(N__43060),
            .I(N__43057));
    LocalMux I__8198 (
            .O(N__43057),
            .I(N__43054));
    Span4Mux_v I__8197 (
            .O(N__43054),
            .I(N__43051));
    Odrv4 I__8196 (
            .O(N__43051),
            .I(\c0.n99_adj_3424 ));
    InMux I__8195 (
            .O(N__43048),
            .I(N__43045));
    LocalMux I__8194 (
            .O(N__43045),
            .I(\c0.n77_adj_3415 ));
    CascadeMux I__8193 (
            .O(N__43042),
            .I(N__43038));
    CascadeMux I__8192 (
            .O(N__43041),
            .I(N__43035));
    InMux I__8191 (
            .O(N__43038),
            .I(N__43027));
    InMux I__8190 (
            .O(N__43035),
            .I(N__43027));
    InMux I__8189 (
            .O(N__43034),
            .I(N__43027));
    LocalMux I__8188 (
            .O(N__43027),
            .I(\c0.data_in_frame_10_2 ));
    InMux I__8187 (
            .O(N__43024),
            .I(N__43018));
    InMux I__8186 (
            .O(N__43023),
            .I(N__43018));
    LocalMux I__8185 (
            .O(N__43018),
            .I(N__43015));
    Odrv4 I__8184 (
            .O(N__43015),
            .I(\c0.n14_adj_3007 ));
    InMux I__8183 (
            .O(N__43012),
            .I(N__43009));
    LocalMux I__8182 (
            .O(N__43009),
            .I(N__43006));
    Span12Mux_v I__8181 (
            .O(N__43006),
            .I(N__43003));
    Odrv12 I__8180 (
            .O(N__43003),
            .I(\c0.n31_adj_3121 ));
    InMux I__8179 (
            .O(N__43000),
            .I(N__42997));
    LocalMux I__8178 (
            .O(N__42997),
            .I(N__42994));
    Odrv12 I__8177 (
            .O(N__42994),
            .I(\c0.n27 ));
    CascadeMux I__8176 (
            .O(N__42991),
            .I(\c0.n28_adj_3120_cascade_ ));
    InMux I__8175 (
            .O(N__42988),
            .I(N__42985));
    LocalMux I__8174 (
            .O(N__42985),
            .I(N__42982));
    Odrv4 I__8173 (
            .O(N__42982),
            .I(\c0.n33_adj_3122 ));
    CascadeMux I__8172 (
            .O(N__42979),
            .I(\c0.n20052_cascade_ ));
    CascadeMux I__8171 (
            .O(N__42976),
            .I(\c0.n10_adj_3129_cascade_ ));
    CascadeMux I__8170 (
            .O(N__42973),
            .I(\c0.n18400_cascade_ ));
    InMux I__8169 (
            .O(N__42970),
            .I(N__42965));
    InMux I__8168 (
            .O(N__42969),
            .I(N__42962));
    CascadeMux I__8167 (
            .O(N__42968),
            .I(N__42959));
    LocalMux I__8166 (
            .O(N__42965),
            .I(N__42956));
    LocalMux I__8165 (
            .O(N__42962),
            .I(N__42953));
    InMux I__8164 (
            .O(N__42959),
            .I(N__42950));
    Odrv4 I__8163 (
            .O(N__42956),
            .I(\c0.n20088 ));
    Odrv4 I__8162 (
            .O(N__42953),
            .I(\c0.n20088 ));
    LocalMux I__8161 (
            .O(N__42950),
            .I(\c0.n20088 ));
    CascadeMux I__8160 (
            .O(N__42943),
            .I(\c0.n20055_cascade_ ));
    CascadeMux I__8159 (
            .O(N__42940),
            .I(N__42937));
    InMux I__8158 (
            .O(N__42937),
            .I(N__42934));
    LocalMux I__8157 (
            .O(N__42934),
            .I(N__42930));
    InMux I__8156 (
            .O(N__42933),
            .I(N__42927));
    Span4Mux_h I__8155 (
            .O(N__42930),
            .I(N__42923));
    LocalMux I__8154 (
            .O(N__42927),
            .I(N__42920));
    InMux I__8153 (
            .O(N__42926),
            .I(N__42917));
    Span4Mux_v I__8152 (
            .O(N__42923),
            .I(N__42914));
    Sp12to4 I__8151 (
            .O(N__42920),
            .I(N__42909));
    LocalMux I__8150 (
            .O(N__42917),
            .I(N__42909));
    Odrv4 I__8149 (
            .O(N__42914),
            .I(\c0.n5_adj_3099 ));
    Odrv12 I__8148 (
            .O(N__42909),
            .I(\c0.n5_adj_3099 ));
    CascadeMux I__8147 (
            .O(N__42904),
            .I(\c0.n37_adj_3110_cascade_ ));
    InMux I__8146 (
            .O(N__42901),
            .I(N__42897));
    InMux I__8145 (
            .O(N__42900),
            .I(N__42894));
    LocalMux I__8144 (
            .O(N__42897),
            .I(\c0.n22_adj_3115 ));
    LocalMux I__8143 (
            .O(N__42894),
            .I(\c0.n22_adj_3115 ));
    CascadeMux I__8142 (
            .O(N__42889),
            .I(\c0.n6_adj_3024_cascade_ ));
    CascadeMux I__8141 (
            .O(N__42886),
            .I(\c0.n18435_cascade_ ));
    InMux I__8140 (
            .O(N__42883),
            .I(N__42880));
    LocalMux I__8139 (
            .O(N__42880),
            .I(\c0.n28_adj_3519 ));
    CascadeMux I__8138 (
            .O(N__42877),
            .I(\c0.n16_adj_3416_cascade_ ));
    InMux I__8137 (
            .O(N__42874),
            .I(N__42871));
    LocalMux I__8136 (
            .O(N__42871),
            .I(\c0.n16_adj_3542 ));
    CascadeMux I__8135 (
            .O(N__42868),
            .I(N__42865));
    InMux I__8134 (
            .O(N__42865),
            .I(N__42862));
    LocalMux I__8133 (
            .O(N__42862),
            .I(N__42858));
    InMux I__8132 (
            .O(N__42861),
            .I(N__42855));
    Odrv4 I__8131 (
            .O(N__42858),
            .I(\c0.n5_adj_3528 ));
    LocalMux I__8130 (
            .O(N__42855),
            .I(\c0.n5_adj_3528 ));
    CascadeMux I__8129 (
            .O(N__42850),
            .I(\c0.n78_cascade_ ));
    CascadeMux I__8128 (
            .O(N__42847),
            .I(\c0.n30_adj_3119_cascade_ ));
    CascadeMux I__8127 (
            .O(N__42844),
            .I(N__42841));
    InMux I__8126 (
            .O(N__42841),
            .I(N__42838));
    LocalMux I__8125 (
            .O(N__42838),
            .I(N__42835));
    Span4Mux_h I__8124 (
            .O(N__42835),
            .I(N__42832));
    Span4Mux_v I__8123 (
            .O(N__42832),
            .I(N__42829));
    Odrv4 I__8122 (
            .O(N__42829),
            .I(\c0.n6_adj_3453 ));
    CascadeMux I__8121 (
            .O(N__42826),
            .I(\c0.n39_adj_3398_cascade_ ));
    InMux I__8120 (
            .O(N__42823),
            .I(N__42820));
    LocalMux I__8119 (
            .O(N__42820),
            .I(\c0.n13_adj_3526 ));
    InMux I__8118 (
            .O(N__42817),
            .I(N__42813));
    InMux I__8117 (
            .O(N__42816),
            .I(N__42810));
    LocalMux I__8116 (
            .O(N__42813),
            .I(\c0.n14_adj_3525 ));
    LocalMux I__8115 (
            .O(N__42810),
            .I(\c0.n14_adj_3525 ));
    InMux I__8114 (
            .O(N__42805),
            .I(N__42802));
    LocalMux I__8113 (
            .O(N__42802),
            .I(\c0.n15_adj_3543 ));
    CascadeMux I__8112 (
            .O(N__42799),
            .I(\c0.n13_adj_3526_cascade_ ));
    CascadeMux I__8111 (
            .O(N__42796),
            .I(N__42793));
    InMux I__8110 (
            .O(N__42793),
            .I(N__42787));
    InMux I__8109 (
            .O(N__42792),
            .I(N__42787));
    LocalMux I__8108 (
            .O(N__42787),
            .I(\c0.n11_adj_3394 ));
    InMux I__8107 (
            .O(N__42784),
            .I(N__42780));
    InMux I__8106 (
            .O(N__42783),
            .I(N__42777));
    LocalMux I__8105 (
            .O(N__42780),
            .I(\c0.n11516 ));
    LocalMux I__8104 (
            .O(N__42777),
            .I(\c0.n11516 ));
    InMux I__8103 (
            .O(N__42772),
            .I(N__42769));
    LocalMux I__8102 (
            .O(N__42769),
            .I(\c0.n14_adj_3480 ));
    CascadeMux I__8101 (
            .O(N__42766),
            .I(\c0.n13_adj_3490_cascade_ ));
    InMux I__8100 (
            .O(N__42763),
            .I(N__42760));
    LocalMux I__8099 (
            .O(N__42760),
            .I(\c0.n13_adj_3546 ));
    InMux I__8098 (
            .O(N__42757),
            .I(N__42753));
    CascadeMux I__8097 (
            .O(N__42756),
            .I(N__42750));
    LocalMux I__8096 (
            .O(N__42753),
            .I(N__42747));
    InMux I__8095 (
            .O(N__42750),
            .I(N__42744));
    Span4Mux_h I__8094 (
            .O(N__42747),
            .I(N__42741));
    LocalMux I__8093 (
            .O(N__42744),
            .I(N__42738));
    Odrv4 I__8092 (
            .O(N__42741),
            .I(\c0.n15497 ));
    Odrv4 I__8091 (
            .O(N__42738),
            .I(\c0.n15497 ));
    InMux I__8090 (
            .O(N__42733),
            .I(N__42730));
    LocalMux I__8089 (
            .O(N__42730),
            .I(N__42727));
    Odrv4 I__8088 (
            .O(N__42727),
            .I(\c0.n14_adj_3459 ));
    InMux I__8087 (
            .O(N__42724),
            .I(N__42721));
    LocalMux I__8086 (
            .O(N__42721),
            .I(\c0.n10_adj_3068 ));
    CascadeMux I__8085 (
            .O(N__42718),
            .I(N__42714));
    InMux I__8084 (
            .O(N__42717),
            .I(N__42709));
    InMux I__8083 (
            .O(N__42714),
            .I(N__42709));
    LocalMux I__8082 (
            .O(N__42709),
            .I(N__42706));
    Odrv4 I__8081 (
            .O(N__42706),
            .I(\c0.n22_adj_3041 ));
    CascadeMux I__8080 (
            .O(N__42703),
            .I(N__42700));
    InMux I__8079 (
            .O(N__42700),
            .I(N__42697));
    LocalMux I__8078 (
            .O(N__42697),
            .I(N__42694));
    Odrv4 I__8077 (
            .O(N__42694),
            .I(\c0.n21079 ));
    InMux I__8076 (
            .O(N__42691),
            .I(N__42687));
    InMux I__8075 (
            .O(N__42690),
            .I(N__42684));
    LocalMux I__8074 (
            .O(N__42687),
            .I(N__42681));
    LocalMux I__8073 (
            .O(N__42684),
            .I(N__42676));
    Span4Mux_h I__8072 (
            .O(N__42681),
            .I(N__42676));
    Odrv4 I__8071 (
            .O(N__42676),
            .I(\c0.n26 ));
    InMux I__8070 (
            .O(N__42673),
            .I(N__42668));
    InMux I__8069 (
            .O(N__42672),
            .I(N__42665));
    InMux I__8068 (
            .O(N__42671),
            .I(N__42662));
    LocalMux I__8067 (
            .O(N__42668),
            .I(N__42659));
    LocalMux I__8066 (
            .O(N__42665),
            .I(N__42654));
    LocalMux I__8065 (
            .O(N__42662),
            .I(N__42654));
    Odrv4 I__8064 (
            .O(N__42659),
            .I(\c0.n5_adj_3044 ));
    Odrv12 I__8063 (
            .O(N__42654),
            .I(\c0.n5_adj_3044 ));
    InMux I__8062 (
            .O(N__42649),
            .I(N__42646));
    LocalMux I__8061 (
            .O(N__42646),
            .I(\c0.n25_adj_3045 ));
    CascadeMux I__8060 (
            .O(N__42643),
            .I(\c0.n14_adj_3073_cascade_ ));
    InMux I__8059 (
            .O(N__42640),
            .I(N__42637));
    LocalMux I__8058 (
            .O(N__42637),
            .I(N__42633));
    CascadeMux I__8057 (
            .O(N__42636),
            .I(N__42629));
    Span4Mux_v I__8056 (
            .O(N__42633),
            .I(N__42625));
    InMux I__8055 (
            .O(N__42632),
            .I(N__42622));
    InMux I__8054 (
            .O(N__42629),
            .I(N__42619));
    InMux I__8053 (
            .O(N__42628),
            .I(N__42616));
    Odrv4 I__8052 (
            .O(N__42625),
            .I(data_in_2_0));
    LocalMux I__8051 (
            .O(N__42622),
            .I(data_in_2_0));
    LocalMux I__8050 (
            .O(N__42619),
            .I(data_in_2_0));
    LocalMux I__8049 (
            .O(N__42616),
            .I(data_in_2_0));
    InMux I__8048 (
            .O(N__42607),
            .I(N__42599));
    InMux I__8047 (
            .O(N__42606),
            .I(N__42599));
    InMux I__8046 (
            .O(N__42605),
            .I(N__42594));
    InMux I__8045 (
            .O(N__42604),
            .I(N__42594));
    LocalMux I__8044 (
            .O(N__42599),
            .I(data_in_1_0));
    LocalMux I__8043 (
            .O(N__42594),
            .I(data_in_1_0));
    InMux I__8042 (
            .O(N__42589),
            .I(N__42586));
    LocalMux I__8041 (
            .O(N__42586),
            .I(N__42583));
    Span4Mux_v I__8040 (
            .O(N__42583),
            .I(N__42580));
    Odrv4 I__8039 (
            .O(N__42580),
            .I(\c0.n12_adj_3230 ));
    InMux I__8038 (
            .O(N__42577),
            .I(N__42571));
    InMux I__8037 (
            .O(N__42576),
            .I(N__42568));
    InMux I__8036 (
            .O(N__42575),
            .I(N__42565));
    InMux I__8035 (
            .O(N__42574),
            .I(N__42562));
    LocalMux I__8034 (
            .O(N__42571),
            .I(N__42555));
    LocalMux I__8033 (
            .O(N__42568),
            .I(N__42555));
    LocalMux I__8032 (
            .O(N__42565),
            .I(N__42555));
    LocalMux I__8031 (
            .O(N__42562),
            .I(data_in_2_7));
    Odrv12 I__8030 (
            .O(N__42555),
            .I(data_in_2_7));
    InMux I__8029 (
            .O(N__42550),
            .I(N__42547));
    LocalMux I__8028 (
            .O(N__42547),
            .I(\c0.n11443 ));
    InMux I__8027 (
            .O(N__42544),
            .I(N__42541));
    LocalMux I__8026 (
            .O(N__42541),
            .I(N__42537));
    InMux I__8025 (
            .O(N__42540),
            .I(N__42533));
    Span4Mux_h I__8024 (
            .O(N__42537),
            .I(N__42530));
    InMux I__8023 (
            .O(N__42536),
            .I(N__42527));
    LocalMux I__8022 (
            .O(N__42533),
            .I(data_in_0_1));
    Odrv4 I__8021 (
            .O(N__42530),
            .I(data_in_0_1));
    LocalMux I__8020 (
            .O(N__42527),
            .I(data_in_0_1));
    CascadeMux I__8019 (
            .O(N__42520),
            .I(N__42513));
    CascadeMux I__8018 (
            .O(N__42519),
            .I(N__42509));
    InMux I__8017 (
            .O(N__42518),
            .I(N__42501));
    InMux I__8016 (
            .O(N__42517),
            .I(N__42498));
    InMux I__8015 (
            .O(N__42516),
            .I(N__42488));
    InMux I__8014 (
            .O(N__42513),
            .I(N__42488));
    InMux I__8013 (
            .O(N__42512),
            .I(N__42488));
    InMux I__8012 (
            .O(N__42509),
            .I(N__42483));
    InMux I__8011 (
            .O(N__42508),
            .I(N__42483));
    CascadeMux I__8010 (
            .O(N__42507),
            .I(N__42480));
    InMux I__8009 (
            .O(N__42506),
            .I(N__42476));
    InMux I__8008 (
            .O(N__42505),
            .I(N__42473));
    InMux I__8007 (
            .O(N__42504),
            .I(N__42470));
    LocalMux I__8006 (
            .O(N__42501),
            .I(N__42467));
    LocalMux I__8005 (
            .O(N__42498),
            .I(N__42464));
    CascadeMux I__8004 (
            .O(N__42497),
            .I(N__42461));
    CascadeMux I__8003 (
            .O(N__42496),
            .I(N__42456));
    CascadeMux I__8002 (
            .O(N__42495),
            .I(N__42453));
    LocalMux I__8001 (
            .O(N__42488),
            .I(N__42448));
    LocalMux I__8000 (
            .O(N__42483),
            .I(N__42448));
    InMux I__7999 (
            .O(N__42480),
            .I(N__42443));
    InMux I__7998 (
            .O(N__42479),
            .I(N__42443));
    LocalMux I__7997 (
            .O(N__42476),
            .I(N__42438));
    LocalMux I__7996 (
            .O(N__42473),
            .I(N__42438));
    LocalMux I__7995 (
            .O(N__42470),
            .I(N__42435));
    Span4Mux_h I__7994 (
            .O(N__42467),
            .I(N__42430));
    Span4Mux_h I__7993 (
            .O(N__42464),
            .I(N__42430));
    InMux I__7992 (
            .O(N__42461),
            .I(N__42423));
    InMux I__7991 (
            .O(N__42460),
            .I(N__42418));
    InMux I__7990 (
            .O(N__42459),
            .I(N__42418));
    InMux I__7989 (
            .O(N__42456),
            .I(N__42415));
    InMux I__7988 (
            .O(N__42453),
            .I(N__42412));
    Span4Mux_v I__7987 (
            .O(N__42448),
            .I(N__42403));
    LocalMux I__7986 (
            .O(N__42443),
            .I(N__42403));
    Span4Mux_v I__7985 (
            .O(N__42438),
            .I(N__42403));
    Span4Mux_h I__7984 (
            .O(N__42435),
            .I(N__42403));
    Span4Mux_v I__7983 (
            .O(N__42430),
            .I(N__42400));
    InMux I__7982 (
            .O(N__42429),
            .I(N__42393));
    InMux I__7981 (
            .O(N__42428),
            .I(N__42393));
    InMux I__7980 (
            .O(N__42427),
            .I(N__42393));
    InMux I__7979 (
            .O(N__42426),
            .I(N__42390));
    LocalMux I__7978 (
            .O(N__42423),
            .I(N__42385));
    LocalMux I__7977 (
            .O(N__42418),
            .I(N__42385));
    LocalMux I__7976 (
            .O(N__42415),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7975 (
            .O(N__42412),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__7974 (
            .O(N__42403),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__7973 (
            .O(N__42400),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7972 (
            .O(N__42393),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7971 (
            .O(N__42390),
            .I(FRAME_MATCHER_state_1));
    Odrv12 I__7970 (
            .O(N__42385),
            .I(FRAME_MATCHER_state_1));
    InMux I__7969 (
            .O(N__42370),
            .I(N__42365));
    InMux I__7968 (
            .O(N__42369),
            .I(N__42361));
    InMux I__7967 (
            .O(N__42368),
            .I(N__42358));
    LocalMux I__7966 (
            .O(N__42365),
            .I(N__42355));
    InMux I__7965 (
            .O(N__42364),
            .I(N__42352));
    LocalMux I__7964 (
            .O(N__42361),
            .I(N__42349));
    LocalMux I__7963 (
            .O(N__42358),
            .I(N__42346));
    Span4Mux_v I__7962 (
            .O(N__42355),
            .I(N__42343));
    LocalMux I__7961 (
            .O(N__42352),
            .I(N__42338));
    Span4Mux_h I__7960 (
            .O(N__42349),
            .I(N__42338));
    Odrv12 I__7959 (
            .O(N__42346),
            .I(n4_adj_3596));
    Odrv4 I__7958 (
            .O(N__42343),
            .I(n4_adj_3596));
    Odrv4 I__7957 (
            .O(N__42338),
            .I(n4_adj_3596));
    InMux I__7956 (
            .O(N__42331),
            .I(N__42325));
    InMux I__7955 (
            .O(N__42330),
            .I(N__42320));
    InMux I__7954 (
            .O(N__42329),
            .I(N__42317));
    InMux I__7953 (
            .O(N__42328),
            .I(N__42314));
    LocalMux I__7952 (
            .O(N__42325),
            .I(N__42311));
    InMux I__7951 (
            .O(N__42324),
            .I(N__42305));
    InMux I__7950 (
            .O(N__42323),
            .I(N__42305));
    LocalMux I__7949 (
            .O(N__42320),
            .I(N__42302));
    LocalMux I__7948 (
            .O(N__42317),
            .I(N__42299));
    LocalMux I__7947 (
            .O(N__42314),
            .I(N__42294));
    Span4Mux_h I__7946 (
            .O(N__42311),
            .I(N__42294));
    InMux I__7945 (
            .O(N__42310),
            .I(N__42290));
    LocalMux I__7944 (
            .O(N__42305),
            .I(N__42287));
    Span4Mux_h I__7943 (
            .O(N__42302),
            .I(N__42280));
    Span4Mux_h I__7942 (
            .O(N__42299),
            .I(N__42280));
    Span4Mux_v I__7941 (
            .O(N__42294),
            .I(N__42280));
    InMux I__7940 (
            .O(N__42293),
            .I(N__42277));
    LocalMux I__7939 (
            .O(N__42290),
            .I(n11421));
    Odrv12 I__7938 (
            .O(N__42287),
            .I(n11421));
    Odrv4 I__7937 (
            .O(N__42280),
            .I(n11421));
    LocalMux I__7936 (
            .O(N__42277),
            .I(n11421));
    InMux I__7935 (
            .O(N__42268),
            .I(N__42262));
    InMux I__7934 (
            .O(N__42267),
            .I(N__42259));
    InMux I__7933 (
            .O(N__42266),
            .I(N__42256));
    InMux I__7932 (
            .O(N__42265),
            .I(N__42253));
    LocalMux I__7931 (
            .O(N__42262),
            .I(N__42240));
    LocalMux I__7930 (
            .O(N__42259),
            .I(N__42240));
    LocalMux I__7929 (
            .O(N__42256),
            .I(N__42240));
    LocalMux I__7928 (
            .O(N__42253),
            .I(N__42240));
    InMux I__7927 (
            .O(N__42252),
            .I(N__42237));
    InMux I__7926 (
            .O(N__42251),
            .I(N__42234));
    InMux I__7925 (
            .O(N__42250),
            .I(N__42231));
    InMux I__7924 (
            .O(N__42249),
            .I(N__42228));
    Span4Mux_v I__7923 (
            .O(N__42240),
            .I(N__42213));
    LocalMux I__7922 (
            .O(N__42237),
            .I(N__42213));
    LocalMux I__7921 (
            .O(N__42234),
            .I(N__42213));
    LocalMux I__7920 (
            .O(N__42231),
            .I(N__42213));
    LocalMux I__7919 (
            .O(N__42228),
            .I(N__42213));
    InMux I__7918 (
            .O(N__42227),
            .I(N__42210));
    InMux I__7917 (
            .O(N__42226),
            .I(N__42207));
    InMux I__7916 (
            .O(N__42225),
            .I(N__42204));
    InMux I__7915 (
            .O(N__42224),
            .I(N__42201));
    Span4Mux_v I__7914 (
            .O(N__42213),
            .I(N__42184));
    LocalMux I__7913 (
            .O(N__42210),
            .I(N__42184));
    LocalMux I__7912 (
            .O(N__42207),
            .I(N__42184));
    LocalMux I__7911 (
            .O(N__42204),
            .I(N__42184));
    LocalMux I__7910 (
            .O(N__42201),
            .I(N__42184));
    InMux I__7909 (
            .O(N__42200),
            .I(N__42181));
    InMux I__7908 (
            .O(N__42199),
            .I(N__42178));
    InMux I__7907 (
            .O(N__42198),
            .I(N__42175));
    InMux I__7906 (
            .O(N__42197),
            .I(N__42172));
    InMux I__7905 (
            .O(N__42196),
            .I(N__42164));
    InMux I__7904 (
            .O(N__42195),
            .I(N__42164));
    Span4Mux_v I__7903 (
            .O(N__42184),
            .I(N__42153));
    LocalMux I__7902 (
            .O(N__42181),
            .I(N__42153));
    LocalMux I__7901 (
            .O(N__42178),
            .I(N__42153));
    LocalMux I__7900 (
            .O(N__42175),
            .I(N__42153));
    LocalMux I__7899 (
            .O(N__42172),
            .I(N__42153));
    InMux I__7898 (
            .O(N__42171),
            .I(N__42146));
    InMux I__7897 (
            .O(N__42170),
            .I(N__42146));
    InMux I__7896 (
            .O(N__42169),
            .I(N__42146));
    LocalMux I__7895 (
            .O(N__42164),
            .I(N__42133));
    Span4Mux_v I__7894 (
            .O(N__42153),
            .I(N__42133));
    LocalMux I__7893 (
            .O(N__42146),
            .I(N__42133));
    InMux I__7892 (
            .O(N__42145),
            .I(N__42128));
    InMux I__7891 (
            .O(N__42144),
            .I(N__42122));
    InMux I__7890 (
            .O(N__42143),
            .I(N__42118));
    InMux I__7889 (
            .O(N__42142),
            .I(N__42115));
    InMux I__7888 (
            .O(N__42141),
            .I(N__42112));
    InMux I__7887 (
            .O(N__42140),
            .I(N__42109));
    Span4Mux_h I__7886 (
            .O(N__42133),
            .I(N__42106));
    InMux I__7885 (
            .O(N__42132),
            .I(N__42103));
    InMux I__7884 (
            .O(N__42131),
            .I(N__42100));
    LocalMux I__7883 (
            .O(N__42128),
            .I(N__42097));
    InMux I__7882 (
            .O(N__42127),
            .I(N__42094));
    InMux I__7881 (
            .O(N__42126),
            .I(N__42091));
    InMux I__7880 (
            .O(N__42125),
            .I(N__42088));
    LocalMux I__7879 (
            .O(N__42122),
            .I(N__42085));
    InMux I__7878 (
            .O(N__42121),
            .I(N__42082));
    LocalMux I__7877 (
            .O(N__42118),
            .I(N__42075));
    LocalMux I__7876 (
            .O(N__42115),
            .I(N__42075));
    LocalMux I__7875 (
            .O(N__42112),
            .I(N__42075));
    LocalMux I__7874 (
            .O(N__42109),
            .I(N__42072));
    Sp12to4 I__7873 (
            .O(N__42106),
            .I(N__42068));
    LocalMux I__7872 (
            .O(N__42103),
            .I(N__42065));
    LocalMux I__7871 (
            .O(N__42100),
            .I(N__42062));
    Span4Mux_h I__7870 (
            .O(N__42097),
            .I(N__42057));
    LocalMux I__7869 (
            .O(N__42094),
            .I(N__42057));
    LocalMux I__7868 (
            .O(N__42091),
            .I(N__42048));
    LocalMux I__7867 (
            .O(N__42088),
            .I(N__42048));
    Span4Mux_s1_v I__7866 (
            .O(N__42085),
            .I(N__42048));
    LocalMux I__7865 (
            .O(N__42082),
            .I(N__42048));
    Span4Mux_v I__7864 (
            .O(N__42075),
            .I(N__42043));
    Span4Mux_v I__7863 (
            .O(N__42072),
            .I(N__42043));
    InMux I__7862 (
            .O(N__42071),
            .I(N__42040));
    Span12Mux_s7_v I__7861 (
            .O(N__42068),
            .I(N__42037));
    Span12Mux_h I__7860 (
            .O(N__42065),
            .I(N__42034));
    Span4Mux_h I__7859 (
            .O(N__42062),
            .I(N__42031));
    Span4Mux_v I__7858 (
            .O(N__42057),
            .I(N__42026));
    Span4Mux_v I__7857 (
            .O(N__42048),
            .I(N__42026));
    Span4Mux_h I__7856 (
            .O(N__42043),
            .I(N__42021));
    LocalMux I__7855 (
            .O(N__42040),
            .I(N__42021));
    Span12Mux_v I__7854 (
            .O(N__42037),
            .I(N__42018));
    Span12Mux_v I__7853 (
            .O(N__42034),
            .I(N__42015));
    Odrv4 I__7852 (
            .O(N__42031),
            .I(n1295));
    Odrv4 I__7851 (
            .O(N__42026),
            .I(n1295));
    Odrv4 I__7850 (
            .O(N__42021),
            .I(n1295));
    Odrv12 I__7849 (
            .O(N__42018),
            .I(n1295));
    Odrv12 I__7848 (
            .O(N__42015),
            .I(n1295));
    CascadeMux I__7847 (
            .O(N__42004),
            .I(N__41999));
    InMux I__7846 (
            .O(N__42003),
            .I(N__41995));
    InMux I__7845 (
            .O(N__42002),
            .I(N__41992));
    InMux I__7844 (
            .O(N__41999),
            .I(N__41987));
    InMux I__7843 (
            .O(N__41998),
            .I(N__41987));
    LocalMux I__7842 (
            .O(N__41995),
            .I(N__41982));
    LocalMux I__7841 (
            .O(N__41992),
            .I(N__41982));
    LocalMux I__7840 (
            .O(N__41987),
            .I(\c0.data_in_frame_27_7 ));
    Odrv12 I__7839 (
            .O(N__41982),
            .I(\c0.data_in_frame_27_7 ));
    InMux I__7838 (
            .O(N__41977),
            .I(N__41974));
    LocalMux I__7837 (
            .O(N__41974),
            .I(N__41968));
    InMux I__7836 (
            .O(N__41973),
            .I(N__41965));
    InMux I__7835 (
            .O(N__41972),
            .I(N__41960));
    InMux I__7834 (
            .O(N__41971),
            .I(N__41960));
    Sp12to4 I__7833 (
            .O(N__41968),
            .I(N__41955));
    LocalMux I__7832 (
            .O(N__41965),
            .I(N__41955));
    LocalMux I__7831 (
            .O(N__41960),
            .I(\c0.data_in_frame_27_6 ));
    Odrv12 I__7830 (
            .O(N__41955),
            .I(\c0.data_in_frame_27_6 ));
    CascadeMux I__7829 (
            .O(N__41950),
            .I(N__41946));
    CascadeMux I__7828 (
            .O(N__41949),
            .I(N__41943));
    InMux I__7827 (
            .O(N__41946),
            .I(N__41939));
    InMux I__7826 (
            .O(N__41943),
            .I(N__41934));
    InMux I__7825 (
            .O(N__41942),
            .I(N__41934));
    LocalMux I__7824 (
            .O(N__41939),
            .I(\c0.data_in_frame_26_4 ));
    LocalMux I__7823 (
            .O(N__41934),
            .I(\c0.data_in_frame_26_4 ));
    InMux I__7822 (
            .O(N__41929),
            .I(N__41923));
    InMux I__7821 (
            .O(N__41928),
            .I(N__41918));
    InMux I__7820 (
            .O(N__41927),
            .I(N__41918));
    InMux I__7819 (
            .O(N__41926),
            .I(N__41915));
    LocalMux I__7818 (
            .O(N__41923),
            .I(data_in_2_2));
    LocalMux I__7817 (
            .O(N__41918),
            .I(data_in_2_2));
    LocalMux I__7816 (
            .O(N__41915),
            .I(data_in_2_2));
    InMux I__7815 (
            .O(N__41908),
            .I(N__41905));
    LocalMux I__7814 (
            .O(N__41905),
            .I(\c0.n10_adj_3238 ));
    InMux I__7813 (
            .O(N__41902),
            .I(N__41899));
    LocalMux I__7812 (
            .O(N__41899),
            .I(N__41896));
    Span4Mux_v I__7811 (
            .O(N__41896),
            .I(N__41892));
    InMux I__7810 (
            .O(N__41895),
            .I(N__41889));
    Odrv4 I__7809 (
            .O(N__41892),
            .I(\c0.n110 ));
    LocalMux I__7808 (
            .O(N__41889),
            .I(\c0.n110 ));
    InMux I__7807 (
            .O(N__41884),
            .I(N__41881));
    LocalMux I__7806 (
            .O(N__41881),
            .I(N__41878));
    Span4Mux_v I__7805 (
            .O(N__41878),
            .I(N__41872));
    InMux I__7804 (
            .O(N__41877),
            .I(N__41869));
    InMux I__7803 (
            .O(N__41876),
            .I(N__41866));
    InMux I__7802 (
            .O(N__41875),
            .I(N__41863));
    Odrv4 I__7801 (
            .O(N__41872),
            .I(data_in_2_5));
    LocalMux I__7800 (
            .O(N__41869),
            .I(data_in_2_5));
    LocalMux I__7799 (
            .O(N__41866),
            .I(data_in_2_5));
    LocalMux I__7798 (
            .O(N__41863),
            .I(data_in_2_5));
    InMux I__7797 (
            .O(N__41854),
            .I(N__41848));
    InMux I__7796 (
            .O(N__41853),
            .I(N__41845));
    InMux I__7795 (
            .O(N__41852),
            .I(N__41840));
    InMux I__7794 (
            .O(N__41851),
            .I(N__41840));
    LocalMux I__7793 (
            .O(N__41848),
            .I(data_in_1_5));
    LocalMux I__7792 (
            .O(N__41845),
            .I(data_in_1_5));
    LocalMux I__7791 (
            .O(N__41840),
            .I(data_in_1_5));
    InMux I__7790 (
            .O(N__41833),
            .I(N__41830));
    LocalMux I__7789 (
            .O(N__41830),
            .I(N__41826));
    CascadeMux I__7788 (
            .O(N__41829),
            .I(N__41823));
    Span12Mux_s9_v I__7787 (
            .O(N__41826),
            .I(N__41820));
    InMux I__7786 (
            .O(N__41823),
            .I(N__41817));
    Span12Mux_h I__7785 (
            .O(N__41820),
            .I(N__41814));
    LocalMux I__7784 (
            .O(N__41817),
            .I(N__41811));
    Span12Mux_v I__7783 (
            .O(N__41814),
            .I(N__41808));
    Span4Mux_v I__7782 (
            .O(N__41811),
            .I(N__41805));
    Odrv12 I__7781 (
            .O(N__41808),
            .I(\c0.n160 ));
    Odrv4 I__7780 (
            .O(N__41805),
            .I(\c0.n160 ));
    InMux I__7779 (
            .O(N__41800),
            .I(N__41794));
    InMux I__7778 (
            .O(N__41799),
            .I(N__41794));
    LocalMux I__7777 (
            .O(N__41794),
            .I(\c0.data_in_frame_29_0 ));
    CascadeMux I__7776 (
            .O(N__41791),
            .I(\c0.n21117_cascade_ ));
    InMux I__7775 (
            .O(N__41788),
            .I(N__41785));
    LocalMux I__7774 (
            .O(N__41785),
            .I(\c0.n18 ));
    InMux I__7773 (
            .O(N__41782),
            .I(N__41779));
    LocalMux I__7772 (
            .O(N__41779),
            .I(\c0.n5_adj_3142 ));
    CascadeMux I__7771 (
            .O(N__41776),
            .I(\c0.n5_adj_3142_cascade_ ));
    CascadeMux I__7770 (
            .O(N__41773),
            .I(\c0.n22_adj_3305_cascade_ ));
    CascadeMux I__7769 (
            .O(N__41770),
            .I(\c0.n37_adj_3309_cascade_ ));
    CascadeMux I__7768 (
            .O(N__41767),
            .I(\c0.n21099_cascade_ ));
    InMux I__7767 (
            .O(N__41764),
            .I(N__41761));
    LocalMux I__7766 (
            .O(N__41761),
            .I(\c0.n18_adj_3314 ));
    CascadeMux I__7765 (
            .O(N__41758),
            .I(\c0.n10_adj_3353_cascade_ ));
    InMux I__7764 (
            .O(N__41755),
            .I(N__41752));
    LocalMux I__7763 (
            .O(N__41752),
            .I(N__41749));
    Span12Mux_v I__7762 (
            .O(N__41749),
            .I(N__41746));
    Odrv12 I__7761 (
            .O(N__41746),
            .I(\c0.n21111 ));
    CascadeMux I__7760 (
            .O(N__41743),
            .I(\c0.n9_adj_3352_cascade_ ));
    InMux I__7759 (
            .O(N__41740),
            .I(N__41737));
    LocalMux I__7758 (
            .O(N__41737),
            .I(\c0.n21051 ));
    InMux I__7757 (
            .O(N__41734),
            .I(N__41731));
    LocalMux I__7756 (
            .O(N__41731),
            .I(N__41728));
    Span4Mux_v I__7755 (
            .O(N__41728),
            .I(N__41725));
    Odrv4 I__7754 (
            .O(N__41725),
            .I(\c0.n18537 ));
    InMux I__7753 (
            .O(N__41722),
            .I(N__41718));
    InMux I__7752 (
            .O(N__41721),
            .I(N__41715));
    LocalMux I__7751 (
            .O(N__41718),
            .I(\c0.n20370 ));
    LocalMux I__7750 (
            .O(N__41715),
            .I(\c0.n20370 ));
    CascadeMux I__7749 (
            .O(N__41710),
            .I(N__41707));
    InMux I__7748 (
            .O(N__41707),
            .I(N__41703));
    InMux I__7747 (
            .O(N__41706),
            .I(N__41700));
    LocalMux I__7746 (
            .O(N__41703),
            .I(\c0.data_in_frame_29_7 ));
    LocalMux I__7745 (
            .O(N__41700),
            .I(\c0.data_in_frame_29_7 ));
    CascadeMux I__7744 (
            .O(N__41695),
            .I(N__41691));
    CascadeMux I__7743 (
            .O(N__41694),
            .I(N__41688));
    InMux I__7742 (
            .O(N__41691),
            .I(N__41685));
    InMux I__7741 (
            .O(N__41688),
            .I(N__41682));
    LocalMux I__7740 (
            .O(N__41685),
            .I(\c0.data_in_frame_29_6 ));
    LocalMux I__7739 (
            .O(N__41682),
            .I(\c0.data_in_frame_29_6 ));
    CascadeMux I__7738 (
            .O(N__41677),
            .I(\c0.n10_adj_3152_cascade_ ));
    InMux I__7737 (
            .O(N__41674),
            .I(N__41671));
    LocalMux I__7736 (
            .O(N__41671),
            .I(\c0.n21117 ));
    CascadeMux I__7735 (
            .O(N__41668),
            .I(\c0.n61_cascade_ ));
    InMux I__7734 (
            .O(N__41665),
            .I(N__41662));
    LocalMux I__7733 (
            .O(N__41662),
            .I(\c0.n50 ));
    InMux I__7732 (
            .O(N__41659),
            .I(N__41656));
    LocalMux I__7731 (
            .O(N__41656),
            .I(\c0.n61 ));
    CascadeMux I__7730 (
            .O(N__41653),
            .I(\c0.n86_adj_3393_cascade_ ));
    CascadeMux I__7729 (
            .O(N__41650),
            .I(\c0.n95_cascade_ ));
    InMux I__7728 (
            .O(N__41647),
            .I(N__41644));
    LocalMux I__7727 (
            .O(N__41644),
            .I(N__41641));
    Span4Mux_v I__7726 (
            .O(N__41641),
            .I(N__41638));
    Odrv4 I__7725 (
            .O(N__41638),
            .I(\c0.n15_adj_3441 ));
    InMux I__7724 (
            .O(N__41635),
            .I(N__41632));
    LocalMux I__7723 (
            .O(N__41632),
            .I(N__41628));
    InMux I__7722 (
            .O(N__41631),
            .I(N__41625));
    Span4Mux_v I__7721 (
            .O(N__41628),
            .I(N__41620));
    LocalMux I__7720 (
            .O(N__41625),
            .I(N__41617));
    InMux I__7719 (
            .O(N__41624),
            .I(N__41612));
    InMux I__7718 (
            .O(N__41623),
            .I(N__41612));
    Odrv4 I__7717 (
            .O(N__41620),
            .I(data_in_3_7));
    Odrv4 I__7716 (
            .O(N__41617),
            .I(data_in_3_7));
    LocalMux I__7715 (
            .O(N__41612),
            .I(data_in_3_7));
    CascadeMux I__7714 (
            .O(N__41605),
            .I(N__41601));
    CascadeMux I__7713 (
            .O(N__41604),
            .I(N__41597));
    InMux I__7712 (
            .O(N__41601),
            .I(N__41594));
    InMux I__7711 (
            .O(N__41600),
            .I(N__41591));
    InMux I__7710 (
            .O(N__41597),
            .I(N__41588));
    LocalMux I__7709 (
            .O(N__41594),
            .I(N__41585));
    LocalMux I__7708 (
            .O(N__41591),
            .I(data_in_frame_16_6));
    LocalMux I__7707 (
            .O(N__41588),
            .I(data_in_frame_16_6));
    Odrv12 I__7706 (
            .O(N__41585),
            .I(data_in_frame_16_6));
    InMux I__7705 (
            .O(N__41578),
            .I(N__41574));
    InMux I__7704 (
            .O(N__41577),
            .I(N__41571));
    LocalMux I__7703 (
            .O(N__41574),
            .I(\c0.data_in_frame_28_4 ));
    LocalMux I__7702 (
            .O(N__41571),
            .I(\c0.data_in_frame_28_4 ));
    InMux I__7701 (
            .O(N__41566),
            .I(N__41563));
    LocalMux I__7700 (
            .O(N__41563),
            .I(N__41560));
    Span4Mux_h I__7699 (
            .O(N__41560),
            .I(N__41557));
    Span4Mux_v I__7698 (
            .O(N__41557),
            .I(N__41554));
    Odrv4 I__7697 (
            .O(N__41554),
            .I(\c0.n20931 ));
    InMux I__7696 (
            .O(N__41551),
            .I(N__41548));
    LocalMux I__7695 (
            .O(N__41548),
            .I(N__41544));
    InMux I__7694 (
            .O(N__41547),
            .I(N__41541));
    Span4Mux_v I__7693 (
            .O(N__41544),
            .I(N__41538));
    LocalMux I__7692 (
            .O(N__41541),
            .I(data_in_frame_18_6));
    Odrv4 I__7691 (
            .O(N__41538),
            .I(data_in_frame_18_6));
    InMux I__7690 (
            .O(N__41533),
            .I(N__41530));
    LocalMux I__7689 (
            .O(N__41530),
            .I(N__41526));
    InMux I__7688 (
            .O(N__41529),
            .I(N__41523));
    Odrv4 I__7687 (
            .O(N__41526),
            .I(n4_adj_3595));
    LocalMux I__7686 (
            .O(N__41523),
            .I(n4_adj_3595));
    InMux I__7685 (
            .O(N__41518),
            .I(N__41515));
    LocalMux I__7684 (
            .O(N__41515),
            .I(N__41512));
    Span4Mux_v I__7683 (
            .O(N__41512),
            .I(N__41509));
    Odrv4 I__7682 (
            .O(N__41509),
            .I(\c0.n14_adj_3434 ));
    InMux I__7681 (
            .O(N__41506),
            .I(N__41500));
    InMux I__7680 (
            .O(N__41505),
            .I(N__41500));
    LocalMux I__7679 (
            .O(N__41500),
            .I(N__41497));
    Span4Mux_v I__7678 (
            .O(N__41497),
            .I(N__41492));
    InMux I__7677 (
            .O(N__41496),
            .I(N__41489));
    InMux I__7676 (
            .O(N__41495),
            .I(N__41486));
    Span4Mux_h I__7675 (
            .O(N__41492),
            .I(N__41483));
    LocalMux I__7674 (
            .O(N__41489),
            .I(\c0.FRAME_MATCHER_state_12 ));
    LocalMux I__7673 (
            .O(N__41486),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv4 I__7672 (
            .O(N__41483),
            .I(\c0.FRAME_MATCHER_state_12 ));
    InMux I__7671 (
            .O(N__41476),
            .I(N__41473));
    LocalMux I__7670 (
            .O(N__41473),
            .I(N__41453));
    InMux I__7669 (
            .O(N__41472),
            .I(N__41450));
    InMux I__7668 (
            .O(N__41471),
            .I(N__41444));
    InMux I__7667 (
            .O(N__41470),
            .I(N__41444));
    InMux I__7666 (
            .O(N__41469),
            .I(N__41441));
    InMux I__7665 (
            .O(N__41468),
            .I(N__41436));
    InMux I__7664 (
            .O(N__41467),
            .I(N__41436));
    InMux I__7663 (
            .O(N__41466),
            .I(N__41430));
    InMux I__7662 (
            .O(N__41465),
            .I(N__41423));
    InMux I__7661 (
            .O(N__41464),
            .I(N__41423));
    InMux I__7660 (
            .O(N__41463),
            .I(N__41414));
    InMux I__7659 (
            .O(N__41462),
            .I(N__41414));
    InMux I__7658 (
            .O(N__41461),
            .I(N__41414));
    InMux I__7657 (
            .O(N__41460),
            .I(N__41414));
    InMux I__7656 (
            .O(N__41459),
            .I(N__41405));
    InMux I__7655 (
            .O(N__41458),
            .I(N__41405));
    InMux I__7654 (
            .O(N__41457),
            .I(N__41405));
    InMux I__7653 (
            .O(N__41456),
            .I(N__41405));
    Span4Mux_v I__7652 (
            .O(N__41453),
            .I(N__41400));
    LocalMux I__7651 (
            .O(N__41450),
            .I(N__41397));
    InMux I__7650 (
            .O(N__41449),
            .I(N__41394));
    LocalMux I__7649 (
            .O(N__41444),
            .I(N__41390));
    LocalMux I__7648 (
            .O(N__41441),
            .I(N__41387));
    LocalMux I__7647 (
            .O(N__41436),
            .I(N__41384));
    InMux I__7646 (
            .O(N__41435),
            .I(N__41381));
    InMux I__7645 (
            .O(N__41434),
            .I(N__41378));
    InMux I__7644 (
            .O(N__41433),
            .I(N__41375));
    LocalMux I__7643 (
            .O(N__41430),
            .I(N__41372));
    InMux I__7642 (
            .O(N__41429),
            .I(N__41369));
    InMux I__7641 (
            .O(N__41428),
            .I(N__41366));
    LocalMux I__7640 (
            .O(N__41423),
            .I(N__41358));
    LocalMux I__7639 (
            .O(N__41414),
            .I(N__41358));
    LocalMux I__7638 (
            .O(N__41405),
            .I(N__41358));
    InMux I__7637 (
            .O(N__41404),
            .I(N__41355));
    InMux I__7636 (
            .O(N__41403),
            .I(N__41352));
    Span4Mux_v I__7635 (
            .O(N__41400),
            .I(N__41345));
    Span4Mux_v I__7634 (
            .O(N__41397),
            .I(N__41345));
    LocalMux I__7633 (
            .O(N__41394),
            .I(N__41345));
    InMux I__7632 (
            .O(N__41393),
            .I(N__41342));
    Span4Mux_h I__7631 (
            .O(N__41390),
            .I(N__41339));
    Span4Mux_h I__7630 (
            .O(N__41387),
            .I(N__41330));
    Span4Mux_v I__7629 (
            .O(N__41384),
            .I(N__41330));
    LocalMux I__7628 (
            .O(N__41381),
            .I(N__41330));
    LocalMux I__7627 (
            .O(N__41378),
            .I(N__41330));
    LocalMux I__7626 (
            .O(N__41375),
            .I(N__41327));
    Span4Mux_h I__7625 (
            .O(N__41372),
            .I(N__41320));
    LocalMux I__7624 (
            .O(N__41369),
            .I(N__41320));
    LocalMux I__7623 (
            .O(N__41366),
            .I(N__41320));
    InMux I__7622 (
            .O(N__41365),
            .I(N__41317));
    Span4Mux_v I__7621 (
            .O(N__41358),
            .I(N__41310));
    LocalMux I__7620 (
            .O(N__41355),
            .I(N__41310));
    LocalMux I__7619 (
            .O(N__41352),
            .I(N__41310));
    Sp12to4 I__7618 (
            .O(N__41345),
            .I(N__41305));
    LocalMux I__7617 (
            .O(N__41342),
            .I(N__41305));
    Span4Mux_h I__7616 (
            .O(N__41339),
            .I(N__41298));
    Span4Mux_h I__7615 (
            .O(N__41330),
            .I(N__41298));
    Span4Mux_h I__7614 (
            .O(N__41327),
            .I(N__41298));
    Span4Mux_v I__7613 (
            .O(N__41320),
            .I(N__41291));
    LocalMux I__7612 (
            .O(N__41317),
            .I(N__41291));
    Span4Mux_h I__7611 (
            .O(N__41310),
            .I(N__41291));
    Odrv12 I__7610 (
            .O(N__41305),
            .I(\c0.n14 ));
    Odrv4 I__7609 (
            .O(N__41298),
            .I(\c0.n14 ));
    Odrv4 I__7608 (
            .O(N__41291),
            .I(\c0.n14 ));
    SRMux I__7607 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__7606 (
            .O(N__41281),
            .I(N__41278));
    Odrv12 I__7605 (
            .O(N__41278),
            .I(\c0.n18667 ));
    CascadeMux I__7604 (
            .O(N__41275),
            .I(N__41272));
    InMux I__7603 (
            .O(N__41272),
            .I(N__41269));
    LocalMux I__7602 (
            .O(N__41269),
            .I(N__41266));
    Span4Mux_h I__7601 (
            .O(N__41266),
            .I(N__41263));
    Odrv4 I__7600 (
            .O(N__41263),
            .I(\c0.n94 ));
    InMux I__7599 (
            .O(N__41260),
            .I(N__41257));
    LocalMux I__7598 (
            .O(N__41257),
            .I(\c0.n12_adj_3004 ));
    InMux I__7597 (
            .O(N__41254),
            .I(N__41251));
    LocalMux I__7596 (
            .O(N__41251),
            .I(\c0.n20_adj_3539 ));
    CascadeMux I__7595 (
            .O(N__41248),
            .I(\c0.n12_adj_3001_cascade_ ));
    CascadeMux I__7594 (
            .O(N__41245),
            .I(\c0.n20403_cascade_ ));
    InMux I__7593 (
            .O(N__41242),
            .I(N__41239));
    LocalMux I__7592 (
            .O(N__41239),
            .I(\c0.n10_adj_3514 ));
    CascadeMux I__7591 (
            .O(N__41236),
            .I(\c0.n20398_cascade_ ));
    CascadeMux I__7590 (
            .O(N__41233),
            .I(N__41229));
    InMux I__7589 (
            .O(N__41232),
            .I(N__41224));
    InMux I__7588 (
            .O(N__41229),
            .I(N__41224));
    LocalMux I__7587 (
            .O(N__41224),
            .I(N__41221));
    Odrv4 I__7586 (
            .O(N__41221),
            .I(\c0.n4_adj_3071 ));
    InMux I__7585 (
            .O(N__41218),
            .I(N__41213));
    InMux I__7584 (
            .O(N__41217),
            .I(N__41208));
    InMux I__7583 (
            .O(N__41216),
            .I(N__41208));
    LocalMux I__7582 (
            .O(N__41213),
            .I(\c0.n5_adj_3003 ));
    LocalMux I__7581 (
            .O(N__41208),
            .I(\c0.n5_adj_3003 ));
    CascadeMux I__7580 (
            .O(N__41203),
            .I(\c0.n36_adj_3267_cascade_ ));
    InMux I__7579 (
            .O(N__41200),
            .I(N__41197));
    LocalMux I__7578 (
            .O(N__41197),
            .I(\c0.n6_adj_3005 ));
    CascadeMux I__7577 (
            .O(N__41194),
            .I(N__41191));
    InMux I__7576 (
            .O(N__41191),
            .I(N__41185));
    InMux I__7575 (
            .O(N__41190),
            .I(N__41185));
    LocalMux I__7574 (
            .O(N__41185),
            .I(\c0.n13 ));
    CascadeMux I__7573 (
            .O(N__41182),
            .I(\c0.n36_adj_3547_cascade_ ));
    InMux I__7572 (
            .O(N__41179),
            .I(N__41176));
    LocalMux I__7571 (
            .O(N__41176),
            .I(N__41173));
    Span4Mux_v I__7570 (
            .O(N__41173),
            .I(N__41170));
    Odrv4 I__7569 (
            .O(N__41170),
            .I(\c0.n63_adj_3417 ));
    CascadeMux I__7568 (
            .O(N__41167),
            .I(\c0.n38_adj_3548_cascade_ ));
    InMux I__7567 (
            .O(N__41164),
            .I(N__41161));
    LocalMux I__7566 (
            .O(N__41161),
            .I(N__41158));
    Span4Mux_h I__7565 (
            .O(N__41158),
            .I(N__41155));
    Odrv4 I__7564 (
            .O(N__41155),
            .I(\c0.n34_adj_3411 ));
    CascadeMux I__7563 (
            .O(N__41152),
            .I(\c0.n18443_cascade_ ));
    InMux I__7562 (
            .O(N__41149),
            .I(N__41146));
    LocalMux I__7561 (
            .O(N__41146),
            .I(\c0.n25_adj_3495 ));
    InMux I__7560 (
            .O(N__41143),
            .I(N__41138));
    InMux I__7559 (
            .O(N__41142),
            .I(N__41135));
    InMux I__7558 (
            .O(N__41141),
            .I(N__41132));
    LocalMux I__7557 (
            .O(N__41138),
            .I(N__41128));
    LocalMux I__7556 (
            .O(N__41135),
            .I(N__41125));
    LocalMux I__7555 (
            .O(N__41132),
            .I(N__41121));
    InMux I__7554 (
            .O(N__41131),
            .I(N__41118));
    Span4Mux_v I__7553 (
            .O(N__41128),
            .I(N__41113));
    Span4Mux_v I__7552 (
            .O(N__41125),
            .I(N__41113));
    InMux I__7551 (
            .O(N__41124),
            .I(N__41110));
    Odrv4 I__7550 (
            .O(N__41121),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__7549 (
            .O(N__41118),
            .I(\c0.data_in_frame_9_4 ));
    Odrv4 I__7548 (
            .O(N__41113),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__7547 (
            .O(N__41110),
            .I(\c0.data_in_frame_9_4 ));
    CascadeMux I__7546 (
            .O(N__41101),
            .I(\c0.n25_adj_3495_cascade_ ));
    CascadeMux I__7545 (
            .O(N__41098),
            .I(N__41091));
    CascadeMux I__7544 (
            .O(N__41097),
            .I(N__41088));
    InMux I__7543 (
            .O(N__41096),
            .I(N__41083));
    InMux I__7542 (
            .O(N__41095),
            .I(N__41080));
    InMux I__7541 (
            .O(N__41094),
            .I(N__41077));
    InMux I__7540 (
            .O(N__41091),
            .I(N__41068));
    InMux I__7539 (
            .O(N__41088),
            .I(N__41068));
    InMux I__7538 (
            .O(N__41087),
            .I(N__41068));
    InMux I__7537 (
            .O(N__41086),
            .I(N__41068));
    LocalMux I__7536 (
            .O(N__41083),
            .I(n21222));
    LocalMux I__7535 (
            .O(N__41080),
            .I(n21222));
    LocalMux I__7534 (
            .O(N__41077),
            .I(n21222));
    LocalMux I__7533 (
            .O(N__41068),
            .I(n21222));
    InMux I__7532 (
            .O(N__41059),
            .I(N__41056));
    LocalMux I__7531 (
            .O(N__41056),
            .I(N__41053));
    Span4Mux_h I__7530 (
            .O(N__41053),
            .I(N__41050));
    Span4Mux_h I__7529 (
            .O(N__41050),
            .I(N__41046));
    InMux I__7528 (
            .O(N__41049),
            .I(N__41043));
    Odrv4 I__7527 (
            .O(N__41046),
            .I(control_mode_1));
    LocalMux I__7526 (
            .O(N__41043),
            .I(control_mode_1));
    InMux I__7525 (
            .O(N__41038),
            .I(N__41035));
    LocalMux I__7524 (
            .O(N__41035),
            .I(\c0.n16_adj_3018 ));
    CascadeMux I__7523 (
            .O(N__41032),
            .I(\c0.n32_adj_3493_cascade_ ));
    InMux I__7522 (
            .O(N__41029),
            .I(N__41024));
    InMux I__7521 (
            .O(N__41028),
            .I(N__41019));
    InMux I__7520 (
            .O(N__41027),
            .I(N__41019));
    LocalMux I__7519 (
            .O(N__41024),
            .I(\c0.n20209 ));
    LocalMux I__7518 (
            .O(N__41019),
            .I(\c0.n20209 ));
    InMux I__7517 (
            .O(N__41014),
            .I(N__41011));
    LocalMux I__7516 (
            .O(N__41011),
            .I(N__41008));
    Odrv4 I__7515 (
            .O(N__41008),
            .I(\c0.n20204 ));
    CascadeMux I__7514 (
            .O(N__41005),
            .I(\c0.n19217_cascade_ ));
    InMux I__7513 (
            .O(N__41002),
            .I(N__40996));
    InMux I__7512 (
            .O(N__41001),
            .I(N__40996));
    LocalMux I__7511 (
            .O(N__40996),
            .I(N__40992));
    InMux I__7510 (
            .O(N__40995),
            .I(N__40989));
    Odrv12 I__7509 (
            .O(N__40992),
            .I(\c0.n66 ));
    LocalMux I__7508 (
            .O(N__40989),
            .I(\c0.n66 ));
    CascadeMux I__7507 (
            .O(N__40984),
            .I(\c0.data_out_frame_28__0__N_708_cascade_ ));
    InMux I__7506 (
            .O(N__40981),
            .I(N__40978));
    LocalMux I__7505 (
            .O(N__40978),
            .I(\c0.data_out_frame_28__0__N_708 ));
    InMux I__7504 (
            .O(N__40975),
            .I(N__40972));
    LocalMux I__7503 (
            .O(N__40972),
            .I(N__40969));
    Span12Mux_v I__7502 (
            .O(N__40969),
            .I(N__40966));
    Odrv12 I__7501 (
            .O(N__40966),
            .I(\c0.data_out_frame_29_0 ));
    InMux I__7500 (
            .O(N__40963),
            .I(N__40960));
    LocalMux I__7499 (
            .O(N__40960),
            .I(\c0.data_out_frame_29_1 ));
    InMux I__7498 (
            .O(N__40957),
            .I(N__40953));
    InMux I__7497 (
            .O(N__40956),
            .I(N__40950));
    LocalMux I__7496 (
            .O(N__40953),
            .I(N__40945));
    LocalMux I__7495 (
            .O(N__40950),
            .I(N__40945));
    Odrv4 I__7494 (
            .O(N__40945),
            .I(data_out_frame_28_1));
    InMux I__7493 (
            .O(N__40942),
            .I(N__40939));
    LocalMux I__7492 (
            .O(N__40939),
            .I(N__40932));
    InMux I__7491 (
            .O(N__40938),
            .I(N__40927));
    InMux I__7490 (
            .O(N__40937),
            .I(N__40927));
    CascadeMux I__7489 (
            .O(N__40936),
            .I(N__40920));
    InMux I__7488 (
            .O(N__40935),
            .I(N__40916));
    Span4Mux_v I__7487 (
            .O(N__40932),
            .I(N__40909));
    LocalMux I__7486 (
            .O(N__40927),
            .I(N__40909));
    InMux I__7485 (
            .O(N__40926),
            .I(N__40901));
    InMux I__7484 (
            .O(N__40925),
            .I(N__40897));
    InMux I__7483 (
            .O(N__40924),
            .I(N__40894));
    InMux I__7482 (
            .O(N__40923),
            .I(N__40887));
    InMux I__7481 (
            .O(N__40920),
            .I(N__40887));
    InMux I__7480 (
            .O(N__40919),
            .I(N__40877));
    LocalMux I__7479 (
            .O(N__40916),
            .I(N__40874));
    InMux I__7478 (
            .O(N__40915),
            .I(N__40869));
    InMux I__7477 (
            .O(N__40914),
            .I(N__40869));
    Span4Mux_v I__7476 (
            .O(N__40909),
            .I(N__40866));
    InMux I__7475 (
            .O(N__40908),
            .I(N__40861));
    InMux I__7474 (
            .O(N__40907),
            .I(N__40861));
    InMux I__7473 (
            .O(N__40906),
            .I(N__40858));
    InMux I__7472 (
            .O(N__40905),
            .I(N__40850));
    InMux I__7471 (
            .O(N__40904),
            .I(N__40847));
    LocalMux I__7470 (
            .O(N__40901),
            .I(N__40841));
    InMux I__7469 (
            .O(N__40900),
            .I(N__40838));
    LocalMux I__7468 (
            .O(N__40897),
            .I(N__40833));
    LocalMux I__7467 (
            .O(N__40894),
            .I(N__40833));
    InMux I__7466 (
            .O(N__40893),
            .I(N__40830));
    InMux I__7465 (
            .O(N__40892),
            .I(N__40827));
    LocalMux I__7464 (
            .O(N__40887),
            .I(N__40820));
    InMux I__7463 (
            .O(N__40886),
            .I(N__40817));
    InMux I__7462 (
            .O(N__40885),
            .I(N__40814));
    InMux I__7461 (
            .O(N__40884),
            .I(N__40811));
    InMux I__7460 (
            .O(N__40883),
            .I(N__40806));
    InMux I__7459 (
            .O(N__40882),
            .I(N__40806));
    InMux I__7458 (
            .O(N__40881),
            .I(N__40801));
    InMux I__7457 (
            .O(N__40880),
            .I(N__40801));
    LocalMux I__7456 (
            .O(N__40877),
            .I(N__40794));
    Span4Mux_v I__7455 (
            .O(N__40874),
            .I(N__40794));
    LocalMux I__7454 (
            .O(N__40869),
            .I(N__40794));
    Span4Mux_h I__7453 (
            .O(N__40866),
            .I(N__40787));
    LocalMux I__7452 (
            .O(N__40861),
            .I(N__40787));
    LocalMux I__7451 (
            .O(N__40858),
            .I(N__40787));
    InMux I__7450 (
            .O(N__40857),
            .I(N__40784));
    InMux I__7449 (
            .O(N__40856),
            .I(N__40781));
    InMux I__7448 (
            .O(N__40855),
            .I(N__40774));
    InMux I__7447 (
            .O(N__40854),
            .I(N__40774));
    InMux I__7446 (
            .O(N__40853),
            .I(N__40774));
    LocalMux I__7445 (
            .O(N__40850),
            .I(N__40771));
    LocalMux I__7444 (
            .O(N__40847),
            .I(N__40768));
    InMux I__7443 (
            .O(N__40846),
            .I(N__40761));
    InMux I__7442 (
            .O(N__40845),
            .I(N__40761));
    InMux I__7441 (
            .O(N__40844),
            .I(N__40761));
    Span4Mux_h I__7440 (
            .O(N__40841),
            .I(N__40754));
    LocalMux I__7439 (
            .O(N__40838),
            .I(N__40754));
    Span4Mux_v I__7438 (
            .O(N__40833),
            .I(N__40754));
    LocalMux I__7437 (
            .O(N__40830),
            .I(N__40749));
    LocalMux I__7436 (
            .O(N__40827),
            .I(N__40749));
    InMux I__7435 (
            .O(N__40826),
            .I(N__40746));
    CascadeMux I__7434 (
            .O(N__40825),
            .I(N__40743));
    InMux I__7433 (
            .O(N__40824),
            .I(N__40740));
    InMux I__7432 (
            .O(N__40823),
            .I(N__40735));
    Span4Mux_v I__7431 (
            .O(N__40820),
            .I(N__40732));
    LocalMux I__7430 (
            .O(N__40817),
            .I(N__40729));
    LocalMux I__7429 (
            .O(N__40814),
            .I(N__40716));
    LocalMux I__7428 (
            .O(N__40811),
            .I(N__40716));
    LocalMux I__7427 (
            .O(N__40806),
            .I(N__40716));
    LocalMux I__7426 (
            .O(N__40801),
            .I(N__40716));
    Span4Mux_h I__7425 (
            .O(N__40794),
            .I(N__40716));
    Span4Mux_h I__7424 (
            .O(N__40787),
            .I(N__40716));
    LocalMux I__7423 (
            .O(N__40784),
            .I(N__40707));
    LocalMux I__7422 (
            .O(N__40781),
            .I(N__40707));
    LocalMux I__7421 (
            .O(N__40774),
            .I(N__40707));
    Span4Mux_v I__7420 (
            .O(N__40771),
            .I(N__40707));
    Span4Mux_v I__7419 (
            .O(N__40768),
            .I(N__40696));
    LocalMux I__7418 (
            .O(N__40761),
            .I(N__40696));
    Span4Mux_v I__7417 (
            .O(N__40754),
            .I(N__40696));
    Span4Mux_h I__7416 (
            .O(N__40749),
            .I(N__40696));
    LocalMux I__7415 (
            .O(N__40746),
            .I(N__40696));
    InMux I__7414 (
            .O(N__40743),
            .I(N__40693));
    LocalMux I__7413 (
            .O(N__40740),
            .I(N__40690));
    InMux I__7412 (
            .O(N__40739),
            .I(N__40687));
    InMux I__7411 (
            .O(N__40738),
            .I(N__40684));
    LocalMux I__7410 (
            .O(N__40735),
            .I(N__40679));
    Span4Mux_h I__7409 (
            .O(N__40732),
            .I(N__40679));
    Span4Mux_h I__7408 (
            .O(N__40729),
            .I(N__40674));
    Span4Mux_v I__7407 (
            .O(N__40716),
            .I(N__40674));
    Span4Mux_v I__7406 (
            .O(N__40707),
            .I(N__40669));
    Span4Mux_v I__7405 (
            .O(N__40696),
            .I(N__40669));
    LocalMux I__7404 (
            .O(N__40693),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7403 (
            .O(N__40690),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__7402 (
            .O(N__40687),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__7401 (
            .O(N__40684),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7400 (
            .O(N__40679),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7399 (
            .O(N__40674),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__7398 (
            .O(N__40669),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__7397 (
            .O(N__40654),
            .I(N__40651));
    LocalMux I__7396 (
            .O(N__40651),
            .I(N__40648));
    Span4Mux_v I__7395 (
            .O(N__40648),
            .I(N__40645));
    Odrv4 I__7394 (
            .O(N__40645),
            .I(\c0.n26_adj_3103 ));
    CascadeMux I__7393 (
            .O(N__40642),
            .I(\c0.n20246_cascade_ ));
    CascadeMux I__7392 (
            .O(N__40639),
            .I(N__40636));
    InMux I__7391 (
            .O(N__40636),
            .I(N__40633));
    LocalMux I__7390 (
            .O(N__40633),
            .I(\c0.n24_adj_3327 ));
    CascadeMux I__7389 (
            .O(N__40630),
            .I(\c0.n23_adj_3039_cascade_ ));
    InMux I__7388 (
            .O(N__40627),
            .I(N__40624));
    LocalMux I__7387 (
            .O(N__40624),
            .I(\c0.n23_adj_3039 ));
    InMux I__7386 (
            .O(N__40621),
            .I(N__40618));
    LocalMux I__7385 (
            .O(N__40618),
            .I(\c0.n30_adj_3042 ));
    CascadeMux I__7384 (
            .O(N__40615),
            .I(N__40611));
    InMux I__7383 (
            .O(N__40614),
            .I(N__40608));
    InMux I__7382 (
            .O(N__40611),
            .I(N__40605));
    LocalMux I__7381 (
            .O(N__40608),
            .I(data_out_frame_29_2));
    LocalMux I__7380 (
            .O(N__40605),
            .I(data_out_frame_29_2));
    CascadeMux I__7379 (
            .O(N__40600),
            .I(\c0.n18428_cascade_ ));
    InMux I__7378 (
            .O(N__40597),
            .I(N__40594));
    LocalMux I__7377 (
            .O(N__40594),
            .I(\c0.n29_adj_3446 ));
    InMux I__7376 (
            .O(N__40591),
            .I(N__40587));
    InMux I__7375 (
            .O(N__40590),
            .I(N__40584));
    LocalMux I__7374 (
            .O(N__40587),
            .I(data_out_frame_28_2));
    LocalMux I__7373 (
            .O(N__40584),
            .I(data_out_frame_28_2));
    InMux I__7372 (
            .O(N__40579),
            .I(N__40576));
    LocalMux I__7371 (
            .O(N__40576),
            .I(N__40570));
    InMux I__7370 (
            .O(N__40575),
            .I(N__40567));
    InMux I__7369 (
            .O(N__40574),
            .I(N__40562));
    InMux I__7368 (
            .O(N__40573),
            .I(N__40562));
    Odrv4 I__7367 (
            .O(N__40570),
            .I(data_in_0_5));
    LocalMux I__7366 (
            .O(N__40567),
            .I(data_in_0_5));
    LocalMux I__7365 (
            .O(N__40562),
            .I(data_in_0_5));
    InMux I__7364 (
            .O(N__40555),
            .I(N__40537));
    InMux I__7363 (
            .O(N__40554),
            .I(N__40534));
    InMux I__7362 (
            .O(N__40553),
            .I(N__40530));
    InMux I__7361 (
            .O(N__40552),
            .I(N__40519));
    InMux I__7360 (
            .O(N__40551),
            .I(N__40516));
    InMux I__7359 (
            .O(N__40550),
            .I(N__40512));
    InMux I__7358 (
            .O(N__40549),
            .I(N__40509));
    InMux I__7357 (
            .O(N__40548),
            .I(N__40506));
    InMux I__7356 (
            .O(N__40547),
            .I(N__40503));
    InMux I__7355 (
            .O(N__40546),
            .I(N__40500));
    InMux I__7354 (
            .O(N__40545),
            .I(N__40497));
    InMux I__7353 (
            .O(N__40544),
            .I(N__40494));
    InMux I__7352 (
            .O(N__40543),
            .I(N__40491));
    InMux I__7351 (
            .O(N__40542),
            .I(N__40487));
    InMux I__7350 (
            .O(N__40541),
            .I(N__40484));
    InMux I__7349 (
            .O(N__40540),
            .I(N__40481));
    LocalMux I__7348 (
            .O(N__40537),
            .I(N__40477));
    LocalMux I__7347 (
            .O(N__40534),
            .I(N__40474));
    InMux I__7346 (
            .O(N__40533),
            .I(N__40471));
    LocalMux I__7345 (
            .O(N__40530),
            .I(N__40468));
    InMux I__7344 (
            .O(N__40529),
            .I(N__40465));
    InMux I__7343 (
            .O(N__40528),
            .I(N__40462));
    InMux I__7342 (
            .O(N__40527),
            .I(N__40459));
    InMux I__7341 (
            .O(N__40526),
            .I(N__40456));
    InMux I__7340 (
            .O(N__40525),
            .I(N__40453));
    InMux I__7339 (
            .O(N__40524),
            .I(N__40450));
    InMux I__7338 (
            .O(N__40523),
            .I(N__40447));
    InMux I__7337 (
            .O(N__40522),
            .I(N__40444));
    LocalMux I__7336 (
            .O(N__40519),
            .I(N__40440));
    LocalMux I__7335 (
            .O(N__40516),
            .I(N__40437));
    InMux I__7334 (
            .O(N__40515),
            .I(N__40434));
    LocalMux I__7333 (
            .O(N__40512),
            .I(N__40423));
    LocalMux I__7332 (
            .O(N__40509),
            .I(N__40423));
    LocalMux I__7331 (
            .O(N__40506),
            .I(N__40423));
    LocalMux I__7330 (
            .O(N__40503),
            .I(N__40423));
    LocalMux I__7329 (
            .O(N__40500),
            .I(N__40423));
    LocalMux I__7328 (
            .O(N__40497),
            .I(N__40420));
    LocalMux I__7327 (
            .O(N__40494),
            .I(N__40415));
    LocalMux I__7326 (
            .O(N__40491),
            .I(N__40415));
    InMux I__7325 (
            .O(N__40490),
            .I(N__40412));
    LocalMux I__7324 (
            .O(N__40487),
            .I(N__40409));
    LocalMux I__7323 (
            .O(N__40484),
            .I(N__40404));
    LocalMux I__7322 (
            .O(N__40481),
            .I(N__40404));
    InMux I__7321 (
            .O(N__40480),
            .I(N__40401));
    Span4Mux_v I__7320 (
            .O(N__40477),
            .I(N__40396));
    Span4Mux_v I__7319 (
            .O(N__40474),
            .I(N__40396));
    LocalMux I__7318 (
            .O(N__40471),
            .I(N__40393));
    Span4Mux_v I__7317 (
            .O(N__40468),
            .I(N__40374));
    LocalMux I__7316 (
            .O(N__40465),
            .I(N__40374));
    LocalMux I__7315 (
            .O(N__40462),
            .I(N__40374));
    LocalMux I__7314 (
            .O(N__40459),
            .I(N__40374));
    LocalMux I__7313 (
            .O(N__40456),
            .I(N__40374));
    LocalMux I__7312 (
            .O(N__40453),
            .I(N__40374));
    LocalMux I__7311 (
            .O(N__40450),
            .I(N__40374));
    LocalMux I__7310 (
            .O(N__40447),
            .I(N__40374));
    LocalMux I__7309 (
            .O(N__40444),
            .I(N__40374));
    InMux I__7308 (
            .O(N__40443),
            .I(N__40371));
    Span12Mux_s11_v I__7307 (
            .O(N__40440),
            .I(N__40368));
    Span4Mux_h I__7306 (
            .O(N__40437),
            .I(N__40365));
    LocalMux I__7305 (
            .O(N__40434),
            .I(N__40362));
    Span4Mux_v I__7304 (
            .O(N__40423),
            .I(N__40353));
    Span4Mux_h I__7303 (
            .O(N__40420),
            .I(N__40353));
    Span4Mux_h I__7302 (
            .O(N__40415),
            .I(N__40353));
    LocalMux I__7301 (
            .O(N__40412),
            .I(N__40353));
    Span4Mux_v I__7300 (
            .O(N__40409),
            .I(N__40346));
    Span4Mux_v I__7299 (
            .O(N__40404),
            .I(N__40346));
    LocalMux I__7298 (
            .O(N__40401),
            .I(N__40346));
    Span4Mux_h I__7297 (
            .O(N__40396),
            .I(N__40337));
    Span4Mux_v I__7296 (
            .O(N__40393),
            .I(N__40337));
    Span4Mux_v I__7295 (
            .O(N__40374),
            .I(N__40337));
    LocalMux I__7294 (
            .O(N__40371),
            .I(N__40337));
    Odrv12 I__7293 (
            .O(N__40368),
            .I(\c0.n5_adj_2999 ));
    Odrv4 I__7292 (
            .O(N__40365),
            .I(\c0.n5_adj_2999 ));
    Odrv12 I__7291 (
            .O(N__40362),
            .I(\c0.n5_adj_2999 ));
    Odrv4 I__7290 (
            .O(N__40353),
            .I(\c0.n5_adj_2999 ));
    Odrv4 I__7289 (
            .O(N__40346),
            .I(\c0.n5_adj_2999 ));
    Odrv4 I__7288 (
            .O(N__40337),
            .I(\c0.n5_adj_2999 ));
    InMux I__7287 (
            .O(N__40324),
            .I(N__40321));
    LocalMux I__7286 (
            .O(N__40321),
            .I(N__40318));
    Span4Mux_v I__7285 (
            .O(N__40318),
            .I(N__40313));
    InMux I__7284 (
            .O(N__40317),
            .I(N__40310));
    InMux I__7283 (
            .O(N__40316),
            .I(N__40307));
    Span4Mux_h I__7282 (
            .O(N__40313),
            .I(N__40304));
    LocalMux I__7281 (
            .O(N__40310),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__7280 (
            .O(N__40307),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__7279 (
            .O(N__40304),
            .I(\c0.FRAME_MATCHER_state_18 ));
    SRMux I__7278 (
            .O(N__40297),
            .I(N__40294));
    LocalMux I__7277 (
            .O(N__40294),
            .I(N__40291));
    Odrv12 I__7276 (
            .O(N__40291),
            .I(\c0.n18655 ));
    InMux I__7275 (
            .O(N__40288),
            .I(N__40281));
    InMux I__7274 (
            .O(N__40287),
            .I(N__40277));
    InMux I__7273 (
            .O(N__40286),
            .I(N__40274));
    InMux I__7272 (
            .O(N__40285),
            .I(N__40271));
    InMux I__7271 (
            .O(N__40284),
            .I(N__40268));
    LocalMux I__7270 (
            .O(N__40281),
            .I(N__40262));
    InMux I__7269 (
            .O(N__40280),
            .I(N__40259));
    LocalMux I__7268 (
            .O(N__40277),
            .I(N__40252));
    LocalMux I__7267 (
            .O(N__40274),
            .I(N__40252));
    LocalMux I__7266 (
            .O(N__40271),
            .I(N__40252));
    LocalMux I__7265 (
            .O(N__40268),
            .I(N__40249));
    InMux I__7264 (
            .O(N__40267),
            .I(N__40246));
    InMux I__7263 (
            .O(N__40266),
            .I(N__40243));
    CascadeMux I__7262 (
            .O(N__40265),
            .I(N__40240));
    Span4Mux_h I__7261 (
            .O(N__40262),
            .I(N__40237));
    LocalMux I__7260 (
            .O(N__40259),
            .I(N__40232));
    Span4Mux_v I__7259 (
            .O(N__40252),
            .I(N__40232));
    Span4Mux_h I__7258 (
            .O(N__40249),
            .I(N__40227));
    LocalMux I__7257 (
            .O(N__40246),
            .I(N__40227));
    LocalMux I__7256 (
            .O(N__40243),
            .I(N__40224));
    InMux I__7255 (
            .O(N__40240),
            .I(N__40221));
    Span4Mux_v I__7254 (
            .O(N__40237),
            .I(N__40216));
    Span4Mux_v I__7253 (
            .O(N__40232),
            .I(N__40216));
    Span4Mux_v I__7252 (
            .O(N__40227),
            .I(N__40213));
    Sp12to4 I__7251 (
            .O(N__40224),
            .I(N__40210));
    LocalMux I__7250 (
            .O(N__40221),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv4 I__7249 (
            .O(N__40216),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv4 I__7248 (
            .O(N__40213),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv12 I__7247 (
            .O(N__40210),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__7246 (
            .O(N__40201),
            .I(N__40196));
    InMux I__7245 (
            .O(N__40200),
            .I(N__40193));
    InMux I__7244 (
            .O(N__40199),
            .I(N__40190));
    LocalMux I__7243 (
            .O(N__40196),
            .I(N__40187));
    LocalMux I__7242 (
            .O(N__40193),
            .I(N__40182));
    LocalMux I__7241 (
            .O(N__40190),
            .I(N__40179));
    Span4Mux_v I__7240 (
            .O(N__40187),
            .I(N__40176));
    InMux I__7239 (
            .O(N__40186),
            .I(N__40170));
    InMux I__7238 (
            .O(N__40185),
            .I(N__40170));
    Span4Mux_h I__7237 (
            .O(N__40182),
            .I(N__40165));
    Span4Mux_h I__7236 (
            .O(N__40179),
            .I(N__40165));
    Span4Mux_v I__7235 (
            .O(N__40176),
            .I(N__40161));
    InMux I__7234 (
            .O(N__40175),
            .I(N__40158));
    LocalMux I__7233 (
            .O(N__40170),
            .I(N__40155));
    Sp12to4 I__7232 (
            .O(N__40165),
            .I(N__40152));
    InMux I__7231 (
            .O(N__40164),
            .I(N__40149));
    Span4Mux_v I__7230 (
            .O(N__40161),
            .I(N__40146));
    LocalMux I__7229 (
            .O(N__40158),
            .I(N__40143));
    Span4Mux_h I__7228 (
            .O(N__40155),
            .I(N__40140));
    Span12Mux_v I__7227 (
            .O(N__40152),
            .I(N__40137));
    LocalMux I__7226 (
            .O(N__40149),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv4 I__7225 (
            .O(N__40146),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv12 I__7224 (
            .O(N__40143),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv4 I__7223 (
            .O(N__40140),
            .I(\c0.FRAME_MATCHER_i_6 ));
    Odrv12 I__7222 (
            .O(N__40137),
            .I(\c0.FRAME_MATCHER_i_6 ));
    CascadeMux I__7221 (
            .O(N__40126),
            .I(N__40122));
    InMux I__7220 (
            .O(N__40125),
            .I(N__40119));
    InMux I__7219 (
            .O(N__40122),
            .I(N__40115));
    LocalMux I__7218 (
            .O(N__40119),
            .I(N__40112));
    CascadeMux I__7217 (
            .O(N__40118),
            .I(N__40107));
    LocalMux I__7216 (
            .O(N__40115),
            .I(N__40102));
    Span4Mux_v I__7215 (
            .O(N__40112),
            .I(N__40102));
    InMux I__7214 (
            .O(N__40111),
            .I(N__40099));
    InMux I__7213 (
            .O(N__40110),
            .I(N__40096));
    InMux I__7212 (
            .O(N__40107),
            .I(N__40093));
    Span4Mux_v I__7211 (
            .O(N__40102),
            .I(N__40085));
    LocalMux I__7210 (
            .O(N__40099),
            .I(N__40085));
    LocalMux I__7209 (
            .O(N__40096),
            .I(N__40085));
    LocalMux I__7208 (
            .O(N__40093),
            .I(N__40081));
    InMux I__7207 (
            .O(N__40092),
            .I(N__40078));
    Span4Mux_h I__7206 (
            .O(N__40085),
            .I(N__40075));
    CascadeMux I__7205 (
            .O(N__40084),
            .I(N__40072));
    Span4Mux_h I__7204 (
            .O(N__40081),
            .I(N__40068));
    LocalMux I__7203 (
            .O(N__40078),
            .I(N__40063));
    Sp12to4 I__7202 (
            .O(N__40075),
            .I(N__40063));
    InMux I__7201 (
            .O(N__40072),
            .I(N__40057));
    InMux I__7200 (
            .O(N__40071),
            .I(N__40057));
    Span4Mux_h I__7199 (
            .O(N__40068),
            .I(N__40054));
    Span12Mux_v I__7198 (
            .O(N__40063),
            .I(N__40051));
    InMux I__7197 (
            .O(N__40062),
            .I(N__40048));
    LocalMux I__7196 (
            .O(N__40057),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__7195 (
            .O(N__40054),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__7194 (
            .O(N__40051),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__7193 (
            .O(N__40048),
            .I(\c0.FRAME_MATCHER_i_3 ));
    CascadeMux I__7192 (
            .O(N__40039),
            .I(\c0.n20224_cascade_ ));
    CascadeMux I__7191 (
            .O(N__40036),
            .I(\c0.n19_cascade_ ));
    InMux I__7190 (
            .O(N__40033),
            .I(N__40027));
    InMux I__7189 (
            .O(N__40032),
            .I(N__40027));
    LocalMux I__7188 (
            .O(N__40027),
            .I(N__40022));
    InMux I__7187 (
            .O(N__40026),
            .I(N__40017));
    InMux I__7186 (
            .O(N__40025),
            .I(N__40017));
    Odrv4 I__7185 (
            .O(N__40022),
            .I(data_in_2_3));
    LocalMux I__7184 (
            .O(N__40017),
            .I(data_in_2_3));
    InMux I__7183 (
            .O(N__40012),
            .I(N__40009));
    LocalMux I__7182 (
            .O(N__40009),
            .I(N__40005));
    InMux I__7181 (
            .O(N__40008),
            .I(N__40000));
    Span4Mux_h I__7180 (
            .O(N__40005),
            .I(N__39997));
    InMux I__7179 (
            .O(N__40004),
            .I(N__39994));
    InMux I__7178 (
            .O(N__40003),
            .I(N__39991));
    LocalMux I__7177 (
            .O(N__40000),
            .I(data_in_1_3));
    Odrv4 I__7176 (
            .O(N__39997),
            .I(data_in_1_3));
    LocalMux I__7175 (
            .O(N__39994),
            .I(data_in_1_3));
    LocalMux I__7174 (
            .O(N__39991),
            .I(data_in_1_3));
    CascadeMux I__7173 (
            .O(N__39982),
            .I(N__39977));
    InMux I__7172 (
            .O(N__39981),
            .I(N__39974));
    InMux I__7171 (
            .O(N__39980),
            .I(N__39971));
    InMux I__7170 (
            .O(N__39977),
            .I(N__39968));
    LocalMux I__7169 (
            .O(N__39974),
            .I(data_in_0_6));
    LocalMux I__7168 (
            .O(N__39971),
            .I(data_in_0_6));
    LocalMux I__7167 (
            .O(N__39968),
            .I(data_in_0_6));
    InMux I__7166 (
            .O(N__39961),
            .I(N__39955));
    InMux I__7165 (
            .O(N__39960),
            .I(N__39955));
    LocalMux I__7164 (
            .O(N__39955),
            .I(N__39951));
    InMux I__7163 (
            .O(N__39954),
            .I(N__39948));
    Span4Mux_h I__7162 (
            .O(N__39951),
            .I(N__39945));
    LocalMux I__7161 (
            .O(N__39948),
            .I(data_in_0_3));
    Odrv4 I__7160 (
            .O(N__39945),
            .I(data_in_0_3));
    InMux I__7159 (
            .O(N__39940),
            .I(N__39937));
    LocalMux I__7158 (
            .O(N__39937),
            .I(\c0.n18_adj_3246 ));
    CascadeMux I__7157 (
            .O(N__39934),
            .I(\c0.n20_cascade_ ));
    InMux I__7156 (
            .O(N__39931),
            .I(N__39928));
    LocalMux I__7155 (
            .O(N__39928),
            .I(\c0.n16_adj_3247 ));
    InMux I__7154 (
            .O(N__39925),
            .I(N__39919));
    InMux I__7153 (
            .O(N__39924),
            .I(N__39919));
    LocalMux I__7152 (
            .O(N__39919),
            .I(\c0.n11311 ));
    CascadeMux I__7151 (
            .O(N__39916),
            .I(N__39910));
    InMux I__7150 (
            .O(N__39915),
            .I(N__39905));
    InMux I__7149 (
            .O(N__39914),
            .I(N__39905));
    InMux I__7148 (
            .O(N__39913),
            .I(N__39900));
    InMux I__7147 (
            .O(N__39910),
            .I(N__39900));
    LocalMux I__7146 (
            .O(N__39905),
            .I(data_in_3_2));
    LocalMux I__7145 (
            .O(N__39900),
            .I(data_in_3_2));
    CascadeMux I__7144 (
            .O(N__39895),
            .I(N__39892));
    InMux I__7143 (
            .O(N__39892),
            .I(N__39888));
    InMux I__7142 (
            .O(N__39891),
            .I(N__39885));
    LocalMux I__7141 (
            .O(N__39888),
            .I(N__39880));
    LocalMux I__7140 (
            .O(N__39885),
            .I(N__39880));
    Span4Mux_h I__7139 (
            .O(N__39880),
            .I(N__39876));
    InMux I__7138 (
            .O(N__39879),
            .I(N__39873));
    Odrv4 I__7137 (
            .O(N__39876),
            .I(\c0.n105 ));
    LocalMux I__7136 (
            .O(N__39873),
            .I(\c0.n105 ));
    InMux I__7135 (
            .O(N__39868),
            .I(N__39862));
    InMux I__7134 (
            .O(N__39867),
            .I(N__39857));
    InMux I__7133 (
            .O(N__39866),
            .I(N__39857));
    InMux I__7132 (
            .O(N__39865),
            .I(N__39854));
    LocalMux I__7131 (
            .O(N__39862),
            .I(data_in_3_3));
    LocalMux I__7130 (
            .O(N__39857),
            .I(data_in_3_3));
    LocalMux I__7129 (
            .O(N__39854),
            .I(data_in_3_3));
    InMux I__7128 (
            .O(N__39847),
            .I(N__39839));
    InMux I__7127 (
            .O(N__39846),
            .I(N__39839));
    InMux I__7126 (
            .O(N__39845),
            .I(N__39834));
    InMux I__7125 (
            .O(N__39844),
            .I(N__39834));
    LocalMux I__7124 (
            .O(N__39839),
            .I(data_in_3_1));
    LocalMux I__7123 (
            .O(N__39834),
            .I(data_in_3_1));
    CascadeMux I__7122 (
            .O(N__39829),
            .I(N__39825));
    CascadeMux I__7121 (
            .O(N__39828),
            .I(N__39821));
    InMux I__7120 (
            .O(N__39825),
            .I(N__39818));
    InMux I__7119 (
            .O(N__39824),
            .I(N__39813));
    InMux I__7118 (
            .O(N__39821),
            .I(N__39813));
    LocalMux I__7117 (
            .O(N__39818),
            .I(data_in_0_7));
    LocalMux I__7116 (
            .O(N__39813),
            .I(data_in_0_7));
    CascadeMux I__7115 (
            .O(N__39808),
            .I(N__39803));
    InMux I__7114 (
            .O(N__39807),
            .I(N__39799));
    InMux I__7113 (
            .O(N__39806),
            .I(N__39796));
    InMux I__7112 (
            .O(N__39803),
            .I(N__39793));
    InMux I__7111 (
            .O(N__39802),
            .I(N__39790));
    LocalMux I__7110 (
            .O(N__39799),
            .I(N__39787));
    LocalMux I__7109 (
            .O(N__39796),
            .I(N__39782));
    LocalMux I__7108 (
            .O(N__39793),
            .I(N__39782));
    LocalMux I__7107 (
            .O(N__39790),
            .I(data_in_1_6));
    Odrv4 I__7106 (
            .O(N__39787),
            .I(data_in_1_6));
    Odrv12 I__7105 (
            .O(N__39782),
            .I(data_in_1_6));
    InMux I__7104 (
            .O(N__39775),
            .I(N__39772));
    LocalMux I__7103 (
            .O(N__39772),
            .I(\c0.n18_adj_3229 ));
    CascadeMux I__7102 (
            .O(N__39769),
            .I(N__39766));
    InMux I__7101 (
            .O(N__39766),
            .I(N__39760));
    InMux I__7100 (
            .O(N__39765),
            .I(N__39760));
    LocalMux I__7099 (
            .O(N__39760),
            .I(N__39757));
    Odrv4 I__7098 (
            .O(N__39757),
            .I(\c0.n11446 ));
    CascadeMux I__7097 (
            .O(N__39754),
            .I(\c0.n21108_cascade_ ));
    InMux I__7096 (
            .O(N__39751),
            .I(N__39748));
    LocalMux I__7095 (
            .O(N__39748),
            .I(\c0.n12_adj_3248 ));
    InMux I__7094 (
            .O(N__39745),
            .I(N__39740));
    InMux I__7093 (
            .O(N__39744),
            .I(N__39736));
    InMux I__7092 (
            .O(N__39743),
            .I(N__39733));
    LocalMux I__7091 (
            .O(N__39740),
            .I(N__39730));
    InMux I__7090 (
            .O(N__39739),
            .I(N__39727));
    LocalMux I__7089 (
            .O(N__39736),
            .I(N__39724));
    LocalMux I__7088 (
            .O(N__39733),
            .I(N__39717));
    Span4Mux_v I__7087 (
            .O(N__39730),
            .I(N__39717));
    LocalMux I__7086 (
            .O(N__39727),
            .I(N__39717));
    Odrv12 I__7085 (
            .O(N__39724),
            .I(data_in_3_5));
    Odrv4 I__7084 (
            .O(N__39717),
            .I(data_in_3_5));
    InMux I__7083 (
            .O(N__39712),
            .I(N__39706));
    InMux I__7082 (
            .O(N__39711),
            .I(N__39706));
    LocalMux I__7081 (
            .O(N__39706),
            .I(\c0.n20_adj_3250 ));
    InMux I__7080 (
            .O(N__39703),
            .I(N__39699));
    CascadeMux I__7079 (
            .O(N__39702),
            .I(N__39696));
    LocalMux I__7078 (
            .O(N__39699),
            .I(N__39693));
    InMux I__7077 (
            .O(N__39696),
            .I(N__39690));
    Span4Mux_h I__7076 (
            .O(N__39693),
            .I(N__39687));
    LocalMux I__7075 (
            .O(N__39690),
            .I(\c0.data_in_frame_28_6 ));
    Odrv4 I__7074 (
            .O(N__39687),
            .I(\c0.data_in_frame_28_6 ));
    CascadeMux I__7073 (
            .O(N__39682),
            .I(\c0.n17947_cascade_ ));
    InMux I__7072 (
            .O(N__39679),
            .I(N__39676));
    LocalMux I__7071 (
            .O(N__39676),
            .I(N__39673));
    Odrv4 I__7070 (
            .O(N__39673),
            .I(\c0.n20793 ));
    CascadeMux I__7069 (
            .O(N__39670),
            .I(\c0.n10_adj_3242_cascade_ ));
    InMux I__7068 (
            .O(N__39667),
            .I(N__39662));
    InMux I__7067 (
            .O(N__39666),
            .I(N__39659));
    InMux I__7066 (
            .O(N__39665),
            .I(N__39656));
    LocalMux I__7065 (
            .O(N__39662),
            .I(data_in_0_2));
    LocalMux I__7064 (
            .O(N__39659),
            .I(data_in_0_2));
    LocalMux I__7063 (
            .O(N__39656),
            .I(data_in_0_2));
    InMux I__7062 (
            .O(N__39649),
            .I(N__39646));
    LocalMux I__7061 (
            .O(N__39646),
            .I(\c0.n14_adj_3243 ));
    CascadeMux I__7060 (
            .O(N__39643),
            .I(\c0.n36_adj_3277_cascade_ ));
    CascadeMux I__7059 (
            .O(N__39640),
            .I(\c0.n20415_cascade_ ));
    CascadeMux I__7058 (
            .O(N__39637),
            .I(\c0.n14_adj_3407_cascade_ ));
    InMux I__7057 (
            .O(N__39634),
            .I(N__39631));
    LocalMux I__7056 (
            .O(N__39631),
            .I(\c0.n100_adj_3403 ));
    CascadeMux I__7055 (
            .O(N__39628),
            .I(N__39625));
    InMux I__7054 (
            .O(N__39625),
            .I(N__39622));
    LocalMux I__7053 (
            .O(N__39622),
            .I(N__39619));
    Span4Mux_h I__7052 (
            .O(N__39619),
            .I(N__39616));
    Span4Mux_v I__7051 (
            .O(N__39616),
            .I(N__39613));
    Odrv4 I__7050 (
            .O(N__39613),
            .I(\c0.n18_adj_3412 ));
    CascadeMux I__7049 (
            .O(N__39610),
            .I(\c0.n20300_cascade_ ));
    CascadeMux I__7048 (
            .O(N__39607),
            .I(N__39604));
    InMux I__7047 (
            .O(N__39604),
            .I(N__39601));
    LocalMux I__7046 (
            .O(N__39601),
            .I(\c0.n20300 ));
    CascadeMux I__7045 (
            .O(N__39598),
            .I(N__39591));
    CascadeMux I__7044 (
            .O(N__39597),
            .I(N__39587));
    InMux I__7043 (
            .O(N__39596),
            .I(N__39582));
    InMux I__7042 (
            .O(N__39595),
            .I(N__39582));
    InMux I__7041 (
            .O(N__39594),
            .I(N__39577));
    InMux I__7040 (
            .O(N__39591),
            .I(N__39577));
    InMux I__7039 (
            .O(N__39590),
            .I(N__39573));
    InMux I__7038 (
            .O(N__39587),
            .I(N__39570));
    LocalMux I__7037 (
            .O(N__39582),
            .I(N__39564));
    LocalMux I__7036 (
            .O(N__39577),
            .I(N__39561));
    InMux I__7035 (
            .O(N__39576),
            .I(N__39558));
    LocalMux I__7034 (
            .O(N__39573),
            .I(N__39553));
    LocalMux I__7033 (
            .O(N__39570),
            .I(N__39549));
    InMux I__7032 (
            .O(N__39569),
            .I(N__39546));
    InMux I__7031 (
            .O(N__39568),
            .I(N__39543));
    InMux I__7030 (
            .O(N__39567),
            .I(N__39540));
    Span4Mux_v I__7029 (
            .O(N__39564),
            .I(N__39537));
    Span4Mux_h I__7028 (
            .O(N__39561),
            .I(N__39532));
    LocalMux I__7027 (
            .O(N__39558),
            .I(N__39532));
    InMux I__7026 (
            .O(N__39557),
            .I(N__39529));
    InMux I__7025 (
            .O(N__39556),
            .I(N__39526));
    Span4Mux_h I__7024 (
            .O(N__39553),
            .I(N__39523));
    InMux I__7023 (
            .O(N__39552),
            .I(N__39520));
    Span4Mux_h I__7022 (
            .O(N__39549),
            .I(N__39515));
    LocalMux I__7021 (
            .O(N__39546),
            .I(N__39515));
    LocalMux I__7020 (
            .O(N__39543),
            .I(N__39512));
    LocalMux I__7019 (
            .O(N__39540),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7018 (
            .O(N__39537),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7017 (
            .O(N__39532),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7016 (
            .O(N__39529),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7015 (
            .O(N__39526),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7014 (
            .O(N__39523),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7013 (
            .O(N__39520),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7012 (
            .O(N__39515),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7011 (
            .O(N__39512),
            .I(\c0.FRAME_MATCHER_state_0 ));
    InMux I__7010 (
            .O(N__39493),
            .I(N__39487));
    InMux I__7009 (
            .O(N__39492),
            .I(N__39483));
    InMux I__7008 (
            .O(N__39491),
            .I(N__39478));
    InMux I__7007 (
            .O(N__39490),
            .I(N__39478));
    LocalMux I__7006 (
            .O(N__39487),
            .I(N__39475));
    InMux I__7005 (
            .O(N__39486),
            .I(N__39472));
    LocalMux I__7004 (
            .O(N__39483),
            .I(N__39469));
    LocalMux I__7003 (
            .O(N__39478),
            .I(N__39466));
    Span4Mux_v I__7002 (
            .O(N__39475),
            .I(N__39463));
    LocalMux I__7001 (
            .O(N__39472),
            .I(N__39460));
    Span4Mux_h I__7000 (
            .O(N__39469),
            .I(N__39457));
    Sp12to4 I__6999 (
            .O(N__39466),
            .I(N__39454));
    Span4Mux_v I__6998 (
            .O(N__39463),
            .I(N__39449));
    Span4Mux_h I__6997 (
            .O(N__39460),
            .I(N__39449));
    Span4Mux_h I__6996 (
            .O(N__39457),
            .I(N__39446));
    Span12Mux_v I__6995 (
            .O(N__39454),
            .I(N__39443));
    Span4Mux_h I__6994 (
            .O(N__39449),
            .I(N__39440));
    Odrv4 I__6993 (
            .O(N__39446),
            .I(\c0.n3235 ));
    Odrv12 I__6992 (
            .O(N__39443),
            .I(\c0.n3235 ));
    Odrv4 I__6991 (
            .O(N__39440),
            .I(\c0.n3235 ));
    InMux I__6990 (
            .O(N__39433),
            .I(N__39429));
    InMux I__6989 (
            .O(N__39432),
            .I(N__39426));
    LocalMux I__6988 (
            .O(N__39429),
            .I(N__39423));
    LocalMux I__6987 (
            .O(N__39426),
            .I(\c0.rx.n15860 ));
    Odrv4 I__6986 (
            .O(N__39423),
            .I(\c0.rx.n15860 ));
    InMux I__6985 (
            .O(N__39418),
            .I(N__39415));
    LocalMux I__6984 (
            .O(N__39415),
            .I(N__39412));
    Span4Mux_v I__6983 (
            .O(N__39412),
            .I(N__39409));
    Odrv4 I__6982 (
            .O(N__39409),
            .I(\c0.n19449 ));
    InMux I__6981 (
            .O(N__39406),
            .I(N__39403));
    LocalMux I__6980 (
            .O(N__39403),
            .I(N__39398));
    InMux I__6979 (
            .O(N__39402),
            .I(N__39393));
    InMux I__6978 (
            .O(N__39401),
            .I(N__39393));
    Span12Mux_h I__6977 (
            .O(N__39398),
            .I(N__39390));
    LocalMux I__6976 (
            .O(N__39393),
            .I(N__39387));
    Odrv12 I__6975 (
            .O(N__39390),
            .I(n12492));
    Odrv4 I__6974 (
            .O(N__39387),
            .I(n12492));
    CascadeMux I__6973 (
            .O(N__39382),
            .I(N__39379));
    InMux I__6972 (
            .O(N__39379),
            .I(N__39376));
    LocalMux I__6971 (
            .O(N__39376),
            .I(N__39371));
    InMux I__6970 (
            .O(N__39375),
            .I(N__39366));
    InMux I__6969 (
            .O(N__39374),
            .I(N__39366));
    Span4Mux_h I__6968 (
            .O(N__39371),
            .I(N__39363));
    LocalMux I__6967 (
            .O(N__39366),
            .I(N__39360));
    Sp12to4 I__6966 (
            .O(N__39363),
            .I(N__39357));
    Odrv12 I__6965 (
            .O(N__39360),
            .I(n12835));
    Odrv12 I__6964 (
            .O(N__39357),
            .I(n12835));
    InMux I__6963 (
            .O(N__39352),
            .I(N__39349));
    LocalMux I__6962 (
            .O(N__39349),
            .I(N__39346));
    Span4Mux_h I__6961 (
            .O(N__39346),
            .I(N__39339));
    InMux I__6960 (
            .O(N__39345),
            .I(N__39336));
    InMux I__6959 (
            .O(N__39344),
            .I(N__39328));
    InMux I__6958 (
            .O(N__39343),
            .I(N__39328));
    InMux I__6957 (
            .O(N__39342),
            .I(N__39328));
    Span4Mux_v I__6956 (
            .O(N__39339),
            .I(N__39325));
    LocalMux I__6955 (
            .O(N__39336),
            .I(N__39322));
    InMux I__6954 (
            .O(N__39335),
            .I(N__39319));
    LocalMux I__6953 (
            .O(N__39328),
            .I(N__39314));
    Span4Mux_v I__6952 (
            .O(N__39325),
            .I(N__39314));
    Odrv12 I__6951 (
            .O(N__39322),
            .I(r_Bit_Index_0));
    LocalMux I__6950 (
            .O(N__39319),
            .I(r_Bit_Index_0));
    Odrv4 I__6949 (
            .O(N__39314),
            .I(r_Bit_Index_0));
    CascadeMux I__6948 (
            .O(N__39307),
            .I(\c0.n22_adj_3276_cascade_ ));
    InMux I__6947 (
            .O(N__39304),
            .I(N__39301));
    LocalMux I__6946 (
            .O(N__39301),
            .I(N__39298));
    Odrv12 I__6945 (
            .O(N__39298),
            .I(\c0.n21104 ));
    CascadeMux I__6944 (
            .O(N__39295),
            .I(n3846_cascade_));
    InMux I__6943 (
            .O(N__39292),
            .I(N__39286));
    InMux I__6942 (
            .O(N__39291),
            .I(N__39280));
    InMux I__6941 (
            .O(N__39290),
            .I(N__39277));
    InMux I__6940 (
            .O(N__39289),
            .I(N__39274));
    LocalMux I__6939 (
            .O(N__39286),
            .I(N__39271));
    InMux I__6938 (
            .O(N__39285),
            .I(N__39264));
    InMux I__6937 (
            .O(N__39284),
            .I(N__39264));
    InMux I__6936 (
            .O(N__39283),
            .I(N__39264));
    LocalMux I__6935 (
            .O(N__39280),
            .I(N__39261));
    LocalMux I__6934 (
            .O(N__39277),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__6933 (
            .O(N__39274),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__6932 (
            .O(N__39271),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__6931 (
            .O(N__39264),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__6930 (
            .O(N__39261),
            .I(\c0.rx.r_Clock_Count_7 ));
    InMux I__6929 (
            .O(N__39250),
            .I(N__39247));
    LocalMux I__6928 (
            .O(N__39247),
            .I(\c0.rx.n6_adj_2995 ));
    InMux I__6927 (
            .O(N__39244),
            .I(N__39240));
    InMux I__6926 (
            .O(N__39243),
            .I(N__39237));
    LocalMux I__6925 (
            .O(N__39240),
            .I(\c0.rx.n11455 ));
    LocalMux I__6924 (
            .O(N__39237),
            .I(\c0.rx.n11455 ));
    InMux I__6923 (
            .O(N__39232),
            .I(N__39228));
    InMux I__6922 (
            .O(N__39231),
            .I(N__39225));
    LocalMux I__6921 (
            .O(N__39228),
            .I(N__39222));
    LocalMux I__6920 (
            .O(N__39225),
            .I(N__39216));
    Span4Mux_v I__6919 (
            .O(N__39222),
            .I(N__39216));
    InMux I__6918 (
            .O(N__39221),
            .I(N__39213));
    Span4Mux_h I__6917 (
            .O(N__39216),
            .I(N__39210));
    LocalMux I__6916 (
            .O(N__39213),
            .I(\c0.rx.r_SM_Main_2_N_2479_0 ));
    Odrv4 I__6915 (
            .O(N__39210),
            .I(\c0.rx.r_SM_Main_2_N_2479_0 ));
    InMux I__6914 (
            .O(N__39205),
            .I(N__39199));
    InMux I__6913 (
            .O(N__39204),
            .I(N__39199));
    LocalMux I__6912 (
            .O(N__39199),
            .I(N__39196));
    Span4Mux_v I__6911 (
            .O(N__39196),
            .I(N__39187));
    InMux I__6910 (
            .O(N__39195),
            .I(N__39184));
    InMux I__6909 (
            .O(N__39194),
            .I(N__39177));
    InMux I__6908 (
            .O(N__39193),
            .I(N__39177));
    InMux I__6907 (
            .O(N__39192),
            .I(N__39177));
    InMux I__6906 (
            .O(N__39191),
            .I(N__39172));
    InMux I__6905 (
            .O(N__39190),
            .I(N__39172));
    Odrv4 I__6904 (
            .O(N__39187),
            .I(n3792));
    LocalMux I__6903 (
            .O(N__39184),
            .I(n3792));
    LocalMux I__6902 (
            .O(N__39177),
            .I(n3792));
    LocalMux I__6901 (
            .O(N__39172),
            .I(n3792));
    InMux I__6900 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__6899 (
            .O(N__39160),
            .I(N__39157));
    Span4Mux_h I__6898 (
            .O(N__39157),
            .I(N__39154));
    Odrv4 I__6897 (
            .O(N__39154),
            .I(n12911));
    InMux I__6896 (
            .O(N__39151),
            .I(N__39147));
    InMux I__6895 (
            .O(N__39150),
            .I(N__39144));
    LocalMux I__6894 (
            .O(N__39147),
            .I(N__39137));
    LocalMux I__6893 (
            .O(N__39144),
            .I(N__39137));
    CascadeMux I__6892 (
            .O(N__39143),
            .I(N__39133));
    InMux I__6891 (
            .O(N__39142),
            .I(N__39130));
    Span4Mux_h I__6890 (
            .O(N__39137),
            .I(N__39127));
    InMux I__6889 (
            .O(N__39136),
            .I(N__39124));
    InMux I__6888 (
            .O(N__39133),
            .I(N__39121));
    LocalMux I__6887 (
            .O(N__39130),
            .I(\c0.rx.r_Clock_Count_3 ));
    Odrv4 I__6886 (
            .O(N__39127),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__6885 (
            .O(N__39124),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__6884 (
            .O(N__39121),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__6883 (
            .O(N__39112),
            .I(N__39109));
    LocalMux I__6882 (
            .O(N__39109),
            .I(\c0.n16 ));
    InMux I__6881 (
            .O(N__39106),
            .I(N__39103));
    LocalMux I__6880 (
            .O(N__39103),
            .I(\c0.n24 ));
    CascadeMux I__6879 (
            .O(N__39100),
            .I(\c0.n28_cascade_ ));
    CascadeMux I__6878 (
            .O(N__39097),
            .I(\c0.n12026_cascade_ ));
    CascadeMux I__6877 (
            .O(N__39094),
            .I(\c0.n10_cascade_ ));
    CascadeMux I__6876 (
            .O(N__39091),
            .I(\c0.n19449_cascade_ ));
    InMux I__6875 (
            .O(N__39088),
            .I(N__39084));
    InMux I__6874 (
            .O(N__39087),
            .I(N__39081));
    LocalMux I__6873 (
            .O(N__39084),
            .I(control_mode_0));
    LocalMux I__6872 (
            .O(N__39081),
            .I(control_mode_0));
    CascadeMux I__6871 (
            .O(N__39076),
            .I(N__39072));
    InMux I__6870 (
            .O(N__39075),
            .I(N__39068));
    InMux I__6869 (
            .O(N__39072),
            .I(N__39065));
    InMux I__6868 (
            .O(N__39071),
            .I(N__39061));
    LocalMux I__6867 (
            .O(N__39068),
            .I(N__39055));
    LocalMux I__6866 (
            .O(N__39065),
            .I(N__39055));
    InMux I__6865 (
            .O(N__39064),
            .I(N__39052));
    LocalMux I__6864 (
            .O(N__39061),
            .I(N__39049));
    InMux I__6863 (
            .O(N__39060),
            .I(N__39046));
    Span4Mux_v I__6862 (
            .O(N__39055),
            .I(N__39043));
    LocalMux I__6861 (
            .O(N__39052),
            .I(N__39040));
    Span4Mux_h I__6860 (
            .O(N__39049),
            .I(N__39037));
    LocalMux I__6859 (
            .O(N__39046),
            .I(N__39032));
    Span4Mux_h I__6858 (
            .O(N__39043),
            .I(N__39032));
    Span4Mux_v I__6857 (
            .O(N__39040),
            .I(N__39029));
    Sp12to4 I__6856 (
            .O(N__39037),
            .I(N__39026));
    Span4Mux_v I__6855 (
            .O(N__39032),
            .I(N__39023));
    Span4Mux_v I__6854 (
            .O(N__39029),
            .I(N__39020));
    Span12Mux_v I__6853 (
            .O(N__39026),
            .I(N__39017));
    Span4Mux_v I__6852 (
            .O(N__39023),
            .I(N__39014));
    Span4Mux_v I__6851 (
            .O(N__39020),
            .I(N__39011));
    Odrv12 I__6850 (
            .O(N__39017),
            .I(FRAME_MATCHER_state_31_N_1800_2));
    Odrv4 I__6849 (
            .O(N__39014),
            .I(FRAME_MATCHER_state_31_N_1800_2));
    Odrv4 I__6848 (
            .O(N__39011),
            .I(FRAME_MATCHER_state_31_N_1800_2));
    InMux I__6847 (
            .O(N__39004),
            .I(N__38998));
    InMux I__6846 (
            .O(N__39003),
            .I(N__38998));
    LocalMux I__6845 (
            .O(N__38998),
            .I(N__38993));
    InMux I__6844 (
            .O(N__38997),
            .I(N__38990));
    CascadeMux I__6843 (
            .O(N__38996),
            .I(N__38986));
    Span4Mux_h I__6842 (
            .O(N__38993),
            .I(N__38979));
    LocalMux I__6841 (
            .O(N__38990),
            .I(N__38979));
    CascadeMux I__6840 (
            .O(N__38989),
            .I(N__38973));
    InMux I__6839 (
            .O(N__38986),
            .I(N__38969));
    CascadeMux I__6838 (
            .O(N__38985),
            .I(N__38965));
    InMux I__6837 (
            .O(N__38984),
            .I(N__38961));
    Span4Mux_v I__6836 (
            .O(N__38979),
            .I(N__38958));
    InMux I__6835 (
            .O(N__38978),
            .I(N__38955));
    CascadeMux I__6834 (
            .O(N__38977),
            .I(N__38952));
    InMux I__6833 (
            .O(N__38976),
            .I(N__38947));
    InMux I__6832 (
            .O(N__38973),
            .I(N__38947));
    InMux I__6831 (
            .O(N__38972),
            .I(N__38944));
    LocalMux I__6830 (
            .O(N__38969),
            .I(N__38941));
    InMux I__6829 (
            .O(N__38968),
            .I(N__38938));
    InMux I__6828 (
            .O(N__38965),
            .I(N__38935));
    CascadeMux I__6827 (
            .O(N__38964),
            .I(N__38932));
    LocalMux I__6826 (
            .O(N__38961),
            .I(N__38928));
    Span4Mux_v I__6825 (
            .O(N__38958),
            .I(N__38922));
    LocalMux I__6824 (
            .O(N__38955),
            .I(N__38919));
    InMux I__6823 (
            .O(N__38952),
            .I(N__38916));
    LocalMux I__6822 (
            .O(N__38947),
            .I(N__38913));
    LocalMux I__6821 (
            .O(N__38944),
            .I(N__38910));
    Span4Mux_v I__6820 (
            .O(N__38941),
            .I(N__38905));
    LocalMux I__6819 (
            .O(N__38938),
            .I(N__38905));
    LocalMux I__6818 (
            .O(N__38935),
            .I(N__38902));
    InMux I__6817 (
            .O(N__38932),
            .I(N__38897));
    InMux I__6816 (
            .O(N__38931),
            .I(N__38897));
    Span12Mux_v I__6815 (
            .O(N__38928),
            .I(N__38894));
    InMux I__6814 (
            .O(N__38927),
            .I(N__38891));
    InMux I__6813 (
            .O(N__38926),
            .I(N__38888));
    InMux I__6812 (
            .O(N__38925),
            .I(N__38885));
    Span4Mux_h I__6811 (
            .O(N__38922),
            .I(N__38880));
    Span4Mux_h I__6810 (
            .O(N__38919),
            .I(N__38880));
    LocalMux I__6809 (
            .O(N__38916),
            .I(N__38875));
    Span4Mux_h I__6808 (
            .O(N__38913),
            .I(N__38875));
    Span4Mux_v I__6807 (
            .O(N__38910),
            .I(N__38870));
    Span4Mux_v I__6806 (
            .O(N__38905),
            .I(N__38870));
    Span12Mux_v I__6805 (
            .O(N__38902),
            .I(N__38865));
    LocalMux I__6804 (
            .O(N__38897),
            .I(N__38865));
    Odrv12 I__6803 (
            .O(N__38894),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__6802 (
            .O(N__38891),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__6801 (
            .O(N__38888),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__6800 (
            .O(N__38885),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__6799 (
            .O(N__38880),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__6798 (
            .O(N__38875),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__6797 (
            .O(N__38870),
            .I(FRAME_MATCHER_state_2));
    Odrv12 I__6796 (
            .O(N__38865),
            .I(FRAME_MATCHER_state_2));
    InMux I__6795 (
            .O(N__38848),
            .I(N__38845));
    LocalMux I__6794 (
            .O(N__38845),
            .I(N__38842));
    Span4Mux_v I__6793 (
            .O(N__38842),
            .I(N__38838));
    InMux I__6792 (
            .O(N__38841),
            .I(N__38834));
    Span4Mux_h I__6791 (
            .O(N__38838),
            .I(N__38831));
    InMux I__6790 (
            .O(N__38837),
            .I(N__38828));
    LocalMux I__6789 (
            .O(N__38834),
            .I(N__38825));
    Sp12to4 I__6788 (
            .O(N__38831),
            .I(N__38818));
    LocalMux I__6787 (
            .O(N__38828),
            .I(N__38818));
    Span12Mux_h I__6786 (
            .O(N__38825),
            .I(N__38818));
    Span12Mux_v I__6785 (
            .O(N__38818),
            .I(N__38815));
    Odrv12 I__6784 (
            .O(N__38815),
            .I(\c0.n15499 ));
    InMux I__6783 (
            .O(N__38812),
            .I(N__38809));
    LocalMux I__6782 (
            .O(N__38809),
            .I(\c0.n13_adj_3016 ));
    CascadeMux I__6781 (
            .O(N__38806),
            .I(N__38803));
    InMux I__6780 (
            .O(N__38803),
            .I(N__38799));
    InMux I__6779 (
            .O(N__38802),
            .I(N__38796));
    LocalMux I__6778 (
            .O(N__38799),
            .I(N__38793));
    LocalMux I__6777 (
            .O(N__38796),
            .I(N__38790));
    Span4Mux_v I__6776 (
            .O(N__38793),
            .I(N__38787));
    Span4Mux_h I__6775 (
            .O(N__38790),
            .I(N__38783));
    Span4Mux_v I__6774 (
            .O(N__38787),
            .I(N__38780));
    InMux I__6773 (
            .O(N__38786),
            .I(N__38777));
    Odrv4 I__6772 (
            .O(N__38783),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    Odrv4 I__6771 (
            .O(N__38780),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    LocalMux I__6770 (
            .O(N__38777),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    CascadeMux I__6769 (
            .O(N__38770),
            .I(\c0.n19111_cascade_ ));
    InMux I__6768 (
            .O(N__38767),
            .I(N__38764));
    LocalMux I__6767 (
            .O(N__38764),
            .I(N__38760));
    InMux I__6766 (
            .O(N__38763),
            .I(N__38757));
    Odrv12 I__6765 (
            .O(N__38760),
            .I(\c0.n19493 ));
    LocalMux I__6764 (
            .O(N__38757),
            .I(\c0.n19493 ));
    InMux I__6763 (
            .O(N__38752),
            .I(N__38748));
    InMux I__6762 (
            .O(N__38751),
            .I(N__38745));
    LocalMux I__6761 (
            .O(N__38748),
            .I(control_mode_4));
    LocalMux I__6760 (
            .O(N__38745),
            .I(control_mode_4));
    InMux I__6759 (
            .O(N__38740),
            .I(N__38737));
    LocalMux I__6758 (
            .O(N__38737),
            .I(N__38734));
    Span4Mux_v I__6757 (
            .O(N__38734),
            .I(N__38730));
    InMux I__6756 (
            .O(N__38733),
            .I(N__38727));
    Odrv4 I__6755 (
            .O(N__38730),
            .I(control_mode_3));
    LocalMux I__6754 (
            .O(N__38727),
            .I(control_mode_3));
    InMux I__6753 (
            .O(N__38722),
            .I(N__38719));
    LocalMux I__6752 (
            .O(N__38719),
            .I(N__38716));
    Sp12to4 I__6751 (
            .O(N__38716),
            .I(N__38712));
    InMux I__6750 (
            .O(N__38715),
            .I(N__38709));
    Odrv12 I__6749 (
            .O(N__38712),
            .I(control_mode_7));
    LocalMux I__6748 (
            .O(N__38709),
            .I(control_mode_7));
    CascadeMux I__6747 (
            .O(N__38704),
            .I(\c0.n9_cascade_ ));
    CascadeMux I__6746 (
            .O(N__38701),
            .I(\c0.n16_adj_3008_cascade_ ));
    InMux I__6745 (
            .O(N__38698),
            .I(N__38695));
    LocalMux I__6744 (
            .O(N__38695),
            .I(\c0.n9 ));
    CascadeMux I__6743 (
            .O(N__38692),
            .I(\c0.n19115_cascade_ ));
    CascadeMux I__6742 (
            .O(N__38689),
            .I(N__38685));
    InMux I__6741 (
            .O(N__38688),
            .I(N__38682));
    InMux I__6740 (
            .O(N__38685),
            .I(N__38679));
    LocalMux I__6739 (
            .O(N__38682),
            .I(\c0.data_in_frame_10_1 ));
    LocalMux I__6738 (
            .O(N__38679),
            .I(\c0.data_in_frame_10_1 ));
    InMux I__6737 (
            .O(N__38674),
            .I(N__38671));
    LocalMux I__6736 (
            .O(N__38671),
            .I(N__38666));
    InMux I__6735 (
            .O(N__38670),
            .I(N__38663));
    InMux I__6734 (
            .O(N__38669),
            .I(N__38660));
    Span4Mux_h I__6733 (
            .O(N__38666),
            .I(N__38657));
    LocalMux I__6732 (
            .O(N__38663),
            .I(N__38654));
    LocalMux I__6731 (
            .O(N__38660),
            .I(N__38651));
    Span4Mux_v I__6730 (
            .O(N__38657),
            .I(N__38648));
    Span12Mux_v I__6729 (
            .O(N__38654),
            .I(N__38643));
    Span12Mux_h I__6728 (
            .O(N__38651),
            .I(N__38643));
    Odrv4 I__6727 (
            .O(N__38648),
            .I(\c0.n63_adj_3146 ));
    Odrv12 I__6726 (
            .O(N__38643),
            .I(\c0.n63_adj_3146 ));
    CascadeMux I__6725 (
            .O(N__38638),
            .I(\c0.n20_adj_3437_cascade_ ));
    CascadeMux I__6724 (
            .O(N__38635),
            .I(n21222_cascade_));
    InMux I__6723 (
            .O(N__38632),
            .I(N__38628));
    InMux I__6722 (
            .O(N__38631),
            .I(N__38625));
    LocalMux I__6721 (
            .O(N__38628),
            .I(control_mode_6));
    LocalMux I__6720 (
            .O(N__38625),
            .I(control_mode_6));
    InMux I__6719 (
            .O(N__38620),
            .I(N__38616));
    InMux I__6718 (
            .O(N__38619),
            .I(N__38613));
    LocalMux I__6717 (
            .O(N__38616),
            .I(control_mode_2));
    LocalMux I__6716 (
            .O(N__38613),
            .I(control_mode_2));
    CascadeMux I__6715 (
            .O(N__38608),
            .I(N__38604));
    CascadeMux I__6714 (
            .O(N__38607),
            .I(N__38601));
    InMux I__6713 (
            .O(N__38604),
            .I(N__38593));
    InMux I__6712 (
            .O(N__38601),
            .I(N__38593));
    InMux I__6711 (
            .O(N__38600),
            .I(N__38593));
    LocalMux I__6710 (
            .O(N__38593),
            .I(\c0.data_in_frame_5_0 ));
    CascadeMux I__6709 (
            .O(N__38590),
            .I(N__38586));
    CascadeMux I__6708 (
            .O(N__38589),
            .I(N__38583));
    InMux I__6707 (
            .O(N__38586),
            .I(N__38578));
    InMux I__6706 (
            .O(N__38583),
            .I(N__38578));
    LocalMux I__6705 (
            .O(N__38578),
            .I(\c0.data_in_frame_9_7 ));
    InMux I__6704 (
            .O(N__38575),
            .I(N__38572));
    LocalMux I__6703 (
            .O(N__38572),
            .I(\c0.n38_adj_3328 ));
    CascadeMux I__6702 (
            .O(N__38569),
            .I(\c0.n21279_cascade_ ));
    CascadeMux I__6701 (
            .O(N__38566),
            .I(\c0.n21255_cascade_ ));
    InMux I__6700 (
            .O(N__38563),
            .I(N__38560));
    LocalMux I__6699 (
            .O(N__38560),
            .I(\c0.n37_adj_3332 ));
    CascadeMux I__6698 (
            .O(N__38557),
            .I(\c0.n63_adj_3417_cascade_ ));
    CascadeMux I__6697 (
            .O(N__38554),
            .I(\c0.n5_adj_3040_cascade_ ));
    InMux I__6696 (
            .O(N__38551),
            .I(N__38548));
    LocalMux I__6695 (
            .O(N__38548),
            .I(N__38545));
    Odrv4 I__6694 (
            .O(N__38545),
            .I(\c0.n30_adj_3264 ));
    InMux I__6693 (
            .O(N__38542),
            .I(N__38539));
    LocalMux I__6692 (
            .O(N__38539),
            .I(\c0.n26_adj_3107 ));
    CascadeMux I__6691 (
            .O(N__38536),
            .I(\c0.n21281_cascade_ ));
    InMux I__6690 (
            .O(N__38533),
            .I(N__38530));
    LocalMux I__6689 (
            .O(N__38530),
            .I(\c0.n108 ));
    CascadeMux I__6688 (
            .O(N__38527),
            .I(\c0.n108_cascade_ ));
    InMux I__6687 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__6686 (
            .O(N__38521),
            .I(N__38516));
    InMux I__6685 (
            .O(N__38520),
            .I(N__38510));
    InMux I__6684 (
            .O(N__38519),
            .I(N__38510));
    Span4Mux_h I__6683 (
            .O(N__38516),
            .I(N__38507));
    InMux I__6682 (
            .O(N__38515),
            .I(N__38504));
    LocalMux I__6681 (
            .O(N__38510),
            .I(N__38501));
    Odrv4 I__6680 (
            .O(N__38507),
            .I(\c0.n92_adj_3254 ));
    LocalMux I__6679 (
            .O(N__38504),
            .I(\c0.n92_adj_3254 ));
    Odrv4 I__6678 (
            .O(N__38501),
            .I(\c0.n92_adj_3254 ));
    InMux I__6677 (
            .O(N__38494),
            .I(N__38486));
    InMux I__6676 (
            .O(N__38493),
            .I(N__38486));
    InMux I__6675 (
            .O(N__38492),
            .I(N__38481));
    InMux I__6674 (
            .O(N__38491),
            .I(N__38481));
    LocalMux I__6673 (
            .O(N__38486),
            .I(data_in_1_2));
    LocalMux I__6672 (
            .O(N__38481),
            .I(data_in_1_2));
    InMux I__6671 (
            .O(N__38476),
            .I(N__38473));
    LocalMux I__6670 (
            .O(N__38473),
            .I(N__38470));
    Span4Mux_v I__6669 (
            .O(N__38470),
            .I(N__38466));
    InMux I__6668 (
            .O(N__38469),
            .I(N__38463));
    Odrv4 I__6667 (
            .O(N__38466),
            .I(\c0.n121 ));
    LocalMux I__6666 (
            .O(N__38463),
            .I(\c0.n121 ));
    InMux I__6665 (
            .O(N__38458),
            .I(N__38452));
    InMux I__6664 (
            .O(N__38457),
            .I(N__38452));
    LocalMux I__6663 (
            .O(N__38452),
            .I(\c0.n103 ));
    InMux I__6662 (
            .O(N__38449),
            .I(N__38446));
    LocalMux I__6661 (
            .O(N__38446),
            .I(\c0.n63_adj_3084 ));
    InMux I__6660 (
            .O(N__38443),
            .I(N__38440));
    LocalMux I__6659 (
            .O(N__38440),
            .I(\c0.n19_adj_3252 ));
    InMux I__6658 (
            .O(N__38437),
            .I(N__38431));
    InMux I__6657 (
            .O(N__38436),
            .I(N__38431));
    LocalMux I__6656 (
            .O(N__38431),
            .I(\c0.n21_adj_3253 ));
    CascadeMux I__6655 (
            .O(N__38428),
            .I(\c0.n19_adj_3252_cascade_ ));
    InMux I__6654 (
            .O(N__38425),
            .I(N__38419));
    InMux I__6653 (
            .O(N__38424),
            .I(N__38419));
    LocalMux I__6652 (
            .O(N__38419),
            .I(\c0.n63_adj_3083 ));
    InMux I__6651 (
            .O(N__38416),
            .I(N__38408));
    InMux I__6650 (
            .O(N__38415),
            .I(N__38408));
    InMux I__6649 (
            .O(N__38414),
            .I(N__38403));
    InMux I__6648 (
            .O(N__38413),
            .I(N__38403));
    LocalMux I__6647 (
            .O(N__38408),
            .I(\c0.n7804 ));
    LocalMux I__6646 (
            .O(N__38403),
            .I(\c0.n7804 ));
    InMux I__6645 (
            .O(N__38398),
            .I(N__38395));
    LocalMux I__6644 (
            .O(N__38395),
            .I(N__38392));
    Span12Mux_v I__6643 (
            .O(N__38392),
            .I(N__38389));
    Odrv12 I__6642 (
            .O(N__38389),
            .I(\c0.n11_adj_3093 ));
    CascadeMux I__6641 (
            .O(N__38386),
            .I(\c0.n15701_cascade_ ));
    CascadeMux I__6640 (
            .O(N__38383),
            .I(n11421_cascade_));
    InMux I__6639 (
            .O(N__38380),
            .I(N__38377));
    LocalMux I__6638 (
            .O(N__38377),
            .I(N__38374));
    Span4Mux_v I__6637 (
            .O(N__38374),
            .I(N__38370));
    InMux I__6636 (
            .O(N__38373),
            .I(N__38367));
    Odrv4 I__6635 (
            .O(N__38370),
            .I(\c0.n11422 ));
    LocalMux I__6634 (
            .O(N__38367),
            .I(\c0.n11422 ));
    InMux I__6633 (
            .O(N__38362),
            .I(N__38358));
    InMux I__6632 (
            .O(N__38361),
            .I(N__38355));
    LocalMux I__6631 (
            .O(N__38358),
            .I(N__38349));
    LocalMux I__6630 (
            .O(N__38355),
            .I(N__38349));
    InMux I__6629 (
            .O(N__38354),
            .I(N__38345));
    Span4Mux_v I__6628 (
            .O(N__38349),
            .I(N__38342));
    InMux I__6627 (
            .O(N__38348),
            .I(N__38339));
    LocalMux I__6626 (
            .O(N__38345),
            .I(N__38336));
    Span4Mux_h I__6625 (
            .O(N__38342),
            .I(N__38331));
    LocalMux I__6624 (
            .O(N__38339),
            .I(N__38331));
    Odrv4 I__6623 (
            .O(N__38336),
            .I(\c0.n3632 ));
    Odrv4 I__6622 (
            .O(N__38331),
            .I(\c0.n3632 ));
    InMux I__6621 (
            .O(N__38326),
            .I(N__38322));
    InMux I__6620 (
            .O(N__38325),
            .I(N__38318));
    LocalMux I__6619 (
            .O(N__38322),
            .I(N__38314));
    InMux I__6618 (
            .O(N__38321),
            .I(N__38310));
    LocalMux I__6617 (
            .O(N__38318),
            .I(N__38307));
    InMux I__6616 (
            .O(N__38317),
            .I(N__38304));
    Span4Mux_v I__6615 (
            .O(N__38314),
            .I(N__38301));
    InMux I__6614 (
            .O(N__38313),
            .I(N__38298));
    LocalMux I__6613 (
            .O(N__38310),
            .I(N__38293));
    Span4Mux_v I__6612 (
            .O(N__38307),
            .I(N__38293));
    LocalMux I__6611 (
            .O(N__38304),
            .I(\c0.n9389 ));
    Odrv4 I__6610 (
            .O(N__38301),
            .I(\c0.n9389 ));
    LocalMux I__6609 (
            .O(N__38298),
            .I(\c0.n9389 ));
    Odrv4 I__6608 (
            .O(N__38293),
            .I(\c0.n9389 ));
    InMux I__6607 (
            .O(N__38284),
            .I(N__38281));
    LocalMux I__6606 (
            .O(N__38281),
            .I(N__38278));
    Span4Mux_h I__6605 (
            .O(N__38278),
            .I(N__38274));
    InMux I__6604 (
            .O(N__38277),
            .I(N__38271));
    Odrv4 I__6603 (
            .O(N__38274),
            .I(\c0.n3 ));
    LocalMux I__6602 (
            .O(N__38271),
            .I(\c0.n3 ));
    InMux I__6601 (
            .O(N__38266),
            .I(N__38262));
    InMux I__6600 (
            .O(N__38265),
            .I(N__38259));
    LocalMux I__6599 (
            .O(N__38262),
            .I(N__38255));
    LocalMux I__6598 (
            .O(N__38259),
            .I(N__38252));
    InMux I__6597 (
            .O(N__38258),
            .I(N__38249));
    Span4Mux_v I__6596 (
            .O(N__38255),
            .I(N__38238));
    Span4Mux_h I__6595 (
            .O(N__38252),
            .I(N__38238));
    LocalMux I__6594 (
            .O(N__38249),
            .I(N__38238));
    InMux I__6593 (
            .O(N__38248),
            .I(N__38235));
    InMux I__6592 (
            .O(N__38247),
            .I(N__38230));
    InMux I__6591 (
            .O(N__38246),
            .I(N__38230));
    InMux I__6590 (
            .O(N__38245),
            .I(N__38227));
    Span4Mux_h I__6589 (
            .O(N__38238),
            .I(N__38224));
    LocalMux I__6588 (
            .O(N__38235),
            .I(N__38221));
    LocalMux I__6587 (
            .O(N__38230),
            .I(\c0.n11427 ));
    LocalMux I__6586 (
            .O(N__38227),
            .I(\c0.n11427 ));
    Odrv4 I__6585 (
            .O(N__38224),
            .I(\c0.n11427 ));
    Odrv12 I__6584 (
            .O(N__38221),
            .I(\c0.n11427 ));
    InMux I__6583 (
            .O(N__38212),
            .I(N__38208));
    InMux I__6582 (
            .O(N__38211),
            .I(N__38205));
    LocalMux I__6581 (
            .O(N__38208),
            .I(\c0.n15874 ));
    LocalMux I__6580 (
            .O(N__38205),
            .I(\c0.n15874 ));
    InMux I__6579 (
            .O(N__38200),
            .I(N__38197));
    LocalMux I__6578 (
            .O(N__38197),
            .I(n12917));
    InMux I__6577 (
            .O(N__38194),
            .I(N__38190));
    InMux I__6576 (
            .O(N__38193),
            .I(N__38187));
    LocalMux I__6575 (
            .O(N__38190),
            .I(N__38181));
    LocalMux I__6574 (
            .O(N__38187),
            .I(N__38181));
    InMux I__6573 (
            .O(N__38186),
            .I(N__38178));
    Span4Mux_h I__6572 (
            .O(N__38181),
            .I(N__38175));
    LocalMux I__6571 (
            .O(N__38178),
            .I(\c0.n11440 ));
    Odrv4 I__6570 (
            .O(N__38175),
            .I(\c0.n11440 ));
    CascadeMux I__6569 (
            .O(N__38170),
            .I(\c0.n11317_cascade_ ));
    CascadeMux I__6568 (
            .O(N__38167),
            .I(N__38164));
    InMux I__6567 (
            .O(N__38164),
            .I(N__38161));
    LocalMux I__6566 (
            .O(N__38161),
            .I(N__38157));
    InMux I__6565 (
            .O(N__38160),
            .I(N__38154));
    Span4Mux_v I__6564 (
            .O(N__38157),
            .I(N__38150));
    LocalMux I__6563 (
            .O(N__38154),
            .I(N__38147));
    InMux I__6562 (
            .O(N__38153),
            .I(N__38144));
    Span4Mux_v I__6561 (
            .O(N__38150),
            .I(N__38141));
    Span4Mux_h I__6560 (
            .O(N__38147),
            .I(N__38136));
    LocalMux I__6559 (
            .O(N__38144),
            .I(N__38136));
    Span4Mux_v I__6558 (
            .O(N__38141),
            .I(N__38131));
    Sp12to4 I__6557 (
            .O(N__38136),
            .I(N__38128));
    InMux I__6556 (
            .O(N__38135),
            .I(N__38125));
    InMux I__6555 (
            .O(N__38134),
            .I(N__38122));
    Span4Mux_v I__6554 (
            .O(N__38131),
            .I(N__38119));
    Span12Mux_v I__6553 (
            .O(N__38128),
            .I(N__38116));
    LocalMux I__6552 (
            .O(N__38125),
            .I(\c0.FRAME_MATCHER_i_31 ));
    LocalMux I__6551 (
            .O(N__38122),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__6550 (
            .O(N__38119),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv12 I__6549 (
            .O(N__38116),
            .I(\c0.FRAME_MATCHER_i_31 ));
    InMux I__6548 (
            .O(N__38107),
            .I(N__38101));
    InMux I__6547 (
            .O(N__38106),
            .I(N__38098));
    InMux I__6546 (
            .O(N__38105),
            .I(N__38095));
    InMux I__6545 (
            .O(N__38104),
            .I(N__38092));
    LocalMux I__6544 (
            .O(N__38101),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__6543 (
            .O(N__38098),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__6542 (
            .O(N__38095),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__6541 (
            .O(N__38092),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__6540 (
            .O(N__38083),
            .I(N__38077));
    InMux I__6539 (
            .O(N__38082),
            .I(N__38074));
    InMux I__6538 (
            .O(N__38081),
            .I(N__38071));
    InMux I__6537 (
            .O(N__38080),
            .I(N__38068));
    LocalMux I__6536 (
            .O(N__38077),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__6535 (
            .O(N__38074),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__6534 (
            .O(N__38071),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__6533 (
            .O(N__38068),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__6532 (
            .O(N__38059),
            .I(N__38056));
    LocalMux I__6531 (
            .O(N__38056),
            .I(N__38053));
    Odrv4 I__6530 (
            .O(N__38053),
            .I(\c0.rx.n21267 ));
    InMux I__6529 (
            .O(N__38050),
            .I(N__38047));
    LocalMux I__6528 (
            .O(N__38047),
            .I(N__38042));
    InMux I__6527 (
            .O(N__38046),
            .I(N__38039));
    InMux I__6526 (
            .O(N__38045),
            .I(N__38036));
    Span4Mux_h I__6525 (
            .O(N__38042),
            .I(N__38033));
    LocalMux I__6524 (
            .O(N__38039),
            .I(\c0.FRAME_MATCHER_i_18 ));
    LocalMux I__6523 (
            .O(N__38036),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__6522 (
            .O(N__38033),
            .I(\c0.FRAME_MATCHER_i_18 ));
    CascadeMux I__6521 (
            .O(N__38026),
            .I(N__38023));
    InMux I__6520 (
            .O(N__38023),
            .I(N__38020));
    LocalMux I__6519 (
            .O(N__38020),
            .I(N__38015));
    InMux I__6518 (
            .O(N__38019),
            .I(N__38012));
    InMux I__6517 (
            .O(N__38018),
            .I(N__38009));
    Span4Mux_h I__6516 (
            .O(N__38015),
            .I(N__38006));
    LocalMux I__6515 (
            .O(N__38012),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__6514 (
            .O(N__38009),
            .I(\c0.FRAME_MATCHER_i_23 ));
    Odrv4 I__6513 (
            .O(N__38006),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__6512 (
            .O(N__37999),
            .I(N__37996));
    LocalMux I__6511 (
            .O(N__37996),
            .I(N__37993));
    Span4Mux_v I__6510 (
            .O(N__37993),
            .I(N__37989));
    InMux I__6509 (
            .O(N__37992),
            .I(N__37986));
    Span4Mux_v I__6508 (
            .O(N__37989),
            .I(N__37982));
    LocalMux I__6507 (
            .O(N__37986),
            .I(N__37979));
    InMux I__6506 (
            .O(N__37985),
            .I(N__37976));
    Span4Mux_v I__6505 (
            .O(N__37982),
            .I(N__37973));
    Odrv4 I__6504 (
            .O(N__37979),
            .I(\c0.FRAME_MATCHER_i_29 ));
    LocalMux I__6503 (
            .O(N__37976),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv4 I__6502 (
            .O(N__37973),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__6501 (
            .O(N__37966),
            .I(N__37963));
    LocalMux I__6500 (
            .O(N__37963),
            .I(\c0.n42_adj_3256 ));
    InMux I__6499 (
            .O(N__37960),
            .I(N__37956));
    InMux I__6498 (
            .O(N__37959),
            .I(N__37953));
    LocalMux I__6497 (
            .O(N__37956),
            .I(N__37950));
    LocalMux I__6496 (
            .O(N__37953),
            .I(N__37947));
    Odrv4 I__6495 (
            .O(N__37950),
            .I(\c0.n1_adj_3002 ));
    Odrv4 I__6494 (
            .O(N__37947),
            .I(\c0.n1_adj_3002 ));
    InMux I__6493 (
            .O(N__37942),
            .I(N__37939));
    LocalMux I__6492 (
            .O(N__37939),
            .I(N__37936));
    Odrv12 I__6491 (
            .O(N__37936),
            .I(\c0.n21053 ));
    CascadeMux I__6490 (
            .O(N__37933),
            .I(\c0.rx.n35_cascade_ ));
    CascadeMux I__6489 (
            .O(N__37930),
            .I(N__37924));
    CascadeMux I__6488 (
            .O(N__37929),
            .I(N__37917));
    InMux I__6487 (
            .O(N__37928),
            .I(N__37914));
    InMux I__6486 (
            .O(N__37927),
            .I(N__37907));
    InMux I__6485 (
            .O(N__37924),
            .I(N__37907));
    InMux I__6484 (
            .O(N__37923),
            .I(N__37900));
    InMux I__6483 (
            .O(N__37922),
            .I(N__37900));
    InMux I__6482 (
            .O(N__37921),
            .I(N__37900));
    InMux I__6481 (
            .O(N__37920),
            .I(N__37895));
    InMux I__6480 (
            .O(N__37917),
            .I(N__37895));
    LocalMux I__6479 (
            .O(N__37914),
            .I(N__37892));
    InMux I__6478 (
            .O(N__37913),
            .I(N__37887));
    InMux I__6477 (
            .O(N__37912),
            .I(N__37887));
    LocalMux I__6476 (
            .O(N__37907),
            .I(N__37884));
    LocalMux I__6475 (
            .O(N__37900),
            .I(r_SM_Main_0));
    LocalMux I__6474 (
            .O(N__37895),
            .I(r_SM_Main_0));
    Odrv4 I__6473 (
            .O(N__37892),
            .I(r_SM_Main_0));
    LocalMux I__6472 (
            .O(N__37887),
            .I(r_SM_Main_0));
    Odrv4 I__6471 (
            .O(N__37884),
            .I(r_SM_Main_0));
    CascadeMux I__6470 (
            .O(N__37873),
            .I(\c0.rx.n12_cascade_ ));
    InMux I__6469 (
            .O(N__37870),
            .I(N__37867));
    LocalMux I__6468 (
            .O(N__37867),
            .I(N__37864));
    Span4Mux_h I__6467 (
            .O(N__37864),
            .I(N__37859));
    InMux I__6466 (
            .O(N__37863),
            .I(N__37854));
    InMux I__6465 (
            .O(N__37862),
            .I(N__37846));
    Span4Mux_v I__6464 (
            .O(N__37859),
            .I(N__37843));
    InMux I__6463 (
            .O(N__37858),
            .I(N__37838));
    InMux I__6462 (
            .O(N__37857),
            .I(N__37838));
    LocalMux I__6461 (
            .O(N__37854),
            .I(N__37835));
    InMux I__6460 (
            .O(N__37853),
            .I(N__37828));
    InMux I__6459 (
            .O(N__37852),
            .I(N__37828));
    InMux I__6458 (
            .O(N__37851),
            .I(N__37828));
    InMux I__6457 (
            .O(N__37850),
            .I(N__37823));
    InMux I__6456 (
            .O(N__37849),
            .I(N__37823));
    LocalMux I__6455 (
            .O(N__37846),
            .I(r_SM_Main_1));
    Odrv4 I__6454 (
            .O(N__37843),
            .I(r_SM_Main_1));
    LocalMux I__6453 (
            .O(N__37838),
            .I(r_SM_Main_1));
    Odrv4 I__6452 (
            .O(N__37835),
            .I(r_SM_Main_1));
    LocalMux I__6451 (
            .O(N__37828),
            .I(r_SM_Main_1));
    LocalMux I__6450 (
            .O(N__37823),
            .I(r_SM_Main_1));
    InMux I__6449 (
            .O(N__37810),
            .I(N__37807));
    LocalMux I__6448 (
            .O(N__37807),
            .I(N__37802));
    InMux I__6447 (
            .O(N__37806),
            .I(N__37791));
    InMux I__6446 (
            .O(N__37805),
            .I(N__37791));
    Sp12to4 I__6445 (
            .O(N__37802),
            .I(N__37788));
    InMux I__6444 (
            .O(N__37801),
            .I(N__37785));
    InMux I__6443 (
            .O(N__37800),
            .I(N__37780));
    InMux I__6442 (
            .O(N__37799),
            .I(N__37780));
    InMux I__6441 (
            .O(N__37798),
            .I(N__37777));
    InMux I__6440 (
            .O(N__37797),
            .I(N__37772));
    InMux I__6439 (
            .O(N__37796),
            .I(N__37772));
    LocalMux I__6438 (
            .O(N__37791),
            .I(N__37769));
    Odrv12 I__6437 (
            .O(N__37788),
            .I(r_SM_Main_2));
    LocalMux I__6436 (
            .O(N__37785),
            .I(r_SM_Main_2));
    LocalMux I__6435 (
            .O(N__37780),
            .I(r_SM_Main_2));
    LocalMux I__6434 (
            .O(N__37777),
            .I(r_SM_Main_2));
    LocalMux I__6433 (
            .O(N__37772),
            .I(r_SM_Main_2));
    Odrv4 I__6432 (
            .O(N__37769),
            .I(r_SM_Main_2));
    CascadeMux I__6431 (
            .O(N__37756),
            .I(\c0.rx.n21406_cascade_ ));
    CascadeMux I__6430 (
            .O(N__37753),
            .I(N__37750));
    InMux I__6429 (
            .O(N__37750),
            .I(N__37745));
    InMux I__6428 (
            .O(N__37749),
            .I(N__37741));
    InMux I__6427 (
            .O(N__37748),
            .I(N__37738));
    LocalMux I__6426 (
            .O(N__37745),
            .I(N__37735));
    InMux I__6425 (
            .O(N__37744),
            .I(N__37732));
    LocalMux I__6424 (
            .O(N__37741),
            .I(r_SM_Main_2_N_2473_2));
    LocalMux I__6423 (
            .O(N__37738),
            .I(r_SM_Main_2_N_2473_2));
    Odrv4 I__6422 (
            .O(N__37735),
            .I(r_SM_Main_2_N_2473_2));
    LocalMux I__6421 (
            .O(N__37732),
            .I(r_SM_Main_2_N_2473_2));
    InMux I__6420 (
            .O(N__37723),
            .I(N__37719));
    InMux I__6419 (
            .O(N__37722),
            .I(N__37716));
    LocalMux I__6418 (
            .O(N__37719),
            .I(N__37710));
    LocalMux I__6417 (
            .O(N__37716),
            .I(N__37707));
    InMux I__6416 (
            .O(N__37715),
            .I(N__37704));
    InMux I__6415 (
            .O(N__37714),
            .I(N__37699));
    InMux I__6414 (
            .O(N__37713),
            .I(N__37699));
    Sp12to4 I__6413 (
            .O(N__37710),
            .I(N__37690));
    Sp12to4 I__6412 (
            .O(N__37707),
            .I(N__37690));
    LocalMux I__6411 (
            .O(N__37704),
            .I(N__37690));
    LocalMux I__6410 (
            .O(N__37699),
            .I(N__37690));
    Odrv12 I__6409 (
            .O(N__37690),
            .I(\c0.rx.r_Clock_Count_6 ));
    InMux I__6408 (
            .O(N__37687),
            .I(N__37684));
    LocalMux I__6407 (
            .O(N__37684),
            .I(N__37676));
    InMux I__6406 (
            .O(N__37683),
            .I(N__37673));
    InMux I__6405 (
            .O(N__37682),
            .I(N__37670));
    InMux I__6404 (
            .O(N__37681),
            .I(N__37663));
    InMux I__6403 (
            .O(N__37680),
            .I(N__37663));
    InMux I__6402 (
            .O(N__37679),
            .I(N__37663));
    Odrv4 I__6401 (
            .O(N__37676),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__6400 (
            .O(N__37673),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__6399 (
            .O(N__37670),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__6398 (
            .O(N__37663),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__6397 (
            .O(N__37654),
            .I(N__37649));
    CascadeMux I__6396 (
            .O(N__37653),
            .I(N__37644));
    InMux I__6395 (
            .O(N__37652),
            .I(N__37641));
    LocalMux I__6394 (
            .O(N__37649),
            .I(N__37638));
    InMux I__6393 (
            .O(N__37648),
            .I(N__37633));
    InMux I__6392 (
            .O(N__37647),
            .I(N__37633));
    InMux I__6391 (
            .O(N__37644),
            .I(N__37630));
    LocalMux I__6390 (
            .O(N__37641),
            .I(\c0.rx.r_Clock_Count_0 ));
    Odrv4 I__6389 (
            .O(N__37638),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__6388 (
            .O(N__37633),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__6387 (
            .O(N__37630),
            .I(\c0.rx.r_Clock_Count_0 ));
    InMux I__6386 (
            .O(N__37621),
            .I(N__37618));
    LocalMux I__6385 (
            .O(N__37618),
            .I(N__37614));
    InMux I__6384 (
            .O(N__37617),
            .I(N__37611));
    Span4Mux_h I__6383 (
            .O(N__37614),
            .I(N__37603));
    LocalMux I__6382 (
            .O(N__37611),
            .I(N__37603));
    InMux I__6381 (
            .O(N__37610),
            .I(N__37600));
    InMux I__6380 (
            .O(N__37609),
            .I(N__37595));
    InMux I__6379 (
            .O(N__37608),
            .I(N__37595));
    Sp12to4 I__6378 (
            .O(N__37603),
            .I(N__37588));
    LocalMux I__6377 (
            .O(N__37600),
            .I(N__37588));
    LocalMux I__6376 (
            .O(N__37595),
            .I(N__37588));
    Odrv12 I__6375 (
            .O(N__37588),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__6374 (
            .O(N__37585),
            .I(N__37582));
    LocalMux I__6373 (
            .O(N__37582),
            .I(\c0.rx.n8 ));
    InMux I__6372 (
            .O(N__37579),
            .I(N__37576));
    LocalMux I__6371 (
            .O(N__37576),
            .I(n12914));
    CascadeMux I__6370 (
            .O(N__37573),
            .I(\c0.rx.n15906_cascade_ ));
    InMux I__6369 (
            .O(N__37570),
            .I(N__37567));
    LocalMux I__6368 (
            .O(N__37567),
            .I(\c0.rx.n20851 ));
    CascadeMux I__6367 (
            .O(N__37564),
            .I(N__37561));
    InMux I__6366 (
            .O(N__37561),
            .I(N__37558));
    LocalMux I__6365 (
            .O(N__37558),
            .I(\c0.rx.n32 ));
    SRMux I__6364 (
            .O(N__37555),
            .I(N__37552));
    LocalMux I__6363 (
            .O(N__37552),
            .I(\c0.rx.n20964 ));
    InMux I__6362 (
            .O(N__37549),
            .I(N__37543));
    InMux I__6361 (
            .O(N__37548),
            .I(N__37543));
    LocalMux I__6360 (
            .O(N__37543),
            .I(\c0.rx.n15906 ));
    CascadeMux I__6359 (
            .O(N__37540),
            .I(r_SM_Main_2_N_2473_2_cascade_));
    InMux I__6358 (
            .O(N__37537),
            .I(N__37534));
    LocalMux I__6357 (
            .O(N__37534),
            .I(\c0.rx.n15926 ));
    InMux I__6356 (
            .O(N__37531),
            .I(N__37528));
    LocalMux I__6355 (
            .O(N__37528),
            .I(n9));
    InMux I__6354 (
            .O(N__37525),
            .I(N__37519));
    InMux I__6353 (
            .O(N__37524),
            .I(N__37516));
    InMux I__6352 (
            .O(N__37523),
            .I(N__37511));
    InMux I__6351 (
            .O(N__37522),
            .I(N__37511));
    LocalMux I__6350 (
            .O(N__37519),
            .I(N__37506));
    LocalMux I__6349 (
            .O(N__37516),
            .I(N__37506));
    LocalMux I__6348 (
            .O(N__37511),
            .I(N__37503));
    Odrv12 I__6347 (
            .O(N__37506),
            .I(\c0.n9755 ));
    Odrv4 I__6346 (
            .O(N__37503),
            .I(\c0.n9755 ));
    CascadeMux I__6345 (
            .O(N__37498),
            .I(N__37495));
    InMux I__6344 (
            .O(N__37495),
            .I(N__37492));
    LocalMux I__6343 (
            .O(N__37492),
            .I(N__37489));
    Span4Mux_h I__6342 (
            .O(N__37489),
            .I(N__37485));
    InMux I__6341 (
            .O(N__37488),
            .I(N__37482));
    Span4Mux_v I__6340 (
            .O(N__37485),
            .I(N__37479));
    LocalMux I__6339 (
            .O(N__37482),
            .I(data_out_frame_28_5));
    Odrv4 I__6338 (
            .O(N__37479),
            .I(data_out_frame_28_5));
    InMux I__6337 (
            .O(N__37474),
            .I(N__37471));
    LocalMux I__6336 (
            .O(N__37471),
            .I(\c0.n21308 ));
    InMux I__6335 (
            .O(N__37468),
            .I(N__37455));
    InMux I__6334 (
            .O(N__37467),
            .I(N__37455));
    InMux I__6333 (
            .O(N__37466),
            .I(N__37452));
    CascadeMux I__6332 (
            .O(N__37465),
            .I(N__37447));
    InMux I__6331 (
            .O(N__37464),
            .I(N__37444));
    InMux I__6330 (
            .O(N__37463),
            .I(N__37434));
    InMux I__6329 (
            .O(N__37462),
            .I(N__37434));
    InMux I__6328 (
            .O(N__37461),
            .I(N__37434));
    InMux I__6327 (
            .O(N__37460),
            .I(N__37434));
    LocalMux I__6326 (
            .O(N__37455),
            .I(N__37429));
    LocalMux I__6325 (
            .O(N__37452),
            .I(N__37429));
    CascadeMux I__6324 (
            .O(N__37451),
            .I(N__37425));
    InMux I__6323 (
            .O(N__37450),
            .I(N__37419));
    InMux I__6322 (
            .O(N__37447),
            .I(N__37416));
    LocalMux I__6321 (
            .O(N__37444),
            .I(N__37413));
    CascadeMux I__6320 (
            .O(N__37443),
            .I(N__37409));
    LocalMux I__6319 (
            .O(N__37434),
            .I(N__37405));
    Sp12to4 I__6318 (
            .O(N__37429),
            .I(N__37402));
    InMux I__6317 (
            .O(N__37428),
            .I(N__37391));
    InMux I__6316 (
            .O(N__37425),
            .I(N__37391));
    InMux I__6315 (
            .O(N__37424),
            .I(N__37391));
    InMux I__6314 (
            .O(N__37423),
            .I(N__37391));
    InMux I__6313 (
            .O(N__37422),
            .I(N__37391));
    LocalMux I__6312 (
            .O(N__37419),
            .I(N__37388));
    LocalMux I__6311 (
            .O(N__37416),
            .I(N__37385));
    Span4Mux_v I__6310 (
            .O(N__37413),
            .I(N__37382));
    InMux I__6309 (
            .O(N__37412),
            .I(N__37379));
    InMux I__6308 (
            .O(N__37409),
            .I(N__37376));
    InMux I__6307 (
            .O(N__37408),
            .I(N__37373));
    Span4Mux_h I__6306 (
            .O(N__37405),
            .I(N__37370));
    Span12Mux_v I__6305 (
            .O(N__37402),
            .I(N__37367));
    LocalMux I__6304 (
            .O(N__37391),
            .I(N__37356));
    Span4Mux_v I__6303 (
            .O(N__37388),
            .I(N__37356));
    Span4Mux_h I__6302 (
            .O(N__37385),
            .I(N__37356));
    Span4Mux_h I__6301 (
            .O(N__37382),
            .I(N__37356));
    LocalMux I__6300 (
            .O(N__37379),
            .I(N__37356));
    LocalMux I__6299 (
            .O(N__37376),
            .I(byte_transmit_counter_4));
    LocalMux I__6298 (
            .O(N__37373),
            .I(byte_transmit_counter_4));
    Odrv4 I__6297 (
            .O(N__37370),
            .I(byte_transmit_counter_4));
    Odrv12 I__6296 (
            .O(N__37367),
            .I(byte_transmit_counter_4));
    Odrv4 I__6295 (
            .O(N__37356),
            .I(byte_transmit_counter_4));
    InMux I__6294 (
            .O(N__37345),
            .I(N__37337));
    InMux I__6293 (
            .O(N__37344),
            .I(N__37330));
    InMux I__6292 (
            .O(N__37343),
            .I(N__37330));
    InMux I__6291 (
            .O(N__37342),
            .I(N__37323));
    InMux I__6290 (
            .O(N__37341),
            .I(N__37323));
    InMux I__6289 (
            .O(N__37340),
            .I(N__37323));
    LocalMux I__6288 (
            .O(N__37337),
            .I(N__37320));
    InMux I__6287 (
            .O(N__37336),
            .I(N__37317));
    CascadeMux I__6286 (
            .O(N__37335),
            .I(N__37313));
    LocalMux I__6285 (
            .O(N__37330),
            .I(N__37308));
    LocalMux I__6284 (
            .O(N__37323),
            .I(N__37305));
    Span4Mux_h I__6283 (
            .O(N__37320),
            .I(N__37302));
    LocalMux I__6282 (
            .O(N__37317),
            .I(N__37298));
    InMux I__6281 (
            .O(N__37316),
            .I(N__37295));
    InMux I__6280 (
            .O(N__37313),
            .I(N__37292));
    InMux I__6279 (
            .O(N__37312),
            .I(N__37289));
    InMux I__6278 (
            .O(N__37311),
            .I(N__37286));
    Span4Mux_v I__6277 (
            .O(N__37308),
            .I(N__37283));
    Span4Mux_h I__6276 (
            .O(N__37305),
            .I(N__37278));
    Span4Mux_v I__6275 (
            .O(N__37302),
            .I(N__37278));
    InMux I__6274 (
            .O(N__37301),
            .I(N__37275));
    Span4Mux_v I__6273 (
            .O(N__37298),
            .I(N__37268));
    LocalMux I__6272 (
            .O(N__37295),
            .I(N__37268));
    LocalMux I__6271 (
            .O(N__37292),
            .I(N__37268));
    LocalMux I__6270 (
            .O(N__37289),
            .I(byte_transmit_counter_3));
    LocalMux I__6269 (
            .O(N__37286),
            .I(byte_transmit_counter_3));
    Odrv4 I__6268 (
            .O(N__37283),
            .I(byte_transmit_counter_3));
    Odrv4 I__6267 (
            .O(N__37278),
            .I(byte_transmit_counter_3));
    LocalMux I__6266 (
            .O(N__37275),
            .I(byte_transmit_counter_3));
    Odrv4 I__6265 (
            .O(N__37268),
            .I(byte_transmit_counter_3));
    CascadeMux I__6264 (
            .O(N__37255),
            .I(\c0.n21310_cascade_ ));
    InMux I__6263 (
            .O(N__37252),
            .I(N__37249));
    LocalMux I__6262 (
            .O(N__37249),
            .I(N__37246));
    Odrv12 I__6261 (
            .O(N__37246),
            .I(\c0.n21568 ));
    InMux I__6260 (
            .O(N__37243),
            .I(N__37240));
    LocalMux I__6259 (
            .O(N__37240),
            .I(N__37237));
    Span4Mux_v I__6258 (
            .O(N__37237),
            .I(N__37234));
    Odrv4 I__6257 (
            .O(N__37234),
            .I(n9_adj_3590));
    InMux I__6256 (
            .O(N__37231),
            .I(N__37228));
    LocalMux I__6255 (
            .O(N__37228),
            .I(N__37225));
    Span4Mux_v I__6254 (
            .O(N__37225),
            .I(N__37222));
    Odrv4 I__6253 (
            .O(N__37222),
            .I(\c0.rx.n11302 ));
    CascadeMux I__6252 (
            .O(N__37219),
            .I(\c0.rx.n11302_cascade_ ));
    InMux I__6251 (
            .O(N__37216),
            .I(N__37213));
    LocalMux I__6250 (
            .O(N__37213),
            .I(N__37208));
    CascadeMux I__6249 (
            .O(N__37212),
            .I(N__37205));
    InMux I__6248 (
            .O(N__37211),
            .I(N__37202));
    Span4Mux_h I__6247 (
            .O(N__37208),
            .I(N__37199));
    InMux I__6246 (
            .O(N__37205),
            .I(N__37196));
    LocalMux I__6245 (
            .O(N__37202),
            .I(N__37191));
    Span4Mux_v I__6244 (
            .O(N__37199),
            .I(N__37191));
    LocalMux I__6243 (
            .O(N__37196),
            .I(N__37188));
    Odrv4 I__6242 (
            .O(N__37191),
            .I(encoder1_position_0));
    Odrv12 I__6241 (
            .O(N__37188),
            .I(encoder1_position_0));
    InMux I__6240 (
            .O(N__37183),
            .I(N__37179));
    InMux I__6239 (
            .O(N__37182),
            .I(N__37176));
    LocalMux I__6238 (
            .O(N__37179),
            .I(N__37173));
    LocalMux I__6237 (
            .O(N__37176),
            .I(data_out_frame_13_0));
    Odrv12 I__6236 (
            .O(N__37173),
            .I(data_out_frame_13_0));
    CascadeMux I__6235 (
            .O(N__37168),
            .I(\c0.rx.n21451_cascade_ ));
    InMux I__6234 (
            .O(N__37165),
            .I(N__37162));
    LocalMux I__6233 (
            .O(N__37162),
            .I(N__37159));
    Span4Mux_v I__6232 (
            .O(N__37159),
            .I(N__37156));
    Odrv4 I__6231 (
            .O(N__37156),
            .I(n12920));
    InMux I__6230 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__6229 (
            .O(N__37150),
            .I(N__37146));
    InMux I__6228 (
            .O(N__37149),
            .I(N__37143));
    Span12Mux_h I__6227 (
            .O(N__37146),
            .I(N__37138));
    LocalMux I__6226 (
            .O(N__37143),
            .I(N__37138));
    Odrv12 I__6225 (
            .O(N__37138),
            .I(\c0.n70 ));
    InMux I__6224 (
            .O(N__37135),
            .I(N__37132));
    LocalMux I__6223 (
            .O(N__37132),
            .I(N__37129));
    Span4Mux_v I__6222 (
            .O(N__37129),
            .I(N__37125));
    InMux I__6221 (
            .O(N__37128),
            .I(N__37122));
    Span4Mux_v I__6220 (
            .O(N__37125),
            .I(N__37119));
    LocalMux I__6219 (
            .O(N__37122),
            .I(N__37116));
    Odrv4 I__6218 (
            .O(N__37119),
            .I(\c0.n15850 ));
    Odrv4 I__6217 (
            .O(N__37116),
            .I(\c0.n15850 ));
    CascadeMux I__6216 (
            .O(N__37111),
            .I(N__37108));
    InMux I__6215 (
            .O(N__37108),
            .I(N__37105));
    LocalMux I__6214 (
            .O(N__37105),
            .I(N__37102));
    Span4Mux_v I__6213 (
            .O(N__37102),
            .I(N__37099));
    Span4Mux_h I__6212 (
            .O(N__37099),
            .I(N__37096));
    Odrv4 I__6211 (
            .O(N__37096),
            .I(\c0.n21231 ));
    CascadeMux I__6210 (
            .O(N__37093),
            .I(N__37088));
    CascadeMux I__6209 (
            .O(N__37092),
            .I(N__37085));
    InMux I__6208 (
            .O(N__37091),
            .I(N__37082));
    InMux I__6207 (
            .O(N__37088),
            .I(N__37077));
    InMux I__6206 (
            .O(N__37085),
            .I(N__37077));
    LocalMux I__6205 (
            .O(N__37082),
            .I(N__37074));
    LocalMux I__6204 (
            .O(N__37077),
            .I(N__37071));
    Span4Mux_h I__6203 (
            .O(N__37074),
            .I(N__37068));
    Span4Mux_h I__6202 (
            .O(N__37071),
            .I(N__37065));
    Odrv4 I__6201 (
            .O(N__37068),
            .I(\c0.n12254 ));
    Odrv4 I__6200 (
            .O(N__37065),
            .I(\c0.n12254 ));
    CascadeMux I__6199 (
            .O(N__37060),
            .I(N__37056));
    InMux I__6198 (
            .O(N__37059),
            .I(N__37053));
    InMux I__6197 (
            .O(N__37056),
            .I(N__37050));
    LocalMux I__6196 (
            .O(N__37053),
            .I(N__37047));
    LocalMux I__6195 (
            .O(N__37050),
            .I(N__37043));
    Sp12to4 I__6194 (
            .O(N__37047),
            .I(N__37040));
    InMux I__6193 (
            .O(N__37046),
            .I(N__37037));
    Span4Mux_h I__6192 (
            .O(N__37043),
            .I(N__37034));
    Odrv12 I__6191 (
            .O(N__37040),
            .I(encoder1_position_12));
    LocalMux I__6190 (
            .O(N__37037),
            .I(encoder1_position_12));
    Odrv4 I__6189 (
            .O(N__37034),
            .I(encoder1_position_12));
    InMux I__6188 (
            .O(N__37027),
            .I(N__37024));
    LocalMux I__6187 (
            .O(N__37024),
            .I(N__37020));
    InMux I__6186 (
            .O(N__37023),
            .I(N__37017));
    Span4Mux_v I__6185 (
            .O(N__37020),
            .I(N__37014));
    LocalMux I__6184 (
            .O(N__37017),
            .I(N__37009));
    Span4Mux_h I__6183 (
            .O(N__37014),
            .I(N__37009));
    Odrv4 I__6182 (
            .O(N__37009),
            .I(data_out_frame_12_4));
    InMux I__6181 (
            .O(N__37006),
            .I(N__37002));
    InMux I__6180 (
            .O(N__37005),
            .I(N__36999));
    LocalMux I__6179 (
            .O(N__37002),
            .I(data_out_frame_5_7));
    LocalMux I__6178 (
            .O(N__36999),
            .I(data_out_frame_5_7));
    InMux I__6177 (
            .O(N__36994),
            .I(N__36991));
    LocalMux I__6176 (
            .O(N__36991),
            .I(\c0.n5_adj_3475 ));
    CascadeMux I__6175 (
            .O(N__36988),
            .I(N__36983));
    CascadeMux I__6174 (
            .O(N__36987),
            .I(N__36980));
    CascadeMux I__6173 (
            .O(N__36986),
            .I(N__36977));
    InMux I__6172 (
            .O(N__36983),
            .I(N__36973));
    InMux I__6171 (
            .O(N__36980),
            .I(N__36970));
    InMux I__6170 (
            .O(N__36977),
            .I(N__36962));
    InMux I__6169 (
            .O(N__36976),
            .I(N__36955));
    LocalMux I__6168 (
            .O(N__36973),
            .I(N__36944));
    LocalMux I__6167 (
            .O(N__36970),
            .I(N__36944));
    InMux I__6166 (
            .O(N__36969),
            .I(N__36941));
    InMux I__6165 (
            .O(N__36968),
            .I(N__36932));
    InMux I__6164 (
            .O(N__36967),
            .I(N__36932));
    InMux I__6163 (
            .O(N__36966),
            .I(N__36932));
    InMux I__6162 (
            .O(N__36965),
            .I(N__36927));
    LocalMux I__6161 (
            .O(N__36962),
            .I(N__36922));
    InMux I__6160 (
            .O(N__36961),
            .I(N__36917));
    InMux I__6159 (
            .O(N__36960),
            .I(N__36917));
    InMux I__6158 (
            .O(N__36959),
            .I(N__36912));
    InMux I__6157 (
            .O(N__36958),
            .I(N__36912));
    LocalMux I__6156 (
            .O(N__36955),
            .I(N__36909));
    InMux I__6155 (
            .O(N__36954),
            .I(N__36905));
    InMux I__6154 (
            .O(N__36953),
            .I(N__36902));
    InMux I__6153 (
            .O(N__36952),
            .I(N__36897));
    InMux I__6152 (
            .O(N__36951),
            .I(N__36897));
    InMux I__6151 (
            .O(N__36950),
            .I(N__36894));
    InMux I__6150 (
            .O(N__36949),
            .I(N__36891));
    Span4Mux_h I__6149 (
            .O(N__36944),
            .I(N__36886));
    LocalMux I__6148 (
            .O(N__36941),
            .I(N__36886));
    InMux I__6147 (
            .O(N__36940),
            .I(N__36880));
    InMux I__6146 (
            .O(N__36939),
            .I(N__36880));
    LocalMux I__6145 (
            .O(N__36932),
            .I(N__36877));
    InMux I__6144 (
            .O(N__36931),
            .I(N__36871));
    InMux I__6143 (
            .O(N__36930),
            .I(N__36871));
    LocalMux I__6142 (
            .O(N__36927),
            .I(N__36868));
    CascadeMux I__6141 (
            .O(N__36926),
            .I(N__36865));
    InMux I__6140 (
            .O(N__36925),
            .I(N__36861));
    Span4Mux_v I__6139 (
            .O(N__36922),
            .I(N__36858));
    LocalMux I__6138 (
            .O(N__36917),
            .I(N__36853));
    LocalMux I__6137 (
            .O(N__36912),
            .I(N__36853));
    Span4Mux_h I__6136 (
            .O(N__36909),
            .I(N__36850));
    InMux I__6135 (
            .O(N__36908),
            .I(N__36847));
    LocalMux I__6134 (
            .O(N__36905),
            .I(N__36844));
    LocalMux I__6133 (
            .O(N__36902),
            .I(N__36839));
    LocalMux I__6132 (
            .O(N__36897),
            .I(N__36839));
    LocalMux I__6131 (
            .O(N__36894),
            .I(N__36834));
    LocalMux I__6130 (
            .O(N__36891),
            .I(N__36834));
    Span4Mux_v I__6129 (
            .O(N__36886),
            .I(N__36831));
    InMux I__6128 (
            .O(N__36885),
            .I(N__36828));
    LocalMux I__6127 (
            .O(N__36880),
            .I(N__36823));
    Span4Mux_h I__6126 (
            .O(N__36877),
            .I(N__36823));
    InMux I__6125 (
            .O(N__36876),
            .I(N__36820));
    LocalMux I__6124 (
            .O(N__36871),
            .I(N__36815));
    Span4Mux_v I__6123 (
            .O(N__36868),
            .I(N__36815));
    InMux I__6122 (
            .O(N__36865),
            .I(N__36810));
    InMux I__6121 (
            .O(N__36864),
            .I(N__36810));
    LocalMux I__6120 (
            .O(N__36861),
            .I(N__36803));
    Span4Mux_v I__6119 (
            .O(N__36858),
            .I(N__36803));
    Span4Mux_v I__6118 (
            .O(N__36853),
            .I(N__36803));
    Span4Mux_v I__6117 (
            .O(N__36850),
            .I(N__36800));
    LocalMux I__6116 (
            .O(N__36847),
            .I(N__36789));
    Span4Mux_v I__6115 (
            .O(N__36844),
            .I(N__36789));
    Span4Mux_h I__6114 (
            .O(N__36839),
            .I(N__36789));
    Span4Mux_h I__6113 (
            .O(N__36834),
            .I(N__36789));
    Span4Mux_h I__6112 (
            .O(N__36831),
            .I(N__36789));
    LocalMux I__6111 (
            .O(N__36828),
            .I(N__36778));
    Span4Mux_v I__6110 (
            .O(N__36823),
            .I(N__36778));
    LocalMux I__6109 (
            .O(N__36820),
            .I(N__36778));
    Span4Mux_h I__6108 (
            .O(N__36815),
            .I(N__36778));
    LocalMux I__6107 (
            .O(N__36810),
            .I(N__36778));
    Odrv4 I__6106 (
            .O(N__36803),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6105 (
            .O(N__36800),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6104 (
            .O(N__36789),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__6103 (
            .O(N__36778),
            .I(\c0.byte_transmit_counter_2 ));
    CascadeMux I__6102 (
            .O(N__36769),
            .I(\c0.n21576_cascade_ ));
    CascadeMux I__6101 (
            .O(N__36766),
            .I(N__36761));
    InMux I__6100 (
            .O(N__36765),
            .I(N__36750));
    InMux I__6099 (
            .O(N__36764),
            .I(N__36750));
    InMux I__6098 (
            .O(N__36761),
            .I(N__36747));
    CascadeMux I__6097 (
            .O(N__36760),
            .I(N__36743));
    InMux I__6096 (
            .O(N__36759),
            .I(N__36740));
    InMux I__6095 (
            .O(N__36758),
            .I(N__36737));
    CascadeMux I__6094 (
            .O(N__36757),
            .I(N__36732));
    InMux I__6093 (
            .O(N__36756),
            .I(N__36720));
    InMux I__6092 (
            .O(N__36755),
            .I(N__36717));
    LocalMux I__6091 (
            .O(N__36750),
            .I(N__36711));
    LocalMux I__6090 (
            .O(N__36747),
            .I(N__36711));
    InMux I__6089 (
            .O(N__36746),
            .I(N__36708));
    InMux I__6088 (
            .O(N__36743),
            .I(N__36704));
    LocalMux I__6087 (
            .O(N__36740),
            .I(N__36690));
    LocalMux I__6086 (
            .O(N__36737),
            .I(N__36690));
    InMux I__6085 (
            .O(N__36736),
            .I(N__36687));
    InMux I__6084 (
            .O(N__36735),
            .I(N__36684));
    InMux I__6083 (
            .O(N__36732),
            .I(N__36679));
    InMux I__6082 (
            .O(N__36731),
            .I(N__36679));
    InMux I__6081 (
            .O(N__36730),
            .I(N__36670));
    InMux I__6080 (
            .O(N__36729),
            .I(N__36670));
    InMux I__6079 (
            .O(N__36728),
            .I(N__36670));
    InMux I__6078 (
            .O(N__36727),
            .I(N__36670));
    InMux I__6077 (
            .O(N__36726),
            .I(N__36661));
    InMux I__6076 (
            .O(N__36725),
            .I(N__36661));
    InMux I__6075 (
            .O(N__36724),
            .I(N__36661));
    InMux I__6074 (
            .O(N__36723),
            .I(N__36661));
    LocalMux I__6073 (
            .O(N__36720),
            .I(N__36656));
    LocalMux I__6072 (
            .O(N__36717),
            .I(N__36656));
    InMux I__6071 (
            .O(N__36716),
            .I(N__36653));
    Span4Mux_h I__6070 (
            .O(N__36711),
            .I(N__36648));
    LocalMux I__6069 (
            .O(N__36708),
            .I(N__36648));
    InMux I__6068 (
            .O(N__36707),
            .I(N__36645));
    LocalMux I__6067 (
            .O(N__36704),
            .I(N__36642));
    InMux I__6066 (
            .O(N__36703),
            .I(N__36637));
    InMux I__6065 (
            .O(N__36702),
            .I(N__36637));
    InMux I__6064 (
            .O(N__36701),
            .I(N__36634));
    InMux I__6063 (
            .O(N__36700),
            .I(N__36628));
    InMux I__6062 (
            .O(N__36699),
            .I(N__36628));
    InMux I__6061 (
            .O(N__36698),
            .I(N__36625));
    InMux I__6060 (
            .O(N__36697),
            .I(N__36618));
    InMux I__6059 (
            .O(N__36696),
            .I(N__36613));
    InMux I__6058 (
            .O(N__36695),
            .I(N__36613));
    Span4Mux_v I__6057 (
            .O(N__36690),
            .I(N__36608));
    LocalMux I__6056 (
            .O(N__36687),
            .I(N__36608));
    LocalMux I__6055 (
            .O(N__36684),
            .I(N__36595));
    LocalMux I__6054 (
            .O(N__36679),
            .I(N__36595));
    LocalMux I__6053 (
            .O(N__36670),
            .I(N__36595));
    LocalMux I__6052 (
            .O(N__36661),
            .I(N__36595));
    Span4Mux_h I__6051 (
            .O(N__36656),
            .I(N__36595));
    LocalMux I__6050 (
            .O(N__36653),
            .I(N__36595));
    Span4Mux_h I__6049 (
            .O(N__36648),
            .I(N__36590));
    LocalMux I__6048 (
            .O(N__36645),
            .I(N__36590));
    Span4Mux_h I__6047 (
            .O(N__36642),
            .I(N__36585));
    LocalMux I__6046 (
            .O(N__36637),
            .I(N__36580));
    LocalMux I__6045 (
            .O(N__36634),
            .I(N__36580));
    InMux I__6044 (
            .O(N__36633),
            .I(N__36577));
    LocalMux I__6043 (
            .O(N__36628),
            .I(N__36574));
    LocalMux I__6042 (
            .O(N__36625),
            .I(N__36571));
    InMux I__6041 (
            .O(N__36624),
            .I(N__36564));
    InMux I__6040 (
            .O(N__36623),
            .I(N__36564));
    InMux I__6039 (
            .O(N__36622),
            .I(N__36564));
    InMux I__6038 (
            .O(N__36621),
            .I(N__36561));
    LocalMux I__6037 (
            .O(N__36618),
            .I(N__36552));
    LocalMux I__6036 (
            .O(N__36613),
            .I(N__36552));
    Span4Mux_v I__6035 (
            .O(N__36608),
            .I(N__36552));
    Span4Mux_v I__6034 (
            .O(N__36595),
            .I(N__36552));
    Span4Mux_v I__6033 (
            .O(N__36590),
            .I(N__36549));
    InMux I__6032 (
            .O(N__36589),
            .I(N__36546));
    InMux I__6031 (
            .O(N__36588),
            .I(N__36543));
    Span4Mux_v I__6030 (
            .O(N__36585),
            .I(N__36538));
    Span4Mux_h I__6029 (
            .O(N__36580),
            .I(N__36538));
    LocalMux I__6028 (
            .O(N__36577),
            .I(N__36535));
    Span4Mux_h I__6027 (
            .O(N__36574),
            .I(N__36526));
    Span4Mux_v I__6026 (
            .O(N__36571),
            .I(N__36526));
    LocalMux I__6025 (
            .O(N__36564),
            .I(N__36526));
    LocalMux I__6024 (
            .O(N__36561),
            .I(N__36526));
    Span4Mux_v I__6023 (
            .O(N__36552),
            .I(N__36521));
    Span4Mux_h I__6022 (
            .O(N__36549),
            .I(N__36521));
    LocalMux I__6021 (
            .O(N__36546),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__6020 (
            .O(N__36543),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6019 (
            .O(N__36538),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6018 (
            .O(N__36535),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6017 (
            .O(N__36526),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__6016 (
            .O(N__36521),
            .I(\c0.byte_transmit_counter_1 ));
    CascadeMux I__6015 (
            .O(N__36508),
            .I(\c0.n21302_cascade_ ));
    CascadeMux I__6014 (
            .O(N__36505),
            .I(\c0.n21304_cascade_ ));
    InMux I__6013 (
            .O(N__36502),
            .I(N__36499));
    LocalMux I__6012 (
            .O(N__36499),
            .I(N__36496));
    Span4Mux_h I__6011 (
            .O(N__36496),
            .I(N__36493));
    Span4Mux_h I__6010 (
            .O(N__36493),
            .I(N__36490));
    Odrv4 I__6009 (
            .O(N__36490),
            .I(\c0.n21572 ));
    CascadeMux I__6008 (
            .O(N__36487),
            .I(N__36484));
    InMux I__6007 (
            .O(N__36484),
            .I(N__36478));
    InMux I__6006 (
            .O(N__36483),
            .I(N__36478));
    LocalMux I__6005 (
            .O(N__36478),
            .I(data_out_frame_5_4));
    InMux I__6004 (
            .O(N__36475),
            .I(N__36472));
    LocalMux I__6003 (
            .O(N__36472),
            .I(N__36469));
    Span4Mux_v I__6002 (
            .O(N__36469),
            .I(N__36466));
    Span4Mux_h I__6001 (
            .O(N__36466),
            .I(N__36463));
    Odrv4 I__6000 (
            .O(N__36463),
            .I(\c0.n21465 ));
    InMux I__5999 (
            .O(N__36460),
            .I(N__36456));
    InMux I__5998 (
            .O(N__36459),
            .I(N__36453));
    LocalMux I__5997 (
            .O(N__36456),
            .I(\c0.data_out_frame_5_0 ));
    LocalMux I__5996 (
            .O(N__36453),
            .I(\c0.data_out_frame_5_0 ));
    InMux I__5995 (
            .O(N__36448),
            .I(N__36445));
    LocalMux I__5994 (
            .O(N__36445),
            .I(N__36442));
    Span4Mux_v I__5993 (
            .O(N__36442),
            .I(N__36438));
    InMux I__5992 (
            .O(N__36441),
            .I(N__36435));
    Odrv4 I__5991 (
            .O(N__36438),
            .I(control_mode_5));
    LocalMux I__5990 (
            .O(N__36435),
            .I(control_mode_5));
    InMux I__5989 (
            .O(N__36430),
            .I(N__36427));
    LocalMux I__5988 (
            .O(N__36427),
            .I(N__36424));
    Span4Mux_v I__5987 (
            .O(N__36424),
            .I(N__36421));
    Odrv4 I__5986 (
            .O(N__36421),
            .I(\c0.n21638 ));
    CascadeMux I__5985 (
            .O(N__36418),
            .I(N__36415));
    InMux I__5984 (
            .O(N__36415),
            .I(N__36412));
    LocalMux I__5983 (
            .O(N__36412),
            .I(N__36409));
    Span4Mux_h I__5982 (
            .O(N__36409),
            .I(N__36406));
    Odrv4 I__5981 (
            .O(N__36406),
            .I(\c0.n11_adj_3462 ));
    InMux I__5980 (
            .O(N__36403),
            .I(N__36399));
    InMux I__5979 (
            .O(N__36402),
            .I(N__36396));
    LocalMux I__5978 (
            .O(N__36399),
            .I(N__36393));
    LocalMux I__5977 (
            .O(N__36396),
            .I(data_out_frame_5_2));
    Odrv12 I__5976 (
            .O(N__36393),
            .I(data_out_frame_5_2));
    InMux I__5975 (
            .O(N__36388),
            .I(N__36385));
    LocalMux I__5974 (
            .O(N__36385),
            .I(N__36382));
    Span4Mux_h I__5973 (
            .O(N__36382),
            .I(N__36379));
    Odrv4 I__5972 (
            .O(N__36379),
            .I(\c0.rx.n9 ));
    InMux I__5971 (
            .O(N__36376),
            .I(N__36373));
    LocalMux I__5970 (
            .O(N__36373),
            .I(\c0.n11_adj_3325 ));
    InMux I__5969 (
            .O(N__36370),
            .I(N__36366));
    CascadeMux I__5968 (
            .O(N__36369),
            .I(N__36363));
    LocalMux I__5967 (
            .O(N__36366),
            .I(N__36360));
    InMux I__5966 (
            .O(N__36363),
            .I(N__36357));
    Span4Mux_v I__5965 (
            .O(N__36360),
            .I(N__36353));
    LocalMux I__5964 (
            .O(N__36357),
            .I(N__36350));
    InMux I__5963 (
            .O(N__36356),
            .I(N__36347));
    Span4Mux_h I__5962 (
            .O(N__36353),
            .I(N__36344));
    Span4Mux_h I__5961 (
            .O(N__36350),
            .I(N__36341));
    LocalMux I__5960 (
            .O(N__36347),
            .I(encoder1_position_8));
    Odrv4 I__5959 (
            .O(N__36344),
            .I(encoder1_position_8));
    Odrv4 I__5958 (
            .O(N__36341),
            .I(encoder1_position_8));
    CascadeMux I__5957 (
            .O(N__36334),
            .I(N__36331));
    InMux I__5956 (
            .O(N__36331),
            .I(N__36325));
    InMux I__5955 (
            .O(N__36330),
            .I(N__36325));
    LocalMux I__5954 (
            .O(N__36325),
            .I(data_out_frame_12_0));
    CascadeMux I__5953 (
            .O(N__36322),
            .I(N__36319));
    InMux I__5952 (
            .O(N__36319),
            .I(N__36315));
    InMux I__5951 (
            .O(N__36318),
            .I(N__36312));
    LocalMux I__5950 (
            .O(N__36315),
            .I(N__36308));
    LocalMux I__5949 (
            .O(N__36312),
            .I(N__36305));
    InMux I__5948 (
            .O(N__36311),
            .I(N__36302));
    Span4Mux_h I__5947 (
            .O(N__36308),
            .I(N__36299));
    Odrv4 I__5946 (
            .O(N__36305),
            .I(encoder1_position_23));
    LocalMux I__5945 (
            .O(N__36302),
            .I(encoder1_position_23));
    Odrv4 I__5944 (
            .O(N__36299),
            .I(encoder1_position_23));
    CascadeMux I__5943 (
            .O(N__36292),
            .I(N__36288));
    InMux I__5942 (
            .O(N__36291),
            .I(N__36285));
    InMux I__5941 (
            .O(N__36288),
            .I(N__36282));
    LocalMux I__5940 (
            .O(N__36285),
            .I(data_out_frame_11_7));
    LocalMux I__5939 (
            .O(N__36282),
            .I(data_out_frame_11_7));
    InMux I__5938 (
            .O(N__36277),
            .I(N__36274));
    LocalMux I__5937 (
            .O(N__36274),
            .I(N__36271));
    Span4Mux_v I__5936 (
            .O(N__36271),
            .I(N__36268));
    Span4Mux_h I__5935 (
            .O(N__36268),
            .I(N__36265));
    Odrv4 I__5934 (
            .O(N__36265),
            .I(n2317));
    InMux I__5933 (
            .O(N__36262),
            .I(N__36251));
    InMux I__5932 (
            .O(N__36261),
            .I(N__36240));
    InMux I__5931 (
            .O(N__36260),
            .I(N__36240));
    InMux I__5930 (
            .O(N__36259),
            .I(N__36231));
    InMux I__5929 (
            .O(N__36258),
            .I(N__36231));
    InMux I__5928 (
            .O(N__36257),
            .I(N__36231));
    InMux I__5927 (
            .O(N__36256),
            .I(N__36231));
    InMux I__5926 (
            .O(N__36255),
            .I(N__36218));
    InMux I__5925 (
            .O(N__36254),
            .I(N__36215));
    LocalMux I__5924 (
            .O(N__36251),
            .I(N__36212));
    InMux I__5923 (
            .O(N__36250),
            .I(N__36207));
    InMux I__5922 (
            .O(N__36249),
            .I(N__36207));
    InMux I__5921 (
            .O(N__36248),
            .I(N__36204));
    InMux I__5920 (
            .O(N__36247),
            .I(N__36201));
    InMux I__5919 (
            .O(N__36246),
            .I(N__36196));
    InMux I__5918 (
            .O(N__36245),
            .I(N__36196));
    LocalMux I__5917 (
            .O(N__36240),
            .I(N__36191));
    LocalMux I__5916 (
            .O(N__36231),
            .I(N__36191));
    InMux I__5915 (
            .O(N__36230),
            .I(N__36184));
    InMux I__5914 (
            .O(N__36229),
            .I(N__36184));
    InMux I__5913 (
            .O(N__36228),
            .I(N__36184));
    InMux I__5912 (
            .O(N__36227),
            .I(N__36181));
    InMux I__5911 (
            .O(N__36226),
            .I(N__36169));
    InMux I__5910 (
            .O(N__36225),
            .I(N__36169));
    InMux I__5909 (
            .O(N__36224),
            .I(N__36166));
    InMux I__5908 (
            .O(N__36223),
            .I(N__36159));
    InMux I__5907 (
            .O(N__36222),
            .I(N__36159));
    InMux I__5906 (
            .O(N__36221),
            .I(N__36159));
    LocalMux I__5905 (
            .O(N__36218),
            .I(N__36150));
    LocalMux I__5904 (
            .O(N__36215),
            .I(N__36150));
    Span4Mux_v I__5903 (
            .O(N__36212),
            .I(N__36150));
    LocalMux I__5902 (
            .O(N__36207),
            .I(N__36150));
    LocalMux I__5901 (
            .O(N__36204),
            .I(N__36141));
    LocalMux I__5900 (
            .O(N__36201),
            .I(N__36141));
    LocalMux I__5899 (
            .O(N__36196),
            .I(N__36141));
    Span4Mux_v I__5898 (
            .O(N__36191),
            .I(N__36141));
    LocalMux I__5897 (
            .O(N__36184),
            .I(N__36138));
    LocalMux I__5896 (
            .O(N__36181),
            .I(N__36135));
    InMux I__5895 (
            .O(N__36180),
            .I(N__36120));
    InMux I__5894 (
            .O(N__36179),
            .I(N__36120));
    InMux I__5893 (
            .O(N__36178),
            .I(N__36120));
    InMux I__5892 (
            .O(N__36177),
            .I(N__36120));
    InMux I__5891 (
            .O(N__36176),
            .I(N__36120));
    InMux I__5890 (
            .O(N__36175),
            .I(N__36120));
    InMux I__5889 (
            .O(N__36174),
            .I(N__36120));
    LocalMux I__5888 (
            .O(N__36169),
            .I(N__36117));
    LocalMux I__5887 (
            .O(N__36166),
            .I(N__36112));
    LocalMux I__5886 (
            .O(N__36159),
            .I(N__36112));
    Span4Mux_v I__5885 (
            .O(N__36150),
            .I(N__36107));
    Span4Mux_v I__5884 (
            .O(N__36141),
            .I(N__36107));
    Span4Mux_h I__5883 (
            .O(N__36138),
            .I(N__36102));
    Span4Mux_h I__5882 (
            .O(N__36135),
            .I(N__36102));
    LocalMux I__5881 (
            .O(N__36120),
            .I(N__36095));
    Span4Mux_h I__5880 (
            .O(N__36117),
            .I(N__36095));
    Span4Mux_v I__5879 (
            .O(N__36112),
            .I(N__36095));
    Sp12to4 I__5878 (
            .O(N__36107),
            .I(N__36092));
    Span4Mux_v I__5877 (
            .O(N__36102),
            .I(N__36089));
    Odrv4 I__5876 (
            .O(N__36095),
            .I(count_enable_adj_3586));
    Odrv12 I__5875 (
            .O(N__36092),
            .I(count_enable_adj_3586));
    Odrv4 I__5874 (
            .O(N__36089),
            .I(count_enable_adj_3586));
    InMux I__5873 (
            .O(N__36082),
            .I(N__36079));
    LocalMux I__5872 (
            .O(N__36079),
            .I(N__36075));
    InMux I__5871 (
            .O(N__36078),
            .I(N__36071));
    Span4Mux_h I__5870 (
            .O(N__36075),
            .I(N__36068));
    InMux I__5869 (
            .O(N__36074),
            .I(N__36065));
    LocalMux I__5868 (
            .O(N__36071),
            .I(N__36062));
    Span4Mux_h I__5867 (
            .O(N__36068),
            .I(N__36059));
    LocalMux I__5866 (
            .O(N__36065),
            .I(N__36054));
    Span4Mux_v I__5865 (
            .O(N__36062),
            .I(N__36054));
    Odrv4 I__5864 (
            .O(N__36059),
            .I(encoder1_position_28));
    Odrv4 I__5863 (
            .O(N__36054),
            .I(encoder1_position_28));
    InMux I__5862 (
            .O(N__36049),
            .I(N__36045));
    InMux I__5861 (
            .O(N__36048),
            .I(N__36042));
    LocalMux I__5860 (
            .O(N__36045),
            .I(data_out_frame_5_6));
    LocalMux I__5859 (
            .O(N__36042),
            .I(data_out_frame_5_6));
    InMux I__5858 (
            .O(N__36037),
            .I(N__36034));
    LocalMux I__5857 (
            .O(N__36034),
            .I(N__36030));
    InMux I__5856 (
            .O(N__36033),
            .I(N__36027));
    Span4Mux_h I__5855 (
            .O(N__36030),
            .I(N__36024));
    LocalMux I__5854 (
            .O(N__36027),
            .I(data_out_frame_29_3));
    Odrv4 I__5853 (
            .O(N__36024),
            .I(data_out_frame_29_3));
    InMux I__5852 (
            .O(N__36019),
            .I(N__36015));
    InMux I__5851 (
            .O(N__36018),
            .I(N__36012));
    LocalMux I__5850 (
            .O(N__36015),
            .I(\c0.data_out_frame_28_3 ));
    LocalMux I__5849 (
            .O(N__36012),
            .I(\c0.data_out_frame_28_3 ));
    CascadeMux I__5848 (
            .O(N__36007),
            .I(N__36004));
    InMux I__5847 (
            .O(N__36004),
            .I(N__36001));
    LocalMux I__5846 (
            .O(N__36001),
            .I(N__35996));
    InMux I__5845 (
            .O(N__36000),
            .I(N__35993));
    CascadeMux I__5844 (
            .O(N__35999),
            .I(N__35990));
    Span4Mux_v I__5843 (
            .O(N__35996),
            .I(N__35985));
    LocalMux I__5842 (
            .O(N__35993),
            .I(N__35985));
    InMux I__5841 (
            .O(N__35990),
            .I(N__35982));
    Span4Mux_v I__5840 (
            .O(N__35985),
            .I(N__35979));
    LocalMux I__5839 (
            .O(N__35982),
            .I(N__35976));
    Span4Mux_h I__5838 (
            .O(N__35979),
            .I(N__35973));
    Span12Mux_h I__5837 (
            .O(N__35976),
            .I(N__35970));
    Odrv4 I__5836 (
            .O(N__35973),
            .I(\c0.n9753 ));
    Odrv12 I__5835 (
            .O(N__35970),
            .I(\c0.n9753 ));
    CascadeMux I__5834 (
            .O(N__35965),
            .I(\c0.n26_adj_3382_cascade_ ));
    InMux I__5833 (
            .O(N__35962),
            .I(N__35959));
    LocalMux I__5832 (
            .O(N__35959),
            .I(N__35956));
    Odrv4 I__5831 (
            .O(N__35956),
            .I(\c0.n21314 ));
    InMux I__5830 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__5829 (
            .O(N__35950),
            .I(N__35947));
    Span4Mux_v I__5828 (
            .O(N__35947),
            .I(N__35944));
    Odrv4 I__5827 (
            .O(N__35944),
            .I(\c0.n21316 ));
    InMux I__5826 (
            .O(N__35941),
            .I(N__35938));
    LocalMux I__5825 (
            .O(N__35938),
            .I(N__35935));
    Span12Mux_v I__5824 (
            .O(N__35935),
            .I(N__35932));
    Odrv12 I__5823 (
            .O(N__35932),
            .I(\c0.n21562 ));
    CascadeMux I__5822 (
            .O(N__35929),
            .I(\c0.n21322_cascade_ ));
    InMux I__5821 (
            .O(N__35926),
            .I(N__35923));
    LocalMux I__5820 (
            .O(N__35923),
            .I(N__35920));
    Span4Mux_v I__5819 (
            .O(N__35920),
            .I(N__35917));
    Odrv4 I__5818 (
            .O(N__35917),
            .I(n10_adj_3594));
    InMux I__5817 (
            .O(N__35914),
            .I(N__35910));
    InMux I__5816 (
            .O(N__35913),
            .I(N__35907));
    LocalMux I__5815 (
            .O(N__35910),
            .I(data_out_frame_7_2));
    LocalMux I__5814 (
            .O(N__35907),
            .I(data_out_frame_7_2));
    InMux I__5813 (
            .O(N__35902),
            .I(N__35899));
    LocalMux I__5812 (
            .O(N__35899),
            .I(\c0.n5_adj_3106 ));
    InMux I__5811 (
            .O(N__35896),
            .I(N__35892));
    CascadeMux I__5810 (
            .O(N__35895),
            .I(N__35888));
    LocalMux I__5809 (
            .O(N__35892),
            .I(N__35885));
    InMux I__5808 (
            .O(N__35891),
            .I(N__35882));
    InMux I__5807 (
            .O(N__35888),
            .I(N__35879));
    Odrv12 I__5806 (
            .O(N__35885),
            .I(encoder0_position_26));
    LocalMux I__5805 (
            .O(N__35882),
            .I(encoder0_position_26));
    LocalMux I__5804 (
            .O(N__35879),
            .I(encoder0_position_26));
    InMux I__5803 (
            .O(N__35872),
            .I(N__35868));
    InMux I__5802 (
            .O(N__35871),
            .I(N__35865));
    LocalMux I__5801 (
            .O(N__35868),
            .I(data_out_frame_6_2));
    LocalMux I__5800 (
            .O(N__35865),
            .I(data_out_frame_6_2));
    InMux I__5799 (
            .O(N__35860),
            .I(N__35854));
    InMux I__5798 (
            .O(N__35859),
            .I(N__35854));
    LocalMux I__5797 (
            .O(N__35854),
            .I(\c0.data_out_frame_0_2 ));
    CascadeMux I__5796 (
            .O(N__35851),
            .I(\c0.n21473_cascade_ ));
    InMux I__5795 (
            .O(N__35848),
            .I(N__35845));
    LocalMux I__5794 (
            .O(N__35845),
            .I(N__35842));
    Odrv4 I__5793 (
            .O(N__35842),
            .I(\c0.n6_adj_3105 ));
    CascadeMux I__5792 (
            .O(N__35839),
            .I(N__35836));
    InMux I__5791 (
            .O(N__35836),
            .I(N__35833));
    LocalMux I__5790 (
            .O(N__35833),
            .I(N__35830));
    Span4Mux_v I__5789 (
            .O(N__35830),
            .I(N__35826));
    InMux I__5788 (
            .O(N__35829),
            .I(N__35823));
    Span4Mux_h I__5787 (
            .O(N__35826),
            .I(N__35820));
    LocalMux I__5786 (
            .O(N__35823),
            .I(data_out_frame_28_6));
    Odrv4 I__5785 (
            .O(N__35820),
            .I(data_out_frame_28_6));
    InMux I__5784 (
            .O(N__35815),
            .I(N__35811));
    InMux I__5783 (
            .O(N__35814),
            .I(N__35808));
    LocalMux I__5782 (
            .O(N__35811),
            .I(\c0.data_out_frame_0_3 ));
    LocalMux I__5781 (
            .O(N__35808),
            .I(\c0.data_out_frame_0_3 ));
    SRMux I__5780 (
            .O(N__35803),
            .I(N__35800));
    LocalMux I__5779 (
            .O(N__35800),
            .I(N__35797));
    Span4Mux_h I__5778 (
            .O(N__35797),
            .I(N__35794));
    Odrv4 I__5777 (
            .O(N__35794),
            .I(\c0.n6_adj_3150 ));
    InMux I__5776 (
            .O(N__35791),
            .I(N__35788));
    LocalMux I__5775 (
            .O(N__35788),
            .I(N__35785));
    Span4Mux_h I__5774 (
            .O(N__35785),
            .I(N__35782));
    Odrv4 I__5773 (
            .O(N__35782),
            .I(n2333));
    InMux I__5772 (
            .O(N__35779),
            .I(N__35776));
    LocalMux I__5771 (
            .O(N__35776),
            .I(N__35773));
    Span4Mux_h I__5770 (
            .O(N__35773),
            .I(N__35770));
    Odrv4 I__5769 (
            .O(N__35770),
            .I(\c0.n21319 ));
    InMux I__5768 (
            .O(N__35767),
            .I(N__35764));
    LocalMux I__5767 (
            .O(N__35764),
            .I(N__35761));
    Span4Mux_v I__5766 (
            .O(N__35761),
            .I(N__35757));
    CascadeMux I__5765 (
            .O(N__35760),
            .I(N__35753));
    Span4Mux_h I__5764 (
            .O(N__35757),
            .I(N__35750));
    InMux I__5763 (
            .O(N__35756),
            .I(N__35747));
    InMux I__5762 (
            .O(N__35753),
            .I(N__35744));
    Odrv4 I__5761 (
            .O(N__35750),
            .I(encoder0_position_18));
    LocalMux I__5760 (
            .O(N__35747),
            .I(encoder0_position_18));
    LocalMux I__5759 (
            .O(N__35744),
            .I(encoder0_position_18));
    InMux I__5758 (
            .O(N__35737),
            .I(N__35734));
    LocalMux I__5757 (
            .O(N__35734),
            .I(\c0.n21317 ));
    InMux I__5756 (
            .O(N__35731),
            .I(N__35725));
    InMux I__5755 (
            .O(N__35730),
            .I(N__35706));
    InMux I__5754 (
            .O(N__35729),
            .I(N__35701));
    InMux I__5753 (
            .O(N__35728),
            .I(N__35701));
    LocalMux I__5752 (
            .O(N__35725),
            .I(N__35698));
    InMux I__5751 (
            .O(N__35724),
            .I(N__35695));
    InMux I__5750 (
            .O(N__35723),
            .I(N__35692));
    InMux I__5749 (
            .O(N__35722),
            .I(N__35689));
    InMux I__5748 (
            .O(N__35721),
            .I(N__35684));
    InMux I__5747 (
            .O(N__35720),
            .I(N__35681));
    InMux I__5746 (
            .O(N__35719),
            .I(N__35678));
    InMux I__5745 (
            .O(N__35718),
            .I(N__35663));
    InMux I__5744 (
            .O(N__35717),
            .I(N__35663));
    InMux I__5743 (
            .O(N__35716),
            .I(N__35663));
    InMux I__5742 (
            .O(N__35715),
            .I(N__35663));
    InMux I__5741 (
            .O(N__35714),
            .I(N__35663));
    InMux I__5740 (
            .O(N__35713),
            .I(N__35663));
    InMux I__5739 (
            .O(N__35712),
            .I(N__35663));
    InMux I__5738 (
            .O(N__35711),
            .I(N__35656));
    InMux I__5737 (
            .O(N__35710),
            .I(N__35656));
    InMux I__5736 (
            .O(N__35709),
            .I(N__35656));
    LocalMux I__5735 (
            .O(N__35706),
            .I(N__35645));
    LocalMux I__5734 (
            .O(N__35701),
            .I(N__35645));
    Span4Mux_h I__5733 (
            .O(N__35698),
            .I(N__35645));
    LocalMux I__5732 (
            .O(N__35695),
            .I(N__35645));
    LocalMux I__5731 (
            .O(N__35692),
            .I(N__35645));
    LocalMux I__5730 (
            .O(N__35689),
            .I(N__35642));
    InMux I__5729 (
            .O(N__35688),
            .I(N__35629));
    InMux I__5728 (
            .O(N__35687),
            .I(N__35626));
    LocalMux I__5727 (
            .O(N__35684),
            .I(N__35621));
    LocalMux I__5726 (
            .O(N__35681),
            .I(N__35621));
    LocalMux I__5725 (
            .O(N__35678),
            .I(N__35614));
    LocalMux I__5724 (
            .O(N__35663),
            .I(N__35614));
    LocalMux I__5723 (
            .O(N__35656),
            .I(N__35614));
    Span4Mux_v I__5722 (
            .O(N__35645),
            .I(N__35609));
    Span4Mux_h I__5721 (
            .O(N__35642),
            .I(N__35609));
    InMux I__5720 (
            .O(N__35641),
            .I(N__35604));
    InMux I__5719 (
            .O(N__35640),
            .I(N__35604));
    InMux I__5718 (
            .O(N__35639),
            .I(N__35587));
    InMux I__5717 (
            .O(N__35638),
            .I(N__35587));
    InMux I__5716 (
            .O(N__35637),
            .I(N__35587));
    InMux I__5715 (
            .O(N__35636),
            .I(N__35587));
    InMux I__5714 (
            .O(N__35635),
            .I(N__35587));
    InMux I__5713 (
            .O(N__35634),
            .I(N__35587));
    InMux I__5712 (
            .O(N__35633),
            .I(N__35587));
    InMux I__5711 (
            .O(N__35632),
            .I(N__35587));
    LocalMux I__5710 (
            .O(N__35629),
            .I(N__35582));
    LocalMux I__5709 (
            .O(N__35626),
            .I(N__35582));
    Span4Mux_h I__5708 (
            .O(N__35621),
            .I(N__35577));
    Span4Mux_v I__5707 (
            .O(N__35614),
            .I(N__35577));
    Span4Mux_h I__5706 (
            .O(N__35609),
            .I(N__35574));
    LocalMux I__5705 (
            .O(N__35604),
            .I(count_enable));
    LocalMux I__5704 (
            .O(N__35587),
            .I(count_enable));
    Odrv12 I__5703 (
            .O(N__35582),
            .I(count_enable));
    Odrv4 I__5702 (
            .O(N__35577),
            .I(count_enable));
    Odrv4 I__5701 (
            .O(N__35574),
            .I(count_enable));
    InMux I__5700 (
            .O(N__35563),
            .I(N__35560));
    LocalMux I__5699 (
            .O(N__35560),
            .I(N__35557));
    Span4Mux_h I__5698 (
            .O(N__35557),
            .I(N__35554));
    Span4Mux_h I__5697 (
            .O(N__35554),
            .I(N__35551));
    Odrv4 I__5696 (
            .O(N__35551),
            .I(n2252));
    InMux I__5695 (
            .O(N__35548),
            .I(N__35544));
    CascadeMux I__5694 (
            .O(N__35547),
            .I(N__35541));
    LocalMux I__5693 (
            .O(N__35544),
            .I(N__35538));
    InMux I__5692 (
            .O(N__35541),
            .I(N__35535));
    Span4Mux_v I__5691 (
            .O(N__35538),
            .I(N__35530));
    LocalMux I__5690 (
            .O(N__35535),
            .I(N__35530));
    Span4Mux_h I__5689 (
            .O(N__35530),
            .I(N__35526));
    InMux I__5688 (
            .O(N__35529),
            .I(N__35523));
    Span4Mux_h I__5687 (
            .O(N__35526),
            .I(N__35520));
    LocalMux I__5686 (
            .O(N__35523),
            .I(encoder0_position_27));
    Odrv4 I__5685 (
            .O(N__35520),
            .I(encoder0_position_27));
    InMux I__5684 (
            .O(N__35515),
            .I(N__35511));
    InMux I__5683 (
            .O(N__35514),
            .I(N__35508));
    LocalMux I__5682 (
            .O(N__35511),
            .I(data_out_frame_7_3));
    LocalMux I__5681 (
            .O(N__35508),
            .I(data_out_frame_7_3));
    InMux I__5680 (
            .O(N__35503),
            .I(N__35500));
    LocalMux I__5679 (
            .O(N__35500),
            .I(N__35496));
    InMux I__5678 (
            .O(N__35499),
            .I(N__35493));
    Span4Mux_h I__5677 (
            .O(N__35496),
            .I(N__35490));
    LocalMux I__5676 (
            .O(N__35493),
            .I(data_out_frame_6_3));
    Odrv4 I__5675 (
            .O(N__35490),
            .I(data_out_frame_6_3));
    InMux I__5674 (
            .O(N__35485),
            .I(N__35482));
    LocalMux I__5673 (
            .O(N__35482),
            .I(\c0.n5_adj_3380 ));
    InMux I__5672 (
            .O(N__35479),
            .I(N__35476));
    LocalMux I__5671 (
            .O(N__35476),
            .I(\c0.n21320 ));
    InMux I__5670 (
            .O(N__35473),
            .I(N__35468));
    InMux I__5669 (
            .O(N__35472),
            .I(N__35465));
    InMux I__5668 (
            .O(N__35471),
            .I(N__35462));
    LocalMux I__5667 (
            .O(N__35468),
            .I(N__35459));
    LocalMux I__5666 (
            .O(N__35465),
            .I(N__35456));
    LocalMux I__5665 (
            .O(N__35462),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__5664 (
            .O(N__35459),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__5663 (
            .O(N__35456),
            .I(\c0.FRAME_MATCHER_state_8 ));
    SRMux I__5662 (
            .O(N__35449),
            .I(N__35446));
    LocalMux I__5661 (
            .O(N__35446),
            .I(N__35443));
    Span4Mux_h I__5660 (
            .O(N__35443),
            .I(N__35440));
    Odrv4 I__5659 (
            .O(N__35440),
            .I(\c0.n18675 ));
    InMux I__5658 (
            .O(N__35437),
            .I(N__35433));
    InMux I__5657 (
            .O(N__35436),
            .I(N__35430));
    LocalMux I__5656 (
            .O(N__35433),
            .I(N__35427));
    LocalMux I__5655 (
            .O(N__35430),
            .I(N__35424));
    Span4Mux_h I__5654 (
            .O(N__35427),
            .I(N__35420));
    Span4Mux_h I__5653 (
            .O(N__35424),
            .I(N__35415));
    InMux I__5652 (
            .O(N__35423),
            .I(N__35412));
    Sp12to4 I__5651 (
            .O(N__35420),
            .I(N__35409));
    InMux I__5650 (
            .O(N__35419),
            .I(N__35406));
    InMux I__5649 (
            .O(N__35418),
            .I(N__35403));
    Span4Mux_v I__5648 (
            .O(N__35415),
            .I(N__35398));
    LocalMux I__5647 (
            .O(N__35412),
            .I(N__35398));
    Span12Mux_v I__5646 (
            .O(N__35409),
            .I(N__35395));
    LocalMux I__5645 (
            .O(N__35406),
            .I(N__35392));
    LocalMux I__5644 (
            .O(N__35403),
            .I(N__35387));
    Span4Mux_h I__5643 (
            .O(N__35398),
            .I(N__35387));
    Odrv12 I__5642 (
            .O(N__35395),
            .I(n11289));
    Odrv4 I__5641 (
            .O(N__35392),
            .I(n11289));
    Odrv4 I__5640 (
            .O(N__35387),
            .I(n11289));
    InMux I__5639 (
            .O(N__35380),
            .I(N__35377));
    LocalMux I__5638 (
            .O(N__35377),
            .I(N__35372));
    InMux I__5637 (
            .O(N__35376),
            .I(N__35369));
    InMux I__5636 (
            .O(N__35375),
            .I(N__35366));
    Span4Mux_v I__5635 (
            .O(N__35372),
            .I(N__35363));
    LocalMux I__5634 (
            .O(N__35369),
            .I(\c0.FRAME_MATCHER_i_26 ));
    LocalMux I__5633 (
            .O(N__35366),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__5632 (
            .O(N__35363),
            .I(\c0.FRAME_MATCHER_i_26 ));
    CascadeMux I__5631 (
            .O(N__35356),
            .I(n2108_cascade_));
    SRMux I__5630 (
            .O(N__35353),
            .I(N__35350));
    LocalMux I__5629 (
            .O(N__35350),
            .I(N__35347));
    Odrv12 I__5628 (
            .O(N__35347),
            .I(\c0.n6_adj_3170 ));
    SRMux I__5627 (
            .O(N__35344),
            .I(N__35341));
    LocalMux I__5626 (
            .O(N__35341),
            .I(N__35338));
    Span4Mux_h I__5625 (
            .O(N__35338),
            .I(N__35335));
    Odrv4 I__5624 (
            .O(N__35335),
            .I(\c0.n6_adj_3165 ));
    InMux I__5623 (
            .O(N__35332),
            .I(N__35329));
    LocalMux I__5622 (
            .O(N__35329),
            .I(N__35324));
    InMux I__5621 (
            .O(N__35328),
            .I(N__35321));
    InMux I__5620 (
            .O(N__35327),
            .I(N__35318));
    Span4Mux_v I__5619 (
            .O(N__35324),
            .I(N__35315));
    LocalMux I__5618 (
            .O(N__35321),
            .I(\c0.FRAME_MATCHER_i_27 ));
    LocalMux I__5617 (
            .O(N__35318),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv4 I__5616 (
            .O(N__35315),
            .I(\c0.FRAME_MATCHER_i_27 ));
    SRMux I__5615 (
            .O(N__35308),
            .I(N__35305));
    LocalMux I__5614 (
            .O(N__35305),
            .I(\c0.n6_adj_3168 ));
    CascadeMux I__5613 (
            .O(N__35302),
            .I(N__35299));
    InMux I__5612 (
            .O(N__35299),
            .I(N__35296));
    LocalMux I__5611 (
            .O(N__35296),
            .I(N__35293));
    Span4Mux_h I__5610 (
            .O(N__35293),
            .I(N__35288));
    InMux I__5609 (
            .O(N__35292),
            .I(N__35285));
    InMux I__5608 (
            .O(N__35291),
            .I(N__35282));
    Span4Mux_v I__5607 (
            .O(N__35288),
            .I(N__35279));
    LocalMux I__5606 (
            .O(N__35285),
            .I(\c0.FRAME_MATCHER_i_28 ));
    LocalMux I__5605 (
            .O(N__35282),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__5604 (
            .O(N__35279),
            .I(\c0.FRAME_MATCHER_i_28 ));
    SRMux I__5603 (
            .O(N__35272),
            .I(N__35269));
    LocalMux I__5602 (
            .O(N__35269),
            .I(N__35266));
    Odrv12 I__5601 (
            .O(N__35266),
            .I(\c0.n6_adj_3166 ));
    SRMux I__5600 (
            .O(N__35263),
            .I(N__35260));
    LocalMux I__5599 (
            .O(N__35260),
            .I(N__35257));
    Span4Mux_s1_v I__5598 (
            .O(N__35257),
            .I(N__35254));
    Odrv4 I__5597 (
            .O(N__35254),
            .I(\c0.n6_adj_3159 ));
    InMux I__5596 (
            .O(N__35251),
            .I(N__35248));
    LocalMux I__5595 (
            .O(N__35248),
            .I(N__35243));
    InMux I__5594 (
            .O(N__35247),
            .I(N__35240));
    InMux I__5593 (
            .O(N__35246),
            .I(N__35237));
    Span4Mux_v I__5592 (
            .O(N__35243),
            .I(N__35234));
    LocalMux I__5591 (
            .O(N__35240),
            .I(\c0.FRAME_MATCHER_i_30 ));
    LocalMux I__5590 (
            .O(N__35237),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__5589 (
            .O(N__35234),
            .I(\c0.FRAME_MATCHER_i_30 ));
    SRMux I__5588 (
            .O(N__35227),
            .I(N__35224));
    LocalMux I__5587 (
            .O(N__35224),
            .I(N__35221));
    Odrv12 I__5586 (
            .O(N__35221),
            .I(\c0.n6_adj_3164 ));
    SRMux I__5585 (
            .O(N__35218),
            .I(N__35215));
    LocalMux I__5584 (
            .O(N__35215),
            .I(N__35212));
    Odrv12 I__5583 (
            .O(N__35212),
            .I(\c0.n18653 ));
    InMux I__5582 (
            .O(N__35209),
            .I(N__35204));
    InMux I__5581 (
            .O(N__35208),
            .I(N__35201));
    InMux I__5580 (
            .O(N__35207),
            .I(N__35198));
    LocalMux I__5579 (
            .O(N__35204),
            .I(N__35195));
    LocalMux I__5578 (
            .O(N__35201),
            .I(N__35192));
    LocalMux I__5577 (
            .O(N__35198),
            .I(N__35189));
    Span4Mux_v I__5576 (
            .O(N__35195),
            .I(N__35186));
    Span4Mux_h I__5575 (
            .O(N__35192),
            .I(N__35183));
    Span4Mux_h I__5574 (
            .O(N__35189),
            .I(N__35180));
    Odrv4 I__5573 (
            .O(N__35186),
            .I(\c0.FRAME_MATCHER_state_31_N_1736_2 ));
    Odrv4 I__5572 (
            .O(N__35183),
            .I(\c0.FRAME_MATCHER_state_31_N_1736_2 ));
    Odrv4 I__5571 (
            .O(N__35180),
            .I(\c0.FRAME_MATCHER_state_31_N_1736_2 ));
    InMux I__5570 (
            .O(N__35173),
            .I(N__35170));
    LocalMux I__5569 (
            .O(N__35170),
            .I(N__35167));
    Odrv4 I__5568 (
            .O(N__35167),
            .I(\c0.FRAME_MATCHER_state_31_N_1736_1 ));
    SRMux I__5567 (
            .O(N__35164),
            .I(N__35161));
    LocalMux I__5566 (
            .O(N__35161),
            .I(N__35158));
    Odrv4 I__5565 (
            .O(N__35158),
            .I(\c0.n6_adj_3176 ));
    InMux I__5564 (
            .O(N__35155),
            .I(N__35151));
    InMux I__5563 (
            .O(N__35154),
            .I(N__35147));
    LocalMux I__5562 (
            .O(N__35151),
            .I(N__35144));
    InMux I__5561 (
            .O(N__35150),
            .I(N__35141));
    LocalMux I__5560 (
            .O(N__35147),
            .I(\c0.n11433 ));
    Odrv4 I__5559 (
            .O(N__35144),
            .I(\c0.n11433 ));
    LocalMux I__5558 (
            .O(N__35141),
            .I(\c0.n11433 ));
    CascadeMux I__5557 (
            .O(N__35134),
            .I(N__35130));
    CascadeMux I__5556 (
            .O(N__35133),
            .I(N__35127));
    InMux I__5555 (
            .O(N__35130),
            .I(N__35124));
    InMux I__5554 (
            .O(N__35127),
            .I(N__35120));
    LocalMux I__5553 (
            .O(N__35124),
            .I(N__35117));
    InMux I__5552 (
            .O(N__35123),
            .I(N__35114));
    LocalMux I__5551 (
            .O(N__35120),
            .I(N__35111));
    Span4Mux_h I__5550 (
            .O(N__35117),
            .I(N__35104));
    LocalMux I__5549 (
            .O(N__35114),
            .I(N__35104));
    Span4Mux_v I__5548 (
            .O(N__35111),
            .I(N__35104));
    Span4Mux_v I__5547 (
            .O(N__35104),
            .I(N__35101));
    Span4Mux_v I__5546 (
            .O(N__35101),
            .I(N__35098));
    Odrv4 I__5545 (
            .O(N__35098),
            .I(\c0.n700 ));
    InMux I__5544 (
            .O(N__35095),
            .I(N__35092));
    LocalMux I__5543 (
            .O(N__35092),
            .I(N__35089));
    Span4Mux_h I__5542 (
            .O(N__35089),
            .I(N__35086));
    Odrv4 I__5541 (
            .O(N__35086),
            .I(\c0.n1 ));
    InMux I__5540 (
            .O(N__35083),
            .I(N__35080));
    LocalMux I__5539 (
            .O(N__35080),
            .I(N__35075));
    InMux I__5538 (
            .O(N__35079),
            .I(N__35072));
    InMux I__5537 (
            .O(N__35078),
            .I(N__35069));
    Span4Mux_v I__5536 (
            .O(N__35075),
            .I(N__35066));
    LocalMux I__5535 (
            .O(N__35072),
            .I(\c0.FRAME_MATCHER_i_21 ));
    LocalMux I__5534 (
            .O(N__35069),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv4 I__5533 (
            .O(N__35066),
            .I(\c0.FRAME_MATCHER_i_21 ));
    CascadeMux I__5532 (
            .O(N__35059),
            .I(N__35056));
    InMux I__5531 (
            .O(N__35056),
            .I(N__35052));
    InMux I__5530 (
            .O(N__35055),
            .I(N__35049));
    LocalMux I__5529 (
            .O(N__35052),
            .I(N__35046));
    LocalMux I__5528 (
            .O(N__35049),
            .I(N__35043));
    Span4Mux_v I__5527 (
            .O(N__35046),
            .I(N__35039));
    Span4Mux_v I__5526 (
            .O(N__35043),
            .I(N__35036));
    InMux I__5525 (
            .O(N__35042),
            .I(N__35033));
    Span4Mux_v I__5524 (
            .O(N__35039),
            .I(N__35030));
    Odrv4 I__5523 (
            .O(N__35036),
            .I(\c0.FRAME_MATCHER_i_17 ));
    LocalMux I__5522 (
            .O(N__35033),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__5521 (
            .O(N__35030),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__5520 (
            .O(N__35023),
            .I(N__35020));
    LocalMux I__5519 (
            .O(N__35020),
            .I(N__35017));
    Odrv12 I__5518 (
            .O(N__35017),
            .I(\c0.n44_adj_3255 ));
    InMux I__5517 (
            .O(N__35014),
            .I(N__35009));
    InMux I__5516 (
            .O(N__35013),
            .I(N__35006));
    InMux I__5515 (
            .O(N__35012),
            .I(N__35003));
    LocalMux I__5514 (
            .O(N__35009),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__5513 (
            .O(N__35006),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__5512 (
            .O(N__35003),
            .I(\c0.FRAME_MATCHER_i_24 ));
    SRMux I__5511 (
            .O(N__34996),
            .I(N__34993));
    LocalMux I__5510 (
            .O(N__34993),
            .I(N__34990));
    Span4Mux_v I__5509 (
            .O(N__34990),
            .I(N__34987));
    Span4Mux_h I__5508 (
            .O(N__34987),
            .I(N__34984));
    Odrv4 I__5507 (
            .O(N__34984),
            .I(\c0.n6_adj_3174 ));
    InMux I__5506 (
            .O(N__34981),
            .I(N__34978));
    LocalMux I__5505 (
            .O(N__34978),
            .I(N__34975));
    Odrv12 I__5504 (
            .O(N__34975),
            .I(\c0.n21273 ));
    CascadeMux I__5503 (
            .O(N__34972),
            .I(\c0.n5_adj_3306_cascade_ ));
    CascadeMux I__5502 (
            .O(N__34969),
            .I(N__34966));
    InMux I__5501 (
            .O(N__34966),
            .I(N__34960));
    InMux I__5500 (
            .O(N__34965),
            .I(N__34960));
    LocalMux I__5499 (
            .O(N__34960),
            .I(\c0.n2_adj_3302 ));
    CascadeMux I__5498 (
            .O(N__34957),
            .I(\c0.n11433_cascade_ ));
    CascadeMux I__5497 (
            .O(N__34954),
            .I(\c0.n8_adj_3228_cascade_ ));
    InMux I__5496 (
            .O(N__34951),
            .I(N__34947));
    InMux I__5495 (
            .O(N__34950),
            .I(N__34944));
    LocalMux I__5494 (
            .O(N__34947),
            .I(N__34941));
    LocalMux I__5493 (
            .O(N__34944),
            .I(\c0.n2103 ));
    Odrv4 I__5492 (
            .O(N__34941),
            .I(\c0.n2103 ));
    CascadeMux I__5491 (
            .O(N__34936),
            .I(\c0.n2103_cascade_ ));
    InMux I__5490 (
            .O(N__34933),
            .I(N__34928));
    InMux I__5489 (
            .O(N__34932),
            .I(N__34925));
    InMux I__5488 (
            .O(N__34931),
            .I(N__34922));
    LocalMux I__5487 (
            .O(N__34928),
            .I(N__34919));
    LocalMux I__5486 (
            .O(N__34925),
            .I(N__34916));
    LocalMux I__5485 (
            .O(N__34922),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv12 I__5484 (
            .O(N__34919),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv4 I__5483 (
            .O(N__34916),
            .I(\c0.FRAME_MATCHER_state_29 ));
    CascadeMux I__5482 (
            .O(N__34909),
            .I(\c0.n41_adj_3258_cascade_ ));
    InMux I__5481 (
            .O(N__34906),
            .I(N__34903));
    LocalMux I__5480 (
            .O(N__34903),
            .I(\c0.n43_adj_3257 ));
    InMux I__5479 (
            .O(N__34900),
            .I(N__34897));
    LocalMux I__5478 (
            .O(N__34897),
            .I(N__34893));
    InMux I__5477 (
            .O(N__34896),
            .I(N__34889));
    Span4Mux_v I__5476 (
            .O(N__34893),
            .I(N__34886));
    InMux I__5475 (
            .O(N__34892),
            .I(N__34883));
    LocalMux I__5474 (
            .O(N__34889),
            .I(N__34878));
    Span4Mux_v I__5473 (
            .O(N__34886),
            .I(N__34878));
    LocalMux I__5472 (
            .O(N__34883),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv4 I__5471 (
            .O(N__34878),
            .I(\c0.FRAME_MATCHER_i_10 ));
    InMux I__5470 (
            .O(N__34873),
            .I(N__34870));
    LocalMux I__5469 (
            .O(N__34870),
            .I(N__34865));
    InMux I__5468 (
            .O(N__34869),
            .I(N__34862));
    InMux I__5467 (
            .O(N__34868),
            .I(N__34859));
    Span4Mux_v I__5466 (
            .O(N__34865),
            .I(N__34856));
    LocalMux I__5465 (
            .O(N__34862),
            .I(\c0.FRAME_MATCHER_i_15 ));
    LocalMux I__5464 (
            .O(N__34859),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__5463 (
            .O(N__34856),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__5462 (
            .O(N__34849),
            .I(N__34845));
    InMux I__5461 (
            .O(N__34848),
            .I(N__34842));
    LocalMux I__5460 (
            .O(N__34845),
            .I(N__34839));
    LocalMux I__5459 (
            .O(N__34842),
            .I(N__34836));
    Span4Mux_v I__5458 (
            .O(N__34839),
            .I(N__34832));
    Span4Mux_v I__5457 (
            .O(N__34836),
            .I(N__34829));
    InMux I__5456 (
            .O(N__34835),
            .I(N__34826));
    Span4Mux_v I__5455 (
            .O(N__34832),
            .I(N__34823));
    Odrv4 I__5454 (
            .O(N__34829),
            .I(\c0.FRAME_MATCHER_i_13 ));
    LocalMux I__5453 (
            .O(N__34826),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__5452 (
            .O(N__34823),
            .I(\c0.FRAME_MATCHER_i_13 ));
    InMux I__5451 (
            .O(N__34816),
            .I(N__34813));
    LocalMux I__5450 (
            .O(N__34813),
            .I(N__34810));
    Span4Mux_v I__5449 (
            .O(N__34810),
            .I(N__34806));
    InMux I__5448 (
            .O(N__34809),
            .I(N__34803));
    Span4Mux_v I__5447 (
            .O(N__34806),
            .I(N__34799));
    LocalMux I__5446 (
            .O(N__34803),
            .I(N__34796));
    InMux I__5445 (
            .O(N__34802),
            .I(N__34793));
    Span4Mux_v I__5444 (
            .O(N__34799),
            .I(N__34790));
    Odrv4 I__5443 (
            .O(N__34796),
            .I(\c0.FRAME_MATCHER_i_9 ));
    LocalMux I__5442 (
            .O(N__34793),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv4 I__5441 (
            .O(N__34790),
            .I(\c0.FRAME_MATCHER_i_9 ));
    InMux I__5440 (
            .O(N__34783),
            .I(N__34780));
    LocalMux I__5439 (
            .O(N__34780),
            .I(\c0.n40_adj_3259 ));
    InMux I__5438 (
            .O(N__34777),
            .I(N__34774));
    LocalMux I__5437 (
            .O(N__34774),
            .I(\c0.n45_adj_3262 ));
    CascadeMux I__5436 (
            .O(N__34771),
            .I(\c0.n39_adj_3260_cascade_ ));
    InMux I__5435 (
            .O(N__34768),
            .I(N__34765));
    LocalMux I__5434 (
            .O(N__34765),
            .I(\c0.n50_adj_3261 ));
    InMux I__5433 (
            .O(N__34762),
            .I(N__34759));
    LocalMux I__5432 (
            .O(N__34759),
            .I(N__34754));
    InMux I__5431 (
            .O(N__34758),
            .I(N__34749));
    InMux I__5430 (
            .O(N__34757),
            .I(N__34749));
    Odrv4 I__5429 (
            .O(N__34754),
            .I(\c0.n11432 ));
    LocalMux I__5428 (
            .O(N__34749),
            .I(\c0.n11432 ));
    CascadeMux I__5427 (
            .O(N__34744),
            .I(\c0.n14_adj_3080_cascade_ ));
    InMux I__5426 (
            .O(N__34741),
            .I(N__34738));
    LocalMux I__5425 (
            .O(N__34738),
            .I(N__34735));
    Span4Mux_h I__5424 (
            .O(N__34735),
            .I(N__34732));
    Odrv4 I__5423 (
            .O(N__34732),
            .I(\c0.n10_adj_3081 ));
    CascadeMux I__5422 (
            .O(N__34729),
            .I(N__34724));
    InMux I__5421 (
            .O(N__34728),
            .I(N__34721));
    InMux I__5420 (
            .O(N__34727),
            .I(N__34718));
    InMux I__5419 (
            .O(N__34724),
            .I(N__34715));
    LocalMux I__5418 (
            .O(N__34721),
            .I(N__34712));
    LocalMux I__5417 (
            .O(N__34718),
            .I(N__34707));
    LocalMux I__5416 (
            .O(N__34715),
            .I(N__34707));
    Span4Mux_h I__5415 (
            .O(N__34712),
            .I(N__34704));
    Odrv4 I__5414 (
            .O(N__34707),
            .I(\c0.n4812 ));
    Odrv4 I__5413 (
            .O(N__34704),
            .I(\c0.n4812 ));
    InMux I__5412 (
            .O(N__34699),
            .I(N__34696));
    LocalMux I__5411 (
            .O(N__34696),
            .I(\c0.n19119 ));
    CascadeMux I__5410 (
            .O(N__34693),
            .I(\c0.n19119_cascade_ ));
    CascadeMux I__5409 (
            .O(N__34690),
            .I(N__34680));
    CascadeMux I__5408 (
            .O(N__34689),
            .I(N__34677));
    CascadeMux I__5407 (
            .O(N__34688),
            .I(N__34674));
    CascadeMux I__5406 (
            .O(N__34687),
            .I(N__34671));
    CascadeMux I__5405 (
            .O(N__34686),
            .I(N__34668));
    CascadeMux I__5404 (
            .O(N__34685),
            .I(N__34665));
    CascadeMux I__5403 (
            .O(N__34684),
            .I(N__34662));
    CascadeMux I__5402 (
            .O(N__34683),
            .I(N__34659));
    InMux I__5401 (
            .O(N__34680),
            .I(N__34650));
    InMux I__5400 (
            .O(N__34677),
            .I(N__34650));
    InMux I__5399 (
            .O(N__34674),
            .I(N__34650));
    InMux I__5398 (
            .O(N__34671),
            .I(N__34650));
    InMux I__5397 (
            .O(N__34668),
            .I(N__34641));
    InMux I__5396 (
            .O(N__34665),
            .I(N__34641));
    InMux I__5395 (
            .O(N__34662),
            .I(N__34641));
    InMux I__5394 (
            .O(N__34659),
            .I(N__34641));
    LocalMux I__5393 (
            .O(N__34650),
            .I(\c0.rx.n3 ));
    LocalMux I__5392 (
            .O(N__34641),
            .I(\c0.rx.n3 ));
    InMux I__5391 (
            .O(N__34636),
            .I(\c0.rx.n17273 ));
    InMux I__5390 (
            .O(N__34633),
            .I(N__34630));
    LocalMux I__5389 (
            .O(N__34630),
            .I(\c0.rx.n7 ));
    CascadeMux I__5388 (
            .O(N__34627),
            .I(N__34624));
    InMux I__5387 (
            .O(N__34624),
            .I(N__34621));
    LocalMux I__5386 (
            .O(N__34621),
            .I(N__34618));
    Span4Mux_v I__5385 (
            .O(N__34618),
            .I(N__34615));
    Span4Mux_v I__5384 (
            .O(N__34615),
            .I(N__34611));
    InMux I__5383 (
            .O(N__34614),
            .I(N__34607));
    Span4Mux_v I__5382 (
            .O(N__34611),
            .I(N__34604));
    InMux I__5381 (
            .O(N__34610),
            .I(N__34601));
    LocalMux I__5380 (
            .O(N__34607),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv4 I__5379 (
            .O(N__34604),
            .I(\c0.FRAME_MATCHER_i_8 ));
    LocalMux I__5378 (
            .O(N__34601),
            .I(\c0.FRAME_MATCHER_i_8 ));
    InMux I__5377 (
            .O(N__34594),
            .I(N__34591));
    LocalMux I__5376 (
            .O(N__34591),
            .I(N__34586));
    InMux I__5375 (
            .O(N__34590),
            .I(N__34583));
    InMux I__5374 (
            .O(N__34589),
            .I(N__34580));
    Odrv4 I__5373 (
            .O(N__34586),
            .I(\c0.FRAME_MATCHER_i_19 ));
    LocalMux I__5372 (
            .O(N__34583),
            .I(\c0.FRAME_MATCHER_i_19 ));
    LocalMux I__5371 (
            .O(N__34580),
            .I(\c0.FRAME_MATCHER_i_19 ));
    SRMux I__5370 (
            .O(N__34573),
            .I(N__34570));
    LocalMux I__5369 (
            .O(N__34570),
            .I(N__34567));
    Span4Mux_h I__5368 (
            .O(N__34567),
            .I(N__34564));
    Span4Mux_v I__5367 (
            .O(N__34564),
            .I(N__34561));
    Odrv4 I__5366 (
            .O(N__34561),
            .I(\c0.n6_adj_3161 ));
    InMux I__5365 (
            .O(N__34558),
            .I(N__34552));
    InMux I__5364 (
            .O(N__34557),
            .I(N__34552));
    LocalMux I__5363 (
            .O(N__34552),
            .I(N__34548));
    InMux I__5362 (
            .O(N__34551),
            .I(N__34545));
    Span4Mux_v I__5361 (
            .O(N__34548),
            .I(N__34542));
    LocalMux I__5360 (
            .O(N__34545),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__5359 (
            .O(N__34542),
            .I(\c0.FRAME_MATCHER_i_25 ));
    SRMux I__5358 (
            .O(N__34537),
            .I(N__34534));
    LocalMux I__5357 (
            .O(N__34534),
            .I(N__34531));
    Span4Mux_v I__5356 (
            .O(N__34531),
            .I(N__34528));
    Span4Mux_v I__5355 (
            .O(N__34528),
            .I(N__34525));
    Odrv4 I__5354 (
            .O(N__34525),
            .I(\c0.n6_adj_3172 ));
    SRMux I__5353 (
            .O(N__34522),
            .I(N__34519));
    LocalMux I__5352 (
            .O(N__34519),
            .I(N__34516));
    Span4Mux_h I__5351 (
            .O(N__34516),
            .I(N__34513));
    Span4Mux_v I__5350 (
            .O(N__34513),
            .I(N__34510));
    Odrv4 I__5349 (
            .O(N__34510),
            .I(\c0.n6_adj_3194 ));
    InMux I__5348 (
            .O(N__34507),
            .I(N__34501));
    InMux I__5347 (
            .O(N__34506),
            .I(N__34501));
    LocalMux I__5346 (
            .O(N__34501),
            .I(N__34498));
    Span4Mux_v I__5345 (
            .O(N__34498),
            .I(N__34494));
    InMux I__5344 (
            .O(N__34497),
            .I(N__34491));
    Span4Mux_v I__5343 (
            .O(N__34494),
            .I(N__34488));
    LocalMux I__5342 (
            .O(N__34491),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv4 I__5341 (
            .O(N__34488),
            .I(\c0.FRAME_MATCHER_i_12 ));
    InMux I__5340 (
            .O(N__34483),
            .I(N__34478));
    InMux I__5339 (
            .O(N__34482),
            .I(N__34475));
    InMux I__5338 (
            .O(N__34481),
            .I(N__34472));
    LocalMux I__5337 (
            .O(N__34478),
            .I(\c0.FRAME_MATCHER_i_20 ));
    LocalMux I__5336 (
            .O(N__34475),
            .I(\c0.FRAME_MATCHER_i_20 ));
    LocalMux I__5335 (
            .O(N__34472),
            .I(\c0.FRAME_MATCHER_i_20 ));
    CascadeMux I__5334 (
            .O(N__34465),
            .I(N__34461));
    InMux I__5333 (
            .O(N__34464),
            .I(N__34456));
    InMux I__5332 (
            .O(N__34461),
            .I(N__34456));
    LocalMux I__5331 (
            .O(N__34456),
            .I(N__34452));
    InMux I__5330 (
            .O(N__34455),
            .I(N__34449));
    Span4Mux_v I__5329 (
            .O(N__34452),
            .I(N__34446));
    LocalMux I__5328 (
            .O(N__34449),
            .I(\c0.FRAME_MATCHER_i_14 ));
    Odrv4 I__5327 (
            .O(N__34446),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__5326 (
            .O(N__34441),
            .I(N__34437));
    InMux I__5325 (
            .O(N__34440),
            .I(N__34434));
    LocalMux I__5324 (
            .O(N__34437),
            .I(N__34431));
    LocalMux I__5323 (
            .O(N__34434),
            .I(N__34428));
    Span4Mux_v I__5322 (
            .O(N__34431),
            .I(N__34425));
    Span12Mux_h I__5321 (
            .O(N__34428),
            .I(N__34421));
    Span4Mux_v I__5320 (
            .O(N__34425),
            .I(N__34418));
    InMux I__5319 (
            .O(N__34424),
            .I(N__34415));
    Span12Mux_v I__5318 (
            .O(N__34421),
            .I(N__34412));
    Odrv4 I__5317 (
            .O(N__34418),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__5316 (
            .O(N__34415),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv12 I__5315 (
            .O(N__34412),
            .I(\c0.FRAME_MATCHER_i_7 ));
    SRMux I__5314 (
            .O(N__34405),
            .I(N__34402));
    LocalMux I__5313 (
            .O(N__34402),
            .I(N__34399));
    Span4Mux_v I__5312 (
            .O(N__34399),
            .I(N__34396));
    Span4Mux_v I__5311 (
            .O(N__34396),
            .I(N__34393));
    Odrv4 I__5310 (
            .O(N__34393),
            .I(\c0.n6_adj_3160 ));
    InMux I__5309 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__5308 (
            .O(N__34387),
            .I(N__34383));
    InMux I__5307 (
            .O(N__34386),
            .I(N__34379));
    Span4Mux_h I__5306 (
            .O(N__34383),
            .I(N__34376));
    InMux I__5305 (
            .O(N__34382),
            .I(N__34373));
    LocalMux I__5304 (
            .O(N__34379),
            .I(N__34370));
    Odrv4 I__5303 (
            .O(N__34376),
            .I(\c0.FRAME_MATCHER_i_22 ));
    LocalMux I__5302 (
            .O(N__34373),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__5301 (
            .O(N__34370),
            .I(\c0.FRAME_MATCHER_i_22 ));
    CascadeMux I__5300 (
            .O(N__34363),
            .I(N__34360));
    InMux I__5299 (
            .O(N__34360),
            .I(N__34357));
    LocalMux I__5298 (
            .O(N__34357),
            .I(N__34352));
    InMux I__5297 (
            .O(N__34356),
            .I(N__34349));
    InMux I__5296 (
            .O(N__34355),
            .I(N__34346));
    Span4Mux_v I__5295 (
            .O(N__34352),
            .I(N__34343));
    LocalMux I__5294 (
            .O(N__34349),
            .I(\c0.FRAME_MATCHER_i_16 ));
    LocalMux I__5293 (
            .O(N__34346),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__5292 (
            .O(N__34343),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__5291 (
            .O(N__34336),
            .I(N__34332));
    InMux I__5290 (
            .O(N__34335),
            .I(N__34329));
    LocalMux I__5289 (
            .O(N__34332),
            .I(N__34324));
    LocalMux I__5288 (
            .O(N__34329),
            .I(N__34324));
    Span4Mux_v I__5287 (
            .O(N__34324),
            .I(N__34320));
    InMux I__5286 (
            .O(N__34323),
            .I(N__34317));
    Span4Mux_v I__5285 (
            .O(N__34320),
            .I(N__34314));
    LocalMux I__5284 (
            .O(N__34317),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv4 I__5283 (
            .O(N__34314),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__5282 (
            .O(N__34309),
            .I(N__34306));
    LocalMux I__5281 (
            .O(N__34306),
            .I(n13179));
    InMux I__5280 (
            .O(N__34303),
            .I(bfn_15_19_0_));
    InMux I__5279 (
            .O(N__34300),
            .I(\c0.rx.n17267 ));
    InMux I__5278 (
            .O(N__34297),
            .I(N__34294));
    LocalMux I__5277 (
            .O(N__34294),
            .I(n12908));
    InMux I__5276 (
            .O(N__34291),
            .I(\c0.rx.n17268 ));
    InMux I__5275 (
            .O(N__34288),
            .I(\c0.rx.n17269 ));
    InMux I__5274 (
            .O(N__34285),
            .I(\c0.rx.n17270 ));
    InMux I__5273 (
            .O(N__34282),
            .I(\c0.rx.n17271 ));
    InMux I__5272 (
            .O(N__34279),
            .I(\c0.rx.n17272 ));
    CascadeMux I__5271 (
            .O(N__34276),
            .I(\c0.rx.n14601_cascade_ ));
    InMux I__5270 (
            .O(N__34273),
            .I(N__34270));
    LocalMux I__5269 (
            .O(N__34270),
            .I(N__34267));
    Odrv12 I__5268 (
            .O(N__34267),
            .I(n12301));
    InMux I__5267 (
            .O(N__34264),
            .I(N__34261));
    LocalMux I__5266 (
            .O(N__34261),
            .I(N__34258));
    Span4Mux_h I__5265 (
            .O(N__34258),
            .I(N__34255));
    Odrv4 I__5264 (
            .O(N__34255),
            .I(\c0.n15685 ));
    CascadeMux I__5263 (
            .O(N__34252),
            .I(N__34249));
    InMux I__5262 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__5261 (
            .O(N__34246),
            .I(N__34243));
    Span4Mux_h I__5260 (
            .O(N__34243),
            .I(N__34240));
    Odrv4 I__5259 (
            .O(N__34240),
            .I(\c0.rx.n6 ));
    CascadeMux I__5258 (
            .O(N__34237),
            .I(n12492_cascade_));
    InMux I__5257 (
            .O(N__34234),
            .I(N__34230));
    CascadeMux I__5256 (
            .O(N__34233),
            .I(N__34223));
    LocalMux I__5255 (
            .O(N__34230),
            .I(N__34217));
    InMux I__5254 (
            .O(N__34229),
            .I(N__34212));
    InMux I__5253 (
            .O(N__34228),
            .I(N__34212));
    InMux I__5252 (
            .O(N__34227),
            .I(N__34209));
    InMux I__5251 (
            .O(N__34226),
            .I(N__34204));
    InMux I__5250 (
            .O(N__34223),
            .I(N__34204));
    InMux I__5249 (
            .O(N__34222),
            .I(N__34197));
    InMux I__5248 (
            .O(N__34221),
            .I(N__34197));
    InMux I__5247 (
            .O(N__34220),
            .I(N__34197));
    Span4Mux_v I__5246 (
            .O(N__34217),
            .I(N__34194));
    LocalMux I__5245 (
            .O(N__34212),
            .I(\c0.r_Bit_Index_0 ));
    LocalMux I__5244 (
            .O(N__34209),
            .I(\c0.r_Bit_Index_0 ));
    LocalMux I__5243 (
            .O(N__34204),
            .I(\c0.r_Bit_Index_0 ));
    LocalMux I__5242 (
            .O(N__34197),
            .I(\c0.r_Bit_Index_0 ));
    Odrv4 I__5241 (
            .O(N__34194),
            .I(\c0.r_Bit_Index_0 ));
    IoInMux I__5240 (
            .O(N__34183),
            .I(N__34179));
    InMux I__5239 (
            .O(N__34182),
            .I(N__34176));
    LocalMux I__5238 (
            .O(N__34179),
            .I(N__34170));
    LocalMux I__5237 (
            .O(N__34176),
            .I(N__34170));
    InMux I__5236 (
            .O(N__34175),
            .I(N__34165));
    Span4Mux_s3_h I__5235 (
            .O(N__34170),
            .I(N__34162));
    InMux I__5234 (
            .O(N__34169),
            .I(N__34155));
    InMux I__5233 (
            .O(N__34168),
            .I(N__34155));
    LocalMux I__5232 (
            .O(N__34165),
            .I(N__34152));
    Sp12to4 I__5231 (
            .O(N__34162),
            .I(N__34149));
    InMux I__5230 (
            .O(N__34161),
            .I(N__34146));
    InMux I__5229 (
            .O(N__34160),
            .I(N__34143));
    LocalMux I__5228 (
            .O(N__34155),
            .I(N__34138));
    Span4Mux_h I__5227 (
            .O(N__34152),
            .I(N__34138));
    Span12Mux_v I__5226 (
            .O(N__34149),
            .I(N__34135));
    LocalMux I__5225 (
            .O(N__34146),
            .I(N__34130));
    LocalMux I__5224 (
            .O(N__34143),
            .I(N__34130));
    Span4Mux_h I__5223 (
            .O(N__34138),
            .I(N__34127));
    Odrv12 I__5222 (
            .O(N__34135),
            .I(tx_o));
    Odrv4 I__5221 (
            .O(N__34130),
            .I(tx_o));
    Odrv4 I__5220 (
            .O(N__34127),
            .I(tx_o));
    CascadeMux I__5219 (
            .O(N__34120),
            .I(N__34116));
    CascadeMux I__5218 (
            .O(N__34119),
            .I(N__34113));
    InMux I__5217 (
            .O(N__34116),
            .I(N__34110));
    InMux I__5216 (
            .O(N__34113),
            .I(N__34107));
    LocalMux I__5215 (
            .O(N__34110),
            .I(N__34104));
    LocalMux I__5214 (
            .O(N__34107),
            .I(r_Tx_Data_1));
    Odrv4 I__5213 (
            .O(N__34104),
            .I(r_Tx_Data_1));
    InMux I__5212 (
            .O(N__34099),
            .I(N__34089));
    InMux I__5211 (
            .O(N__34098),
            .I(N__34086));
    InMux I__5210 (
            .O(N__34097),
            .I(N__34078));
    InMux I__5209 (
            .O(N__34096),
            .I(N__34078));
    InMux I__5208 (
            .O(N__34095),
            .I(N__34069));
    InMux I__5207 (
            .O(N__34094),
            .I(N__34069));
    InMux I__5206 (
            .O(N__34093),
            .I(N__34069));
    InMux I__5205 (
            .O(N__34092),
            .I(N__34069));
    LocalMux I__5204 (
            .O(N__34089),
            .I(N__34066));
    LocalMux I__5203 (
            .O(N__34086),
            .I(N__34056));
    InMux I__5202 (
            .O(N__34085),
            .I(N__34053));
    InMux I__5201 (
            .O(N__34084),
            .I(N__34050));
    InMux I__5200 (
            .O(N__34083),
            .I(N__34047));
    LocalMux I__5199 (
            .O(N__34078),
            .I(N__34040));
    LocalMux I__5198 (
            .O(N__34069),
            .I(N__34040));
    Span4Mux_h I__5197 (
            .O(N__34066),
            .I(N__34040));
    InMux I__5196 (
            .O(N__34065),
            .I(N__34037));
    InMux I__5195 (
            .O(N__34064),
            .I(N__34034));
    InMux I__5194 (
            .O(N__34063),
            .I(N__34031));
    InMux I__5193 (
            .O(N__34062),
            .I(N__34028));
    InMux I__5192 (
            .O(N__34061),
            .I(N__34021));
    InMux I__5191 (
            .O(N__34060),
            .I(N__34021));
    InMux I__5190 (
            .O(N__34059),
            .I(N__34021));
    Span4Mux_h I__5189 (
            .O(N__34056),
            .I(N__34018));
    LocalMux I__5188 (
            .O(N__34053),
            .I(N__34011));
    LocalMux I__5187 (
            .O(N__34050),
            .I(N__34011));
    LocalMux I__5186 (
            .O(N__34047),
            .I(N__34011));
    Span4Mux_h I__5185 (
            .O(N__34040),
            .I(N__34008));
    LocalMux I__5184 (
            .O(N__34037),
            .I(\c0.r_SM_Main_2 ));
    LocalMux I__5183 (
            .O(N__34034),
            .I(\c0.r_SM_Main_2 ));
    LocalMux I__5182 (
            .O(N__34031),
            .I(\c0.r_SM_Main_2 ));
    LocalMux I__5181 (
            .O(N__34028),
            .I(\c0.r_SM_Main_2 ));
    LocalMux I__5180 (
            .O(N__34021),
            .I(\c0.r_SM_Main_2 ));
    Odrv4 I__5179 (
            .O(N__34018),
            .I(\c0.r_SM_Main_2 ));
    Odrv4 I__5178 (
            .O(N__34011),
            .I(\c0.r_SM_Main_2 ));
    Odrv4 I__5177 (
            .O(N__34008),
            .I(\c0.r_SM_Main_2 ));
    InMux I__5176 (
            .O(N__33991),
            .I(N__33988));
    LocalMux I__5175 (
            .O(N__33988),
            .I(N__33985));
    Span4Mux_v I__5174 (
            .O(N__33985),
            .I(N__33982));
    Odrv4 I__5173 (
            .O(N__33982),
            .I(\c0.n21611 ));
    InMux I__5172 (
            .O(N__33979),
            .I(N__33976));
    LocalMux I__5171 (
            .O(N__33976),
            .I(N__33973));
    Span4Mux_h I__5170 (
            .O(N__33973),
            .I(N__33970));
    Span4Mux_h I__5169 (
            .O(N__33970),
            .I(N__33966));
    CascadeMux I__5168 (
            .O(N__33969),
            .I(N__33962));
    Span4Mux_v I__5167 (
            .O(N__33966),
            .I(N__33959));
    InMux I__5166 (
            .O(N__33965),
            .I(N__33956));
    InMux I__5165 (
            .O(N__33962),
            .I(N__33953));
    Odrv4 I__5164 (
            .O(N__33959),
            .I(encoder0_position_23));
    LocalMux I__5163 (
            .O(N__33956),
            .I(encoder0_position_23));
    LocalMux I__5162 (
            .O(N__33953),
            .I(encoder0_position_23));
    InMux I__5161 (
            .O(N__33946),
            .I(N__33942));
    InMux I__5160 (
            .O(N__33945),
            .I(N__33939));
    LocalMux I__5159 (
            .O(N__33942),
            .I(N__33936));
    LocalMux I__5158 (
            .O(N__33939),
            .I(data_out_frame_7_7));
    Odrv12 I__5157 (
            .O(N__33936),
            .I(data_out_frame_7_7));
    InMux I__5156 (
            .O(N__33931),
            .I(N__33927));
    InMux I__5155 (
            .O(N__33930),
            .I(N__33924));
    LocalMux I__5154 (
            .O(N__33927),
            .I(N__33921));
    LocalMux I__5153 (
            .O(N__33924),
            .I(r_Tx_Data_7));
    Odrv4 I__5152 (
            .O(N__33921),
            .I(r_Tx_Data_7));
    InMux I__5151 (
            .O(N__33916),
            .I(N__33910));
    InMux I__5150 (
            .O(N__33915),
            .I(N__33910));
    LocalMux I__5149 (
            .O(N__33910),
            .I(data_out_frame_7_5));
    InMux I__5148 (
            .O(N__33907),
            .I(N__33903));
    InMux I__5147 (
            .O(N__33906),
            .I(N__33900));
    LocalMux I__5146 (
            .O(N__33903),
            .I(N__33897));
    LocalMux I__5145 (
            .O(N__33900),
            .I(data_out_frame_6_5));
    Odrv4 I__5144 (
            .O(N__33897),
            .I(data_out_frame_6_5));
    InMux I__5143 (
            .O(N__33892),
            .I(N__33889));
    LocalMux I__5142 (
            .O(N__33889),
            .I(\c0.n5_adj_3447 ));
    CascadeMux I__5141 (
            .O(N__33886),
            .I(N__33882));
    CascadeMux I__5140 (
            .O(N__33885),
            .I(N__33874));
    InMux I__5139 (
            .O(N__33882),
            .I(N__33870));
    InMux I__5138 (
            .O(N__33881),
            .I(N__33865));
    InMux I__5137 (
            .O(N__33880),
            .I(N__33865));
    InMux I__5136 (
            .O(N__33879),
            .I(N__33862));
    CascadeMux I__5135 (
            .O(N__33878),
            .I(N__33858));
    CascadeMux I__5134 (
            .O(N__33877),
            .I(N__33855));
    InMux I__5133 (
            .O(N__33874),
            .I(N__33852));
    InMux I__5132 (
            .O(N__33873),
            .I(N__33849));
    LocalMux I__5131 (
            .O(N__33870),
            .I(N__33845));
    LocalMux I__5130 (
            .O(N__33865),
            .I(N__33840));
    LocalMux I__5129 (
            .O(N__33862),
            .I(N__33840));
    InMux I__5128 (
            .O(N__33861),
            .I(N__33835));
    InMux I__5127 (
            .O(N__33858),
            .I(N__33835));
    InMux I__5126 (
            .O(N__33855),
            .I(N__33832));
    LocalMux I__5125 (
            .O(N__33852),
            .I(N__33827));
    LocalMux I__5124 (
            .O(N__33849),
            .I(N__33827));
    InMux I__5123 (
            .O(N__33848),
            .I(N__33824));
    Span4Mux_h I__5122 (
            .O(N__33845),
            .I(N__33821));
    Span4Mux_v I__5121 (
            .O(N__33840),
            .I(N__33818));
    LocalMux I__5120 (
            .O(N__33835),
            .I(byte_transmit_counter_5));
    LocalMux I__5119 (
            .O(N__33832),
            .I(byte_transmit_counter_5));
    Odrv12 I__5118 (
            .O(N__33827),
            .I(byte_transmit_counter_5));
    LocalMux I__5117 (
            .O(N__33824),
            .I(byte_transmit_counter_5));
    Odrv4 I__5116 (
            .O(N__33821),
            .I(byte_transmit_counter_5));
    Odrv4 I__5115 (
            .O(N__33818),
            .I(byte_transmit_counter_5));
    CascadeMux I__5114 (
            .O(N__33805),
            .I(N__33802));
    InMux I__5113 (
            .O(N__33802),
            .I(N__33792));
    InMux I__5112 (
            .O(N__33801),
            .I(N__33792));
    InMux I__5111 (
            .O(N__33800),
            .I(N__33789));
    InMux I__5110 (
            .O(N__33799),
            .I(N__33786));
    InMux I__5109 (
            .O(N__33798),
            .I(N__33780));
    InMux I__5108 (
            .O(N__33797),
            .I(N__33780));
    LocalMux I__5107 (
            .O(N__33792),
            .I(N__33775));
    LocalMux I__5106 (
            .O(N__33789),
            .I(N__33775));
    LocalMux I__5105 (
            .O(N__33786),
            .I(N__33772));
    InMux I__5104 (
            .O(N__33785),
            .I(N__33769));
    LocalMux I__5103 (
            .O(N__33780),
            .I(N__33766));
    Span4Mux_h I__5102 (
            .O(N__33775),
            .I(N__33762));
    Span4Mux_h I__5101 (
            .O(N__33772),
            .I(N__33757));
    LocalMux I__5100 (
            .O(N__33769),
            .I(N__33757));
    Span4Mux_h I__5099 (
            .O(N__33766),
            .I(N__33754));
    InMux I__5098 (
            .O(N__33765),
            .I(N__33751));
    Odrv4 I__5097 (
            .O(N__33762),
            .I(n9377));
    Odrv4 I__5096 (
            .O(N__33757),
            .I(n9377));
    Odrv4 I__5095 (
            .O(N__33754),
            .I(n9377));
    LocalMux I__5094 (
            .O(N__33751),
            .I(n9377));
    CascadeMux I__5093 (
            .O(N__33742),
            .I(N__33739));
    InMux I__5092 (
            .O(N__33739),
            .I(N__33736));
    LocalMux I__5091 (
            .O(N__33736),
            .I(N__33732));
    InMux I__5090 (
            .O(N__33735),
            .I(N__33729));
    Span4Mux_v I__5089 (
            .O(N__33732),
            .I(N__33726));
    LocalMux I__5088 (
            .O(N__33729),
            .I(data_out_frame_5_5));
    Odrv4 I__5087 (
            .O(N__33726),
            .I(data_out_frame_5_5));
    CascadeMux I__5086 (
            .O(N__33721),
            .I(N__33718));
    InMux I__5085 (
            .O(N__33718),
            .I(N__33715));
    LocalMux I__5084 (
            .O(N__33715),
            .I(\c0.n21546 ));
    SRMux I__5083 (
            .O(N__33712),
            .I(N__33709));
    LocalMux I__5082 (
            .O(N__33709),
            .I(N__33706));
    Odrv4 I__5081 (
            .O(N__33706),
            .I(\c0.n6_adj_3192 ));
    InMux I__5080 (
            .O(N__33703),
            .I(N__33699));
    CascadeMux I__5079 (
            .O(N__33702),
            .I(N__33696));
    LocalMux I__5078 (
            .O(N__33699),
            .I(N__33693));
    InMux I__5077 (
            .O(N__33696),
            .I(N__33690));
    Span4Mux_h I__5076 (
            .O(N__33693),
            .I(N__33686));
    LocalMux I__5075 (
            .O(N__33690),
            .I(N__33683));
    InMux I__5074 (
            .O(N__33689),
            .I(N__33680));
    Span4Mux_v I__5073 (
            .O(N__33686),
            .I(N__33675));
    Span4Mux_h I__5072 (
            .O(N__33683),
            .I(N__33675));
    LocalMux I__5071 (
            .O(N__33680),
            .I(encoder1_position_1));
    Odrv4 I__5070 (
            .O(N__33675),
            .I(encoder1_position_1));
    InMux I__5069 (
            .O(N__33670),
            .I(N__33666));
    InMux I__5068 (
            .O(N__33669),
            .I(N__33663));
    LocalMux I__5067 (
            .O(N__33666),
            .I(N__33660));
    LocalMux I__5066 (
            .O(N__33663),
            .I(data_out_frame_13_1));
    Odrv4 I__5065 (
            .O(N__33660),
            .I(data_out_frame_13_1));
    SRMux I__5064 (
            .O(N__33655),
            .I(N__33652));
    LocalMux I__5063 (
            .O(N__33652),
            .I(N__33649));
    Odrv4 I__5062 (
            .O(N__33649),
            .I(\c0.n6_adj_3190 ));
    CascadeMux I__5061 (
            .O(N__33646),
            .I(N__33643));
    InMux I__5060 (
            .O(N__33643),
            .I(N__33639));
    InMux I__5059 (
            .O(N__33642),
            .I(N__33636));
    LocalMux I__5058 (
            .O(N__33639),
            .I(N__33633));
    LocalMux I__5057 (
            .O(N__33636),
            .I(data_out_frame_11_2));
    Odrv12 I__5056 (
            .O(N__33633),
            .I(data_out_frame_11_2));
    InMux I__5055 (
            .O(N__33628),
            .I(N__33624));
    InMux I__5054 (
            .O(N__33627),
            .I(N__33621));
    LocalMux I__5053 (
            .O(N__33624),
            .I(N__33616));
    LocalMux I__5052 (
            .O(N__33621),
            .I(N__33616));
    Odrv4 I__5051 (
            .O(N__33616),
            .I(data_out_frame_10_0));
    CascadeMux I__5050 (
            .O(N__33613),
            .I(N__33610));
    InMux I__5049 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__5048 (
            .O(N__33607),
            .I(N__33603));
    InMux I__5047 (
            .O(N__33606),
            .I(N__33600));
    Span12Mux_h I__5046 (
            .O(N__33603),
            .I(N__33597));
    LocalMux I__5045 (
            .O(N__33600),
            .I(data_out_frame_11_0));
    Odrv12 I__5044 (
            .O(N__33597),
            .I(data_out_frame_11_0));
    InMux I__5043 (
            .O(N__33592),
            .I(N__33588));
    InMux I__5042 (
            .O(N__33591),
            .I(N__33585));
    LocalMux I__5041 (
            .O(N__33588),
            .I(N__33582));
    LocalMux I__5040 (
            .O(N__33585),
            .I(data_out_frame_8_0));
    Odrv4 I__5039 (
            .O(N__33582),
            .I(data_out_frame_8_0));
    CascadeMux I__5038 (
            .O(N__33577),
            .I(\c0.n21617_cascade_ ));
    InMux I__5037 (
            .O(N__33574),
            .I(N__33570));
    InMux I__5036 (
            .O(N__33573),
            .I(N__33567));
    LocalMux I__5035 (
            .O(N__33570),
            .I(N__33564));
    LocalMux I__5034 (
            .O(N__33567),
            .I(data_out_frame_9_0));
    Odrv12 I__5033 (
            .O(N__33564),
            .I(data_out_frame_9_0));
    CascadeMux I__5032 (
            .O(N__33559),
            .I(\c0.n21620_cascade_ ));
    InMux I__5031 (
            .O(N__33556),
            .I(N__33553));
    LocalMux I__5030 (
            .O(N__33553),
            .I(N__33550));
    Span4Mux_h I__5029 (
            .O(N__33550),
            .I(N__33547));
    Odrv4 I__5028 (
            .O(N__33547),
            .I(\c0.n21574 ));
    InMux I__5027 (
            .O(N__33544),
            .I(N__33541));
    LocalMux I__5026 (
            .O(N__33541),
            .I(N__33537));
    InMux I__5025 (
            .O(N__33540),
            .I(N__33534));
    Span4Mux_h I__5024 (
            .O(N__33537),
            .I(N__33531));
    LocalMux I__5023 (
            .O(N__33534),
            .I(\c0.byte_transmit_counter_6 ));
    Odrv4 I__5022 (
            .O(N__33531),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__5021 (
            .O(N__33526),
            .I(N__33523));
    LocalMux I__5020 (
            .O(N__33523),
            .I(N__33519));
    InMux I__5019 (
            .O(N__33522),
            .I(N__33516));
    Span4Mux_h I__5018 (
            .O(N__33519),
            .I(N__33513));
    LocalMux I__5017 (
            .O(N__33516),
            .I(\c0.byte_transmit_counter_7 ));
    Odrv4 I__5016 (
            .O(N__33513),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__5015 (
            .O(N__33508),
            .I(N__33502));
    InMux I__5014 (
            .O(N__33507),
            .I(N__33502));
    LocalMux I__5013 (
            .O(N__33502),
            .I(N__33499));
    Odrv12 I__5012 (
            .O(N__33499),
            .I(\c0.n7235 ));
    InMux I__5011 (
            .O(N__33496),
            .I(N__33493));
    LocalMux I__5010 (
            .O(N__33493),
            .I(N__33490));
    Span4Mux_v I__5009 (
            .O(N__33490),
            .I(N__33487));
    Span4Mux_v I__5008 (
            .O(N__33487),
            .I(N__33484));
    Odrv4 I__5007 (
            .O(N__33484),
            .I(\c0.n2_adj_3147 ));
    SRMux I__5006 (
            .O(N__33481),
            .I(N__33478));
    LocalMux I__5005 (
            .O(N__33478),
            .I(N__33475));
    Span4Mux_h I__5004 (
            .O(N__33475),
            .I(N__33472));
    Span4Mux_v I__5003 (
            .O(N__33472),
            .I(N__33469));
    Odrv4 I__5002 (
            .O(N__33469),
            .I(\c0.n6_adj_3151 ));
    InMux I__5001 (
            .O(N__33466),
            .I(N__33463));
    LocalMux I__5000 (
            .O(N__33463),
            .I(N__33459));
    CascadeMux I__4999 (
            .O(N__33462),
            .I(N__33455));
    Span12Mux_v I__4998 (
            .O(N__33459),
            .I(N__33452));
    InMux I__4997 (
            .O(N__33458),
            .I(N__33449));
    InMux I__4996 (
            .O(N__33455),
            .I(N__33446));
    Odrv12 I__4995 (
            .O(N__33452),
            .I(encoder0_position_21));
    LocalMux I__4994 (
            .O(N__33449),
            .I(encoder0_position_21));
    LocalMux I__4993 (
            .O(N__33446),
            .I(encoder0_position_21));
    InMux I__4992 (
            .O(N__33439),
            .I(N__33436));
    LocalMux I__4991 (
            .O(N__33436),
            .I(N__33433));
    Odrv4 I__4990 (
            .O(N__33433),
            .I(\c0.n21470 ));
    CascadeMux I__4989 (
            .O(N__33430),
            .I(N__33427));
    InMux I__4988 (
            .O(N__33427),
            .I(N__33424));
    LocalMux I__4987 (
            .O(N__33424),
            .I(N__33421));
    Span4Mux_v I__4986 (
            .O(N__33421),
            .I(N__33418));
    Span4Mux_h I__4985 (
            .O(N__33418),
            .I(N__33415));
    Odrv4 I__4984 (
            .O(N__33415),
            .I(\c0.n21542 ));
    InMux I__4983 (
            .O(N__33412),
            .I(N__33409));
    LocalMux I__4982 (
            .O(N__33409),
            .I(N__33406));
    Span4Mux_h I__4981 (
            .O(N__33406),
            .I(N__33403));
    Odrv4 I__4980 (
            .O(N__33403),
            .I(n2316));
    SRMux I__4979 (
            .O(N__33400),
            .I(N__33397));
    LocalMux I__4978 (
            .O(N__33397),
            .I(N__33394));
    Odrv4 I__4977 (
            .O(N__33394),
            .I(\c0.n6_adj_3156 ));
    CascadeMux I__4976 (
            .O(N__33391),
            .I(N__33388));
    InMux I__4975 (
            .O(N__33388),
            .I(N__33385));
    LocalMux I__4974 (
            .O(N__33385),
            .I(N__33380));
    InMux I__4973 (
            .O(N__33384),
            .I(N__33375));
    InMux I__4972 (
            .O(N__33383),
            .I(N__33375));
    Span4Mux_h I__4971 (
            .O(N__33380),
            .I(N__33372));
    LocalMux I__4970 (
            .O(N__33375),
            .I(encoder1_position_29));
    Odrv4 I__4969 (
            .O(N__33372),
            .I(encoder1_position_29));
    InMux I__4968 (
            .O(N__33367),
            .I(N__33363));
    InMux I__4967 (
            .O(N__33366),
            .I(N__33360));
    LocalMux I__4966 (
            .O(N__33363),
            .I(data_out_frame_10_5));
    LocalMux I__4965 (
            .O(N__33360),
            .I(data_out_frame_10_5));
    InMux I__4964 (
            .O(N__33355),
            .I(N__33351));
    CascadeMux I__4963 (
            .O(N__33354),
            .I(N__33347));
    LocalMux I__4962 (
            .O(N__33351),
            .I(N__33344));
    InMux I__4961 (
            .O(N__33350),
            .I(N__33341));
    InMux I__4960 (
            .O(N__33347),
            .I(N__33338));
    Span4Mux_h I__4959 (
            .O(N__33344),
            .I(N__33335));
    LocalMux I__4958 (
            .O(N__33341),
            .I(N__33330));
    LocalMux I__4957 (
            .O(N__33338),
            .I(N__33330));
    Odrv4 I__4956 (
            .O(N__33335),
            .I(encoder0_position_29));
    Odrv4 I__4955 (
            .O(N__33330),
            .I(encoder0_position_29));
    InMux I__4954 (
            .O(N__33325),
            .I(N__33322));
    LocalMux I__4953 (
            .O(N__33322),
            .I(N__33318));
    InMux I__4952 (
            .O(N__33321),
            .I(N__33315));
    Span4Mux_h I__4951 (
            .O(N__33318),
            .I(N__33312));
    LocalMux I__4950 (
            .O(N__33315),
            .I(\c0.data_out_frame_7_0 ));
    Odrv4 I__4949 (
            .O(N__33312),
            .I(\c0.data_out_frame_7_0 ));
    InMux I__4948 (
            .O(N__33307),
            .I(N__33304));
    LocalMux I__4947 (
            .O(N__33304),
            .I(N__33301));
    Span4Mux_v I__4946 (
            .O(N__33301),
            .I(N__33298));
    Odrv4 I__4945 (
            .O(N__33298),
            .I(\c0.n17150 ));
    InMux I__4944 (
            .O(N__33295),
            .I(N__33291));
    CascadeMux I__4943 (
            .O(N__33294),
            .I(N__33287));
    LocalMux I__4942 (
            .O(N__33291),
            .I(N__33284));
    InMux I__4941 (
            .O(N__33290),
            .I(N__33281));
    InMux I__4940 (
            .O(N__33287),
            .I(N__33278));
    Span4Mux_v I__4939 (
            .O(N__33284),
            .I(N__33275));
    LocalMux I__4938 (
            .O(N__33281),
            .I(N__33270));
    LocalMux I__4937 (
            .O(N__33278),
            .I(N__33270));
    Odrv4 I__4936 (
            .O(N__33275),
            .I(encoder1_position_18));
    Odrv4 I__4935 (
            .O(N__33270),
            .I(encoder1_position_18));
    InMux I__4934 (
            .O(N__33265),
            .I(N__33262));
    LocalMux I__4933 (
            .O(N__33262),
            .I(N__33259));
    Span4Mux_h I__4932 (
            .O(N__33259),
            .I(N__33254));
    CascadeMux I__4931 (
            .O(N__33258),
            .I(N__33251));
    InMux I__4930 (
            .O(N__33257),
            .I(N__33248));
    Span4Mux_h I__4929 (
            .O(N__33254),
            .I(N__33245));
    InMux I__4928 (
            .O(N__33251),
            .I(N__33242));
    LocalMux I__4927 (
            .O(N__33248),
            .I(encoder0_position_11));
    Odrv4 I__4926 (
            .O(N__33245),
            .I(encoder0_position_11));
    LocalMux I__4925 (
            .O(N__33242),
            .I(encoder0_position_11));
    InMux I__4924 (
            .O(N__33235),
            .I(N__33232));
    LocalMux I__4923 (
            .O(N__33232),
            .I(N__33228));
    InMux I__4922 (
            .O(N__33231),
            .I(N__33225));
    Span4Mux_h I__4921 (
            .O(N__33228),
            .I(N__33222));
    LocalMux I__4920 (
            .O(N__33225),
            .I(data_out_frame_10_7));
    Odrv4 I__4919 (
            .O(N__33222),
            .I(data_out_frame_10_7));
    InMux I__4918 (
            .O(N__33217),
            .I(N__33214));
    LocalMux I__4917 (
            .O(N__33214),
            .I(N__33211));
    Span4Mux_v I__4916 (
            .O(N__33211),
            .I(N__33208));
    Odrv4 I__4915 (
            .O(N__33208),
            .I(\c0.n21623 ));
    InMux I__4914 (
            .O(N__33205),
            .I(N__33201));
    InMux I__4913 (
            .O(N__33204),
            .I(N__33198));
    LocalMux I__4912 (
            .O(N__33201),
            .I(N__33195));
    LocalMux I__4911 (
            .O(N__33198),
            .I(data_out_frame_9_3));
    Odrv12 I__4910 (
            .O(N__33195),
            .I(data_out_frame_9_3));
    InMux I__4909 (
            .O(N__33190),
            .I(N__33187));
    LocalMux I__4908 (
            .O(N__33187),
            .I(N__33184));
    Span4Mux_h I__4907 (
            .O(N__33184),
            .I(N__33181));
    Odrv4 I__4906 (
            .O(N__33181),
            .I(\c0.n21641 ));
    CascadeMux I__4905 (
            .O(N__33178),
            .I(N__33174));
    CascadeMux I__4904 (
            .O(N__33177),
            .I(N__33171));
    InMux I__4903 (
            .O(N__33174),
            .I(N__33166));
    InMux I__4902 (
            .O(N__33171),
            .I(N__33166));
    LocalMux I__4901 (
            .O(N__33166),
            .I(data_out_frame_8_3));
    InMux I__4900 (
            .O(N__33163),
            .I(N__33160));
    LocalMux I__4899 (
            .O(N__33160),
            .I(N__33157));
    Span4Mux_h I__4898 (
            .O(N__33157),
            .I(N__33154));
    Span4Mux_v I__4897 (
            .O(N__33154),
            .I(N__33151));
    Odrv4 I__4896 (
            .O(N__33151),
            .I(\c0.n21644 ));
    CascadeMux I__4895 (
            .O(N__33148),
            .I(N__33145));
    InMux I__4894 (
            .O(N__33145),
            .I(N__33142));
    LocalMux I__4893 (
            .O(N__33142),
            .I(N__33138));
    InMux I__4892 (
            .O(N__33141),
            .I(N__33135));
    Span4Mux_v I__4891 (
            .O(N__33138),
            .I(N__33132));
    LocalMux I__4890 (
            .O(N__33135),
            .I(data_out_frame_11_5));
    Odrv4 I__4889 (
            .O(N__33132),
            .I(data_out_frame_11_5));
    InMux I__4888 (
            .O(N__33127),
            .I(N__33123));
    InMux I__4887 (
            .O(N__33126),
            .I(N__33120));
    LocalMux I__4886 (
            .O(N__33123),
            .I(N__33117));
    LocalMux I__4885 (
            .O(N__33120),
            .I(data_out_frame_8_5));
    Odrv12 I__4884 (
            .O(N__33117),
            .I(data_out_frame_8_5));
    CascadeMux I__4883 (
            .O(N__33112),
            .I(\c0.n21635_cascade_ ));
    InMux I__4882 (
            .O(N__33109),
            .I(N__33106));
    LocalMux I__4881 (
            .O(N__33106),
            .I(N__33103));
    Span4Mux_h I__4880 (
            .O(N__33103),
            .I(N__33099));
    InMux I__4879 (
            .O(N__33102),
            .I(N__33096));
    Span4Mux_h I__4878 (
            .O(N__33099),
            .I(N__33093));
    LocalMux I__4877 (
            .O(N__33096),
            .I(data_out_frame_9_5));
    Odrv4 I__4876 (
            .O(N__33093),
            .I(data_out_frame_9_5));
    CascadeMux I__4875 (
            .O(N__33088),
            .I(N__33084));
    InMux I__4874 (
            .O(N__33087),
            .I(N__33081));
    InMux I__4873 (
            .O(N__33084),
            .I(N__33078));
    LocalMux I__4872 (
            .O(N__33081),
            .I(data_out_frame_5_3));
    LocalMux I__4871 (
            .O(N__33078),
            .I(data_out_frame_5_3));
    CascadeMux I__4870 (
            .O(N__33073),
            .I(N__33070));
    InMux I__4869 (
            .O(N__33070),
            .I(N__33067));
    LocalMux I__4868 (
            .O(N__33067),
            .I(N__33064));
    Span4Mux_h I__4867 (
            .O(N__33064),
            .I(N__33060));
    InMux I__4866 (
            .O(N__33063),
            .I(N__33057));
    Span4Mux_v I__4865 (
            .O(N__33060),
            .I(N__33054));
    LocalMux I__4864 (
            .O(N__33057),
            .I(data_out_frame_28_4));
    Odrv4 I__4863 (
            .O(N__33054),
            .I(data_out_frame_28_4));
    InMux I__4862 (
            .O(N__33049),
            .I(N__33046));
    LocalMux I__4861 (
            .O(N__33046),
            .I(N__33043));
    Span4Mux_v I__4860 (
            .O(N__33043),
            .I(N__33040));
    Odrv4 I__4859 (
            .O(N__33040),
            .I(n2342));
    CascadeMux I__4858 (
            .O(N__33037),
            .I(N__33033));
    InMux I__4857 (
            .O(N__33036),
            .I(N__33030));
    InMux I__4856 (
            .O(N__33033),
            .I(N__33027));
    LocalMux I__4855 (
            .O(N__33030),
            .I(N__33024));
    LocalMux I__4854 (
            .O(N__33027),
            .I(N__33020));
    Span4Mux_v I__4853 (
            .O(N__33024),
            .I(N__33017));
    InMux I__4852 (
            .O(N__33023),
            .I(N__33014));
    Span4Mux_h I__4851 (
            .O(N__33020),
            .I(N__33011));
    Odrv4 I__4850 (
            .O(N__33017),
            .I(encoder1_position_3));
    LocalMux I__4849 (
            .O(N__33014),
            .I(encoder1_position_3));
    Odrv4 I__4848 (
            .O(N__33011),
            .I(encoder1_position_3));
    InMux I__4847 (
            .O(N__33004),
            .I(N__32999));
    CascadeMux I__4846 (
            .O(N__33003),
            .I(N__32996));
    InMux I__4845 (
            .O(N__33002),
            .I(N__32993));
    LocalMux I__4844 (
            .O(N__32999),
            .I(N__32990));
    InMux I__4843 (
            .O(N__32996),
            .I(N__32987));
    LocalMux I__4842 (
            .O(N__32993),
            .I(encoder0_position_19));
    Odrv12 I__4841 (
            .O(N__32990),
            .I(encoder0_position_19));
    LocalMux I__4840 (
            .O(N__32987),
            .I(encoder0_position_19));
    CascadeMux I__4839 (
            .O(N__32980),
            .I(\c0.n6_adj_3379_cascade_ ));
    InMux I__4838 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__4837 (
            .O(N__32974),
            .I(N__32971));
    Span4Mux_h I__4836 (
            .O(N__32971),
            .I(N__32968));
    Odrv4 I__4835 (
            .O(N__32968),
            .I(n2324));
    CascadeMux I__4834 (
            .O(N__32965),
            .I(N__32961));
    InMux I__4833 (
            .O(N__32964),
            .I(N__32958));
    InMux I__4832 (
            .O(N__32961),
            .I(N__32954));
    LocalMux I__4831 (
            .O(N__32958),
            .I(N__32951));
    InMux I__4830 (
            .O(N__32957),
            .I(N__32948));
    LocalMux I__4829 (
            .O(N__32954),
            .I(N__32945));
    Odrv4 I__4828 (
            .O(N__32951),
            .I(encoder1_position_21));
    LocalMux I__4827 (
            .O(N__32948),
            .I(encoder1_position_21));
    Odrv4 I__4826 (
            .O(N__32945),
            .I(encoder1_position_21));
    InMux I__4825 (
            .O(N__32938),
            .I(N__32935));
    LocalMux I__4824 (
            .O(N__32935),
            .I(N__32932));
    Span4Mux_h I__4823 (
            .O(N__32932),
            .I(N__32929));
    Span4Mux_h I__4822 (
            .O(N__32929),
            .I(N__32926));
    Odrv4 I__4821 (
            .O(N__32926),
            .I(\c0.n21559 ));
    InMux I__4820 (
            .O(N__32923),
            .I(N__32920));
    LocalMux I__4819 (
            .O(N__32920),
            .I(N__32917));
    Span4Mux_h I__4818 (
            .O(N__32917),
            .I(N__32914));
    Odrv4 I__4817 (
            .O(N__32914),
            .I(\c0.n5_adj_3102 ));
    InMux I__4816 (
            .O(N__32911),
            .I(N__32908));
    LocalMux I__4815 (
            .O(N__32908),
            .I(N__32905));
    Span4Mux_v I__4814 (
            .O(N__32905),
            .I(N__32902));
    Span4Mux_v I__4813 (
            .O(N__32902),
            .I(N__32899));
    Odrv4 I__4812 (
            .O(N__32899),
            .I(n2322));
    InMux I__4811 (
            .O(N__32896),
            .I(N__32893));
    LocalMux I__4810 (
            .O(N__32893),
            .I(N__32890));
    Span4Mux_h I__4809 (
            .O(N__32890),
            .I(N__32886));
    CascadeMux I__4808 (
            .O(N__32889),
            .I(N__32882));
    Span4Mux_h I__4807 (
            .O(N__32886),
            .I(N__32879));
    InMux I__4806 (
            .O(N__32885),
            .I(N__32876));
    InMux I__4805 (
            .O(N__32882),
            .I(N__32873));
    Odrv4 I__4804 (
            .O(N__32879),
            .I(encoder0_position_24));
    LocalMux I__4803 (
            .O(N__32876),
            .I(encoder0_position_24));
    LocalMux I__4802 (
            .O(N__32873),
            .I(encoder0_position_24));
    InMux I__4801 (
            .O(N__32866),
            .I(N__32863));
    LocalMux I__4800 (
            .O(N__32863),
            .I(N__32860));
    Odrv4 I__4799 (
            .O(N__32860),
            .I(n2340));
    InMux I__4798 (
            .O(N__32857),
            .I(N__32854));
    LocalMux I__4797 (
            .O(N__32854),
            .I(N__32850));
    CascadeMux I__4796 (
            .O(N__32853),
            .I(N__32847));
    Span4Mux_h I__4795 (
            .O(N__32850),
            .I(N__32844));
    InMux I__4794 (
            .O(N__32847),
            .I(N__32840));
    Sp12to4 I__4793 (
            .O(N__32844),
            .I(N__32837));
    InMux I__4792 (
            .O(N__32843),
            .I(N__32834));
    LocalMux I__4791 (
            .O(N__32840),
            .I(N__32831));
    Odrv12 I__4790 (
            .O(N__32837),
            .I(encoder1_position_5));
    LocalMux I__4789 (
            .O(N__32834),
            .I(encoder1_position_5));
    Odrv4 I__4788 (
            .O(N__32831),
            .I(encoder1_position_5));
    CascadeMux I__4787 (
            .O(N__32824),
            .I(N__32821));
    InMux I__4786 (
            .O(N__32821),
            .I(N__32818));
    LocalMux I__4785 (
            .O(N__32818),
            .I(N__32815));
    Span4Mux_h I__4784 (
            .O(N__32815),
            .I(N__32812));
    Span4Mux_h I__4783 (
            .O(N__32812),
            .I(N__32809));
    Odrv4 I__4782 (
            .O(N__32809),
            .I(\c0.n21647 ));
    InMux I__4781 (
            .O(N__32806),
            .I(N__32803));
    LocalMux I__4780 (
            .O(N__32803),
            .I(N__32800));
    Span4Mux_v I__4779 (
            .O(N__32800),
            .I(N__32795));
    InMux I__4778 (
            .O(N__32799),
            .I(N__32792));
    InMux I__4777 (
            .O(N__32798),
            .I(N__32789));
    Odrv4 I__4776 (
            .O(N__32795),
            .I(encoder1_position_26));
    LocalMux I__4775 (
            .O(N__32792),
            .I(encoder1_position_26));
    LocalMux I__4774 (
            .O(N__32789),
            .I(encoder1_position_26));
    InMux I__4773 (
            .O(N__32782),
            .I(N__32776));
    InMux I__4772 (
            .O(N__32781),
            .I(N__32776));
    LocalMux I__4771 (
            .O(N__32776),
            .I(data_out_frame_10_2));
    SRMux I__4770 (
            .O(N__32773),
            .I(N__32770));
    LocalMux I__4769 (
            .O(N__32770),
            .I(N__32767));
    Odrv4 I__4768 (
            .O(N__32767),
            .I(\c0.n6_adj_3154 ));
    InMux I__4767 (
            .O(N__32764),
            .I(N__32760));
    InMux I__4766 (
            .O(N__32763),
            .I(N__32757));
    LocalMux I__4765 (
            .O(N__32760),
            .I(N__32754));
    LocalMux I__4764 (
            .O(N__32757),
            .I(data_out_frame_6_0));
    Odrv4 I__4763 (
            .O(N__32754),
            .I(data_out_frame_6_0));
    InMux I__4762 (
            .O(N__32749),
            .I(N__32746));
    LocalMux I__4761 (
            .O(N__32746),
            .I(N__32743));
    Span4Mux_h I__4760 (
            .O(N__32743),
            .I(N__32740));
    Odrv4 I__4759 (
            .O(N__32740),
            .I(\c0.n6_adj_3321 ));
    InMux I__4758 (
            .O(N__32737),
            .I(N__32734));
    LocalMux I__4757 (
            .O(N__32734),
            .I(N__32731));
    Span4Mux_h I__4756 (
            .O(N__32731),
            .I(N__32728));
    Odrv4 I__4755 (
            .O(N__32728),
            .I(n2344));
    InMux I__4754 (
            .O(N__32725),
            .I(N__32688));
    InMux I__4753 (
            .O(N__32724),
            .I(N__32688));
    InMux I__4752 (
            .O(N__32723),
            .I(N__32688));
    InMux I__4751 (
            .O(N__32722),
            .I(N__32679));
    InMux I__4750 (
            .O(N__32721),
            .I(N__32679));
    InMux I__4749 (
            .O(N__32720),
            .I(N__32679));
    InMux I__4748 (
            .O(N__32719),
            .I(N__32679));
    InMux I__4747 (
            .O(N__32718),
            .I(N__32672));
    InMux I__4746 (
            .O(N__32717),
            .I(N__32672));
    InMux I__4745 (
            .O(N__32716),
            .I(N__32672));
    InMux I__4744 (
            .O(N__32715),
            .I(N__32663));
    InMux I__4743 (
            .O(N__32714),
            .I(N__32663));
    InMux I__4742 (
            .O(N__32713),
            .I(N__32663));
    InMux I__4741 (
            .O(N__32712),
            .I(N__32663));
    InMux I__4740 (
            .O(N__32711),
            .I(N__32656));
    InMux I__4739 (
            .O(N__32710),
            .I(N__32656));
    InMux I__4738 (
            .O(N__32709),
            .I(N__32656));
    InMux I__4737 (
            .O(N__32708),
            .I(N__32647));
    InMux I__4736 (
            .O(N__32707),
            .I(N__32647));
    InMux I__4735 (
            .O(N__32706),
            .I(N__32647));
    InMux I__4734 (
            .O(N__32705),
            .I(N__32647));
    CascadeMux I__4733 (
            .O(N__32704),
            .I(N__32615));
    CascadeMux I__4732 (
            .O(N__32703),
            .I(N__32610));
    CascadeMux I__4731 (
            .O(N__32702),
            .I(N__32606));
    CascadeMux I__4730 (
            .O(N__32701),
            .I(N__32602));
    CascadeMux I__4729 (
            .O(N__32700),
            .I(N__32597));
    CascadeMux I__4728 (
            .O(N__32699),
            .I(N__32593));
    CascadeMux I__4727 (
            .O(N__32698),
            .I(N__32589));
    CascadeMux I__4726 (
            .O(N__32697),
            .I(N__32575));
    CascadeMux I__4725 (
            .O(N__32696),
            .I(N__32571));
    CascadeMux I__4724 (
            .O(N__32695),
            .I(N__32567));
    LocalMux I__4723 (
            .O(N__32688),
            .I(N__32550));
    LocalMux I__4722 (
            .O(N__32679),
            .I(N__32550));
    LocalMux I__4721 (
            .O(N__32672),
            .I(N__32550));
    LocalMux I__4720 (
            .O(N__32663),
            .I(N__32550));
    LocalMux I__4719 (
            .O(N__32656),
            .I(N__32550));
    LocalMux I__4718 (
            .O(N__32647),
            .I(N__32550));
    InMux I__4717 (
            .O(N__32646),
            .I(N__32543));
    InMux I__4716 (
            .O(N__32645),
            .I(N__32543));
    InMux I__4715 (
            .O(N__32644),
            .I(N__32543));
    InMux I__4714 (
            .O(N__32643),
            .I(N__32534));
    InMux I__4713 (
            .O(N__32642),
            .I(N__32534));
    InMux I__4712 (
            .O(N__32641),
            .I(N__32534));
    InMux I__4711 (
            .O(N__32640),
            .I(N__32534));
    InMux I__4710 (
            .O(N__32639),
            .I(N__32527));
    InMux I__4709 (
            .O(N__32638),
            .I(N__32527));
    InMux I__4708 (
            .O(N__32637),
            .I(N__32527));
    InMux I__4707 (
            .O(N__32636),
            .I(N__32518));
    InMux I__4706 (
            .O(N__32635),
            .I(N__32518));
    InMux I__4705 (
            .O(N__32634),
            .I(N__32518));
    InMux I__4704 (
            .O(N__32633),
            .I(N__32518));
    InMux I__4703 (
            .O(N__32632),
            .I(N__32511));
    InMux I__4702 (
            .O(N__32631),
            .I(N__32511));
    InMux I__4701 (
            .O(N__32630),
            .I(N__32511));
    InMux I__4700 (
            .O(N__32629),
            .I(N__32502));
    InMux I__4699 (
            .O(N__32628),
            .I(N__32502));
    InMux I__4698 (
            .O(N__32627),
            .I(N__32502));
    InMux I__4697 (
            .O(N__32626),
            .I(N__32502));
    InMux I__4696 (
            .O(N__32625),
            .I(N__32495));
    InMux I__4695 (
            .O(N__32624),
            .I(N__32495));
    InMux I__4694 (
            .O(N__32623),
            .I(N__32495));
    InMux I__4693 (
            .O(N__32622),
            .I(N__32486));
    InMux I__4692 (
            .O(N__32621),
            .I(N__32486));
    InMux I__4691 (
            .O(N__32620),
            .I(N__32486));
    InMux I__4690 (
            .O(N__32619),
            .I(N__32486));
    InMux I__4689 (
            .O(N__32618),
            .I(N__32451));
    InMux I__4688 (
            .O(N__32615),
            .I(N__32451));
    InMux I__4687 (
            .O(N__32614),
            .I(N__32451));
    InMux I__4686 (
            .O(N__32613),
            .I(N__32436));
    InMux I__4685 (
            .O(N__32610),
            .I(N__32436));
    InMux I__4684 (
            .O(N__32609),
            .I(N__32436));
    InMux I__4683 (
            .O(N__32606),
            .I(N__32436));
    InMux I__4682 (
            .O(N__32605),
            .I(N__32436));
    InMux I__4681 (
            .O(N__32602),
            .I(N__32436));
    InMux I__4680 (
            .O(N__32601),
            .I(N__32436));
    InMux I__4679 (
            .O(N__32600),
            .I(N__32421));
    InMux I__4678 (
            .O(N__32597),
            .I(N__32421));
    InMux I__4677 (
            .O(N__32596),
            .I(N__32421));
    InMux I__4676 (
            .O(N__32593),
            .I(N__32421));
    InMux I__4675 (
            .O(N__32592),
            .I(N__32421));
    InMux I__4674 (
            .O(N__32589),
            .I(N__32421));
    InMux I__4673 (
            .O(N__32588),
            .I(N__32421));
    CascadeMux I__4672 (
            .O(N__32587),
            .I(N__32417));
    CascadeMux I__4671 (
            .O(N__32586),
            .I(N__32413));
    CascadeMux I__4670 (
            .O(N__32585),
            .I(N__32409));
    CascadeMux I__4669 (
            .O(N__32584),
            .I(N__32404));
    CascadeMux I__4668 (
            .O(N__32583),
            .I(N__32400));
    CascadeMux I__4667 (
            .O(N__32582),
            .I(N__32396));
    CascadeMux I__4666 (
            .O(N__32581),
            .I(N__32391));
    CascadeMux I__4665 (
            .O(N__32580),
            .I(N__32387));
    CascadeMux I__4664 (
            .O(N__32579),
            .I(N__32383));
    InMux I__4663 (
            .O(N__32578),
            .I(N__32361));
    InMux I__4662 (
            .O(N__32575),
            .I(N__32361));
    InMux I__4661 (
            .O(N__32574),
            .I(N__32361));
    InMux I__4660 (
            .O(N__32571),
            .I(N__32361));
    InMux I__4659 (
            .O(N__32570),
            .I(N__32361));
    InMux I__4658 (
            .O(N__32567),
            .I(N__32361));
    InMux I__4657 (
            .O(N__32566),
            .I(N__32361));
    CascadeMux I__4656 (
            .O(N__32565),
            .I(N__32357));
    CascadeMux I__4655 (
            .O(N__32564),
            .I(N__32353));
    CascadeMux I__4654 (
            .O(N__32563),
            .I(N__32349));
    Span4Mux_v I__4653 (
            .O(N__32550),
            .I(N__32329));
    LocalMux I__4652 (
            .O(N__32543),
            .I(N__32329));
    LocalMux I__4651 (
            .O(N__32534),
            .I(N__32329));
    LocalMux I__4650 (
            .O(N__32527),
            .I(N__32329));
    LocalMux I__4649 (
            .O(N__32518),
            .I(N__32329));
    LocalMux I__4648 (
            .O(N__32511),
            .I(N__32329));
    LocalMux I__4647 (
            .O(N__32502),
            .I(N__32329));
    LocalMux I__4646 (
            .O(N__32495),
            .I(N__32329));
    LocalMux I__4645 (
            .O(N__32486),
            .I(N__32329));
    InMux I__4644 (
            .O(N__32485),
            .I(N__32322));
    InMux I__4643 (
            .O(N__32484),
            .I(N__32322));
    InMux I__4642 (
            .O(N__32483),
            .I(N__32322));
    InMux I__4641 (
            .O(N__32482),
            .I(N__32313));
    InMux I__4640 (
            .O(N__32481),
            .I(N__32313));
    InMux I__4639 (
            .O(N__32480),
            .I(N__32313));
    InMux I__4638 (
            .O(N__32479),
            .I(N__32313));
    InMux I__4637 (
            .O(N__32478),
            .I(N__32306));
    InMux I__4636 (
            .O(N__32477),
            .I(N__32306));
    InMux I__4635 (
            .O(N__32476),
            .I(N__32306));
    InMux I__4634 (
            .O(N__32475),
            .I(N__32297));
    InMux I__4633 (
            .O(N__32474),
            .I(N__32297));
    InMux I__4632 (
            .O(N__32473),
            .I(N__32297));
    InMux I__4631 (
            .O(N__32472),
            .I(N__32297));
    InMux I__4630 (
            .O(N__32471),
            .I(N__32290));
    InMux I__4629 (
            .O(N__32470),
            .I(N__32290));
    InMux I__4628 (
            .O(N__32469),
            .I(N__32290));
    InMux I__4627 (
            .O(N__32468),
            .I(N__32281));
    InMux I__4626 (
            .O(N__32467),
            .I(N__32281));
    InMux I__4625 (
            .O(N__32466),
            .I(N__32281));
    InMux I__4624 (
            .O(N__32465),
            .I(N__32281));
    InMux I__4623 (
            .O(N__32464),
            .I(N__32274));
    InMux I__4622 (
            .O(N__32463),
            .I(N__32274));
    InMux I__4621 (
            .O(N__32462),
            .I(N__32274));
    InMux I__4620 (
            .O(N__32461),
            .I(N__32265));
    InMux I__4619 (
            .O(N__32460),
            .I(N__32265));
    InMux I__4618 (
            .O(N__32459),
            .I(N__32265));
    InMux I__4617 (
            .O(N__32458),
            .I(N__32265));
    LocalMux I__4616 (
            .O(N__32451),
            .I(N__32251));
    LocalMux I__4615 (
            .O(N__32436),
            .I(N__32251));
    LocalMux I__4614 (
            .O(N__32421),
            .I(N__32251));
    InMux I__4613 (
            .O(N__32420),
            .I(N__32236));
    InMux I__4612 (
            .O(N__32417),
            .I(N__32236));
    InMux I__4611 (
            .O(N__32416),
            .I(N__32236));
    InMux I__4610 (
            .O(N__32413),
            .I(N__32236));
    InMux I__4609 (
            .O(N__32412),
            .I(N__32236));
    InMux I__4608 (
            .O(N__32409),
            .I(N__32236));
    InMux I__4607 (
            .O(N__32408),
            .I(N__32236));
    InMux I__4606 (
            .O(N__32407),
            .I(N__32221));
    InMux I__4605 (
            .O(N__32404),
            .I(N__32221));
    InMux I__4604 (
            .O(N__32403),
            .I(N__32221));
    InMux I__4603 (
            .O(N__32400),
            .I(N__32221));
    InMux I__4602 (
            .O(N__32399),
            .I(N__32221));
    InMux I__4601 (
            .O(N__32396),
            .I(N__32221));
    InMux I__4600 (
            .O(N__32395),
            .I(N__32221));
    InMux I__4599 (
            .O(N__32394),
            .I(N__32206));
    InMux I__4598 (
            .O(N__32391),
            .I(N__32206));
    InMux I__4597 (
            .O(N__32390),
            .I(N__32206));
    InMux I__4596 (
            .O(N__32387),
            .I(N__32206));
    InMux I__4595 (
            .O(N__32386),
            .I(N__32206));
    InMux I__4594 (
            .O(N__32383),
            .I(N__32206));
    InMux I__4593 (
            .O(N__32382),
            .I(N__32206));
    CascadeMux I__4592 (
            .O(N__32381),
            .I(N__32202));
    CascadeMux I__4591 (
            .O(N__32380),
            .I(N__32198));
    CascadeMux I__4590 (
            .O(N__32379),
            .I(N__32194));
    CascadeMux I__4589 (
            .O(N__32378),
            .I(N__32189));
    CascadeMux I__4588 (
            .O(N__32377),
            .I(N__32185));
    CascadeMux I__4587 (
            .O(N__32376),
            .I(N__32181));
    LocalMux I__4586 (
            .O(N__32361),
            .I(N__32177));
    InMux I__4585 (
            .O(N__32360),
            .I(N__32162));
    InMux I__4584 (
            .O(N__32357),
            .I(N__32162));
    InMux I__4583 (
            .O(N__32356),
            .I(N__32162));
    InMux I__4582 (
            .O(N__32353),
            .I(N__32162));
    InMux I__4581 (
            .O(N__32352),
            .I(N__32162));
    InMux I__4580 (
            .O(N__32349),
            .I(N__32162));
    InMux I__4579 (
            .O(N__32348),
            .I(N__32162));
    Span4Mux_v I__4578 (
            .O(N__32329),
            .I(N__32129));
    LocalMux I__4577 (
            .O(N__32322),
            .I(N__32129));
    LocalMux I__4576 (
            .O(N__32313),
            .I(N__32129));
    LocalMux I__4575 (
            .O(N__32306),
            .I(N__32129));
    LocalMux I__4574 (
            .O(N__32297),
            .I(N__32129));
    LocalMux I__4573 (
            .O(N__32290),
            .I(N__32129));
    LocalMux I__4572 (
            .O(N__32281),
            .I(N__32129));
    LocalMux I__4571 (
            .O(N__32274),
            .I(N__32129));
    LocalMux I__4570 (
            .O(N__32265),
            .I(N__32129));
    InMux I__4569 (
            .O(N__32264),
            .I(N__32122));
    InMux I__4568 (
            .O(N__32263),
            .I(N__32122));
    InMux I__4567 (
            .O(N__32262),
            .I(N__32122));
    InMux I__4566 (
            .O(N__32261),
            .I(N__32113));
    InMux I__4565 (
            .O(N__32260),
            .I(N__32113));
    InMux I__4564 (
            .O(N__32259),
            .I(N__32113));
    InMux I__4563 (
            .O(N__32258),
            .I(N__32113));
    Span4Mux_v I__4562 (
            .O(N__32251),
            .I(N__32104));
    LocalMux I__4561 (
            .O(N__32236),
            .I(N__32104));
    LocalMux I__4560 (
            .O(N__32221),
            .I(N__32104));
    LocalMux I__4559 (
            .O(N__32206),
            .I(N__32104));
    InMux I__4558 (
            .O(N__32205),
            .I(N__32089));
    InMux I__4557 (
            .O(N__32202),
            .I(N__32089));
    InMux I__4556 (
            .O(N__32201),
            .I(N__32089));
    InMux I__4555 (
            .O(N__32198),
            .I(N__32089));
    InMux I__4554 (
            .O(N__32197),
            .I(N__32089));
    InMux I__4553 (
            .O(N__32194),
            .I(N__32089));
    InMux I__4552 (
            .O(N__32193),
            .I(N__32089));
    InMux I__4551 (
            .O(N__32192),
            .I(N__32074));
    InMux I__4550 (
            .O(N__32189),
            .I(N__32074));
    InMux I__4549 (
            .O(N__32188),
            .I(N__32074));
    InMux I__4548 (
            .O(N__32185),
            .I(N__32074));
    InMux I__4547 (
            .O(N__32184),
            .I(N__32074));
    InMux I__4546 (
            .O(N__32181),
            .I(N__32074));
    InMux I__4545 (
            .O(N__32180),
            .I(N__32074));
    Span4Mux_v I__4544 (
            .O(N__32177),
            .I(N__32066));
    LocalMux I__4543 (
            .O(N__32162),
            .I(N__32066));
    InMux I__4542 (
            .O(N__32161),
            .I(N__32059));
    InMux I__4541 (
            .O(N__32160),
            .I(N__32059));
    InMux I__4540 (
            .O(N__32159),
            .I(N__32059));
    InMux I__4539 (
            .O(N__32158),
            .I(N__32050));
    InMux I__4538 (
            .O(N__32157),
            .I(N__32050));
    InMux I__4537 (
            .O(N__32156),
            .I(N__32050));
    InMux I__4536 (
            .O(N__32155),
            .I(N__32050));
    InMux I__4535 (
            .O(N__32154),
            .I(N__32043));
    InMux I__4534 (
            .O(N__32153),
            .I(N__32043));
    InMux I__4533 (
            .O(N__32152),
            .I(N__32043));
    InMux I__4532 (
            .O(N__32151),
            .I(N__32034));
    InMux I__4531 (
            .O(N__32150),
            .I(N__32034));
    InMux I__4530 (
            .O(N__32149),
            .I(N__32034));
    InMux I__4529 (
            .O(N__32148),
            .I(N__32034));
    Span4Mux_v I__4528 (
            .O(N__32129),
            .I(N__32027));
    LocalMux I__4527 (
            .O(N__32122),
            .I(N__32027));
    LocalMux I__4526 (
            .O(N__32113),
            .I(N__32027));
    Span4Mux_v I__4525 (
            .O(N__32104),
            .I(N__32020));
    LocalMux I__4524 (
            .O(N__32089),
            .I(N__32020));
    LocalMux I__4523 (
            .O(N__32074),
            .I(N__32020));
    CascadeMux I__4522 (
            .O(N__32073),
            .I(N__32009));
    CascadeMux I__4521 (
            .O(N__32072),
            .I(N__32005));
    CascadeMux I__4520 (
            .O(N__32071),
            .I(N__32001));
    Span4Mux_v I__4519 (
            .O(N__32066),
            .I(N__31982));
    LocalMux I__4518 (
            .O(N__32059),
            .I(N__31982));
    LocalMux I__4517 (
            .O(N__32050),
            .I(N__31982));
    LocalMux I__4516 (
            .O(N__32043),
            .I(N__31982));
    LocalMux I__4515 (
            .O(N__32034),
            .I(N__31982));
    Span4Mux_v I__4514 (
            .O(N__32027),
            .I(N__31977));
    Span4Mux_v I__4513 (
            .O(N__32020),
            .I(N__31977));
    InMux I__4512 (
            .O(N__32019),
            .I(N__31970));
    InMux I__4511 (
            .O(N__32018),
            .I(N__31970));
    InMux I__4510 (
            .O(N__32017),
            .I(N__31970));
    InMux I__4509 (
            .O(N__32016),
            .I(N__31961));
    InMux I__4508 (
            .O(N__32015),
            .I(N__31961));
    InMux I__4507 (
            .O(N__32014),
            .I(N__31961));
    InMux I__4506 (
            .O(N__32013),
            .I(N__31961));
    InMux I__4505 (
            .O(N__32012),
            .I(N__31946));
    InMux I__4504 (
            .O(N__32009),
            .I(N__31946));
    InMux I__4503 (
            .O(N__32008),
            .I(N__31946));
    InMux I__4502 (
            .O(N__32005),
            .I(N__31946));
    InMux I__4501 (
            .O(N__32004),
            .I(N__31946));
    InMux I__4500 (
            .O(N__32001),
            .I(N__31946));
    InMux I__4499 (
            .O(N__32000),
            .I(N__31946));
    InMux I__4498 (
            .O(N__31999),
            .I(N__31939));
    InMux I__4497 (
            .O(N__31998),
            .I(N__31939));
    InMux I__4496 (
            .O(N__31997),
            .I(N__31939));
    InMux I__4495 (
            .O(N__31996),
            .I(N__31930));
    InMux I__4494 (
            .O(N__31995),
            .I(N__31930));
    InMux I__4493 (
            .O(N__31994),
            .I(N__31930));
    InMux I__4492 (
            .O(N__31993),
            .I(N__31930));
    Odrv4 I__4491 (
            .O(N__31982),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4490 (
            .O(N__31977),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4489 (
            .O(N__31970),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4488 (
            .O(N__31961),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4487 (
            .O(N__31946),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4486 (
            .O(N__31939),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4485 (
            .O(N__31930),
            .I(CONSTANT_ONE_NET));
    InMux I__4484 (
            .O(N__31915),
            .I(bfn_14_32_0_));
    InMux I__4483 (
            .O(N__31912),
            .I(N__31909));
    LocalMux I__4482 (
            .O(N__31909),
            .I(N__31906));
    Span12Mux_h I__4481 (
            .O(N__31906),
            .I(N__31903));
    Span12Mux_v I__4480 (
            .O(N__31903),
            .I(N__31900));
    Odrv12 I__4479 (
            .O(N__31900),
            .I(n20764));
    InMux I__4478 (
            .O(N__31897),
            .I(N__31894));
    LocalMux I__4477 (
            .O(N__31894),
            .I(N__31891));
    Span4Mux_v I__4476 (
            .O(N__31891),
            .I(N__31888));
    Odrv4 I__4475 (
            .O(N__31888),
            .I(n16));
    SRMux I__4474 (
            .O(N__31885),
            .I(N__31882));
    LocalMux I__4473 (
            .O(N__31882),
            .I(N__31879));
    Span4Mux_h I__4472 (
            .O(N__31879),
            .I(N__31876));
    Odrv4 I__4471 (
            .O(N__31876),
            .I(\c0.n6_adj_3155 ));
    InMux I__4470 (
            .O(N__31873),
            .I(bfn_14_31_0_));
    InMux I__4469 (
            .O(N__31870),
            .I(bfn_14_29_0_));
    InMux I__4468 (
            .O(N__31867),
            .I(bfn_14_30_0_));
    InMux I__4467 (
            .O(N__31864),
            .I(bfn_14_28_0_));
    InMux I__4466 (
            .O(N__31861),
            .I(bfn_14_27_0_));
    InMux I__4465 (
            .O(N__31858),
            .I(bfn_14_26_0_));
    InMux I__4464 (
            .O(N__31855),
            .I(bfn_14_25_0_));
    InMux I__4463 (
            .O(N__31852),
            .I(bfn_14_24_0_));
    InMux I__4462 (
            .O(N__31849),
            .I(bfn_14_23_0_));
    SRMux I__4461 (
            .O(N__31846),
            .I(N__31843));
    LocalMux I__4460 (
            .O(N__31843),
            .I(N__31840));
    Span4Mux_h I__4459 (
            .O(N__31840),
            .I(N__31837));
    Odrv4 I__4458 (
            .O(N__31837),
            .I(\c0.n6_adj_3178 ));
    SRMux I__4457 (
            .O(N__31834),
            .I(N__31831));
    LocalMux I__4456 (
            .O(N__31831),
            .I(\c0.n6_adj_3182 ));
    InMux I__4455 (
            .O(N__31828),
            .I(bfn_14_22_0_));
    SRMux I__4454 (
            .O(N__31825),
            .I(N__31822));
    LocalMux I__4453 (
            .O(N__31822),
            .I(N__31819));
    Odrv4 I__4452 (
            .O(N__31819),
            .I(\c0.n6_adj_3180 ));
    InMux I__4451 (
            .O(N__31816),
            .I(bfn_14_20_0_));
    SRMux I__4450 (
            .O(N__31813),
            .I(N__31810));
    LocalMux I__4449 (
            .O(N__31810),
            .I(N__31807));
    Sp12to4 I__4448 (
            .O(N__31807),
            .I(N__31804));
    Odrv12 I__4447 (
            .O(N__31804),
            .I(\c0.n6_adj_3184 ));
    InMux I__4446 (
            .O(N__31801),
            .I(bfn_14_21_0_));
    InMux I__4445 (
            .O(N__31798),
            .I(bfn_14_19_0_));
    SRMux I__4444 (
            .O(N__31795),
            .I(N__31792));
    LocalMux I__4443 (
            .O(N__31792),
            .I(N__31789));
    Odrv4 I__4442 (
            .O(N__31789),
            .I(\c0.n6_adj_3186 ));
    InMux I__4441 (
            .O(N__31786),
            .I(bfn_14_18_0_));
    SRMux I__4440 (
            .O(N__31783),
            .I(N__31780));
    LocalMux I__4439 (
            .O(N__31780),
            .I(N__31777));
    Span4Mux_v I__4438 (
            .O(N__31777),
            .I(N__31774));
    Odrv4 I__4437 (
            .O(N__31774),
            .I(\c0.n6_adj_3188 ));
    InMux I__4436 (
            .O(N__31771),
            .I(bfn_14_17_0_));
    InMux I__4435 (
            .O(N__31768),
            .I(bfn_14_16_0_));
    InMux I__4434 (
            .O(N__31765),
            .I(bfn_14_15_0_));
    InMux I__4433 (
            .O(N__31762),
            .I(bfn_14_14_0_));
    SRMux I__4432 (
            .O(N__31759),
            .I(N__31756));
    LocalMux I__4431 (
            .O(N__31756),
            .I(N__31753));
    Span4Mux_v I__4430 (
            .O(N__31753),
            .I(N__31750));
    Odrv4 I__4429 (
            .O(N__31750),
            .I(\c0.n6_adj_3162 ));
    InMux I__4428 (
            .O(N__31747),
            .I(bfn_14_13_0_));
    InMux I__4427 (
            .O(N__31744),
            .I(bfn_14_11_0_));
    InMux I__4426 (
            .O(N__31741),
            .I(bfn_14_12_0_));
    InMux I__4425 (
            .O(N__31738),
            .I(bfn_14_10_0_));
    InMux I__4424 (
            .O(N__31735),
            .I(bfn_14_9_0_));
    InMux I__4423 (
            .O(N__31732),
            .I(bfn_14_8_0_));
    InMux I__4422 (
            .O(N__31729),
            .I(bfn_14_7_0_));
    InMux I__4421 (
            .O(N__31726),
            .I(\c0.n17177 ));
    InMux I__4420 (
            .O(N__31723),
            .I(N__31720));
    LocalMux I__4419 (
            .O(N__31720),
            .I(\c0.n2_adj_3145 ));
    InMux I__4418 (
            .O(N__31717),
            .I(\c0.n17178 ));
    InMux I__4417 (
            .O(N__31714),
            .I(\c0.n17179 ));
    InMux I__4416 (
            .O(N__31711),
            .I(bfn_14_6_0_));
    InMux I__4415 (
            .O(N__31708),
            .I(N__31705));
    LocalMux I__4414 (
            .O(N__31705),
            .I(N__31702));
    Odrv4 I__4413 (
            .O(N__31702),
            .I(\c0.n19638 ));
    CascadeMux I__4412 (
            .O(N__31699),
            .I(\c0.n6_adj_3515_cascade_ ));
    InMux I__4411 (
            .O(N__31696),
            .I(N__31693));
    LocalMux I__4410 (
            .O(N__31693),
            .I(\c0.n5_adj_3516 ));
    CascadeMux I__4409 (
            .O(N__31690),
            .I(N__31685));
    InMux I__4408 (
            .O(N__31689),
            .I(N__31682));
    InMux I__4407 (
            .O(N__31688),
            .I(N__31677));
    InMux I__4406 (
            .O(N__31685),
            .I(N__31677));
    LocalMux I__4405 (
            .O(N__31682),
            .I(\c0.FRAME_MATCHER_state_5 ));
    LocalMux I__4404 (
            .O(N__31677),
            .I(\c0.FRAME_MATCHER_state_5 ));
    SRMux I__4403 (
            .O(N__31672),
            .I(N__31669));
    LocalMux I__4402 (
            .O(N__31669),
            .I(\c0.n18681 ));
    CascadeMux I__4401 (
            .O(N__31666),
            .I(N__31663));
    InMux I__4400 (
            .O(N__31663),
            .I(N__31659));
    InMux I__4399 (
            .O(N__31662),
            .I(N__31655));
    LocalMux I__4398 (
            .O(N__31659),
            .I(N__31652));
    InMux I__4397 (
            .O(N__31658),
            .I(N__31649));
    LocalMux I__4396 (
            .O(N__31655),
            .I(N__31646));
    Span4Mux_h I__4395 (
            .O(N__31652),
            .I(N__31643));
    LocalMux I__4394 (
            .O(N__31649),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__4393 (
            .O(N__31646),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__4392 (
            .O(N__31643),
            .I(\c0.FRAME_MATCHER_state_17 ));
    SRMux I__4391 (
            .O(N__31636),
            .I(N__31633));
    LocalMux I__4390 (
            .O(N__31633),
            .I(N__31630));
    Odrv4 I__4389 (
            .O(N__31630),
            .I(\c0.n18657 ));
    InMux I__4388 (
            .O(N__31627),
            .I(N__31622));
    InMux I__4387 (
            .O(N__31626),
            .I(N__31619));
    InMux I__4386 (
            .O(N__31625),
            .I(N__31616));
    LocalMux I__4385 (
            .O(N__31622),
            .I(N__31613));
    LocalMux I__4384 (
            .O(N__31619),
            .I(\c0.FRAME_MATCHER_state_4 ));
    LocalMux I__4383 (
            .O(N__31616),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__4382 (
            .O(N__31613),
            .I(\c0.FRAME_MATCHER_state_4 ));
    SRMux I__4381 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__4380 (
            .O(N__31603),
            .I(N__31600));
    Odrv4 I__4379 (
            .O(N__31600),
            .I(\c0.n18629 ));
    InMux I__4378 (
            .O(N__31597),
            .I(\c0.n17176 ));
    InMux I__4377 (
            .O(N__31594),
            .I(N__31591));
    LocalMux I__4376 (
            .O(N__31591),
            .I(\c0.n2_adj_3144 ));
    CascadeMux I__4375 (
            .O(N__31588),
            .I(\c0.n19638_cascade_ ));
    InMux I__4374 (
            .O(N__31585),
            .I(N__31582));
    LocalMux I__4373 (
            .O(N__31582),
            .I(\c0.FRAME_MATCHER_state_31_N_1864_2 ));
    CascadeMux I__4372 (
            .O(N__31579),
            .I(\c0.n6_adj_3521_cascade_ ));
    CascadeMux I__4371 (
            .O(N__31576),
            .I(N__31572));
    InMux I__4370 (
            .O(N__31575),
            .I(N__31568));
    InMux I__4369 (
            .O(N__31572),
            .I(N__31565));
    InMux I__4368 (
            .O(N__31571),
            .I(N__31562));
    LocalMux I__4367 (
            .O(N__31568),
            .I(N__31559));
    LocalMux I__4366 (
            .O(N__31565),
            .I(N__31556));
    LocalMux I__4365 (
            .O(N__31562),
            .I(N__31553));
    Span4Mux_h I__4364 (
            .O(N__31559),
            .I(N__31550));
    Odrv12 I__4363 (
            .O(N__31556),
            .I(\c0.n936 ));
    Odrv4 I__4362 (
            .O(N__31553),
            .I(\c0.n936 ));
    Odrv4 I__4361 (
            .O(N__31550),
            .I(\c0.n936 ));
    InMux I__4360 (
            .O(N__31543),
            .I(N__31540));
    LocalMux I__4359 (
            .O(N__31540),
            .I(\c0.n11_adj_3370 ));
    InMux I__4358 (
            .O(N__31537),
            .I(N__31533));
    InMux I__4357 (
            .O(N__31536),
            .I(N__31530));
    LocalMux I__4356 (
            .O(N__31533),
            .I(N__31527));
    LocalMux I__4355 (
            .O(N__31530),
            .I(N__31524));
    Odrv12 I__4354 (
            .O(N__31527),
            .I(\c0.tx_transmit_N_2443 ));
    Odrv4 I__4353 (
            .O(N__31524),
            .I(\c0.tx_transmit_N_2443 ));
    InMux I__4352 (
            .O(N__31519),
            .I(N__31516));
    LocalMux I__4351 (
            .O(N__31516),
            .I(N__31513));
    Span4Mux_h I__4350 (
            .O(N__31513),
            .I(N__31510));
    Odrv4 I__4349 (
            .O(N__31510),
            .I(\c0.n21420 ));
    InMux I__4348 (
            .O(N__31507),
            .I(N__31503));
    InMux I__4347 (
            .O(N__31506),
            .I(N__31499));
    LocalMux I__4346 (
            .O(N__31503),
            .I(N__31496));
    InMux I__4345 (
            .O(N__31502),
            .I(N__31493));
    LocalMux I__4344 (
            .O(N__31499),
            .I(N__31488));
    Span4Mux_v I__4343 (
            .O(N__31496),
            .I(N__31488));
    LocalMux I__4342 (
            .O(N__31493),
            .I(N__31485));
    Odrv4 I__4341 (
            .O(N__31488),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv4 I__4340 (
            .O(N__31485),
            .I(\c0.FRAME_MATCHER_state_21 ));
    SRMux I__4339 (
            .O(N__31480),
            .I(N__31477));
    LocalMux I__4338 (
            .O(N__31477),
            .I(N__31474));
    Span4Mux_h I__4337 (
            .O(N__31474),
            .I(N__31471));
    Odrv4 I__4336 (
            .O(N__31471),
            .I(\c0.n18627 ));
    InMux I__4335 (
            .O(N__31468),
            .I(N__31465));
    LocalMux I__4334 (
            .O(N__31465),
            .I(N__31462));
    Odrv4 I__4333 (
            .O(N__31462),
            .I(\c0.n19650 ));
    InMux I__4332 (
            .O(N__31459),
            .I(\c0.n17349 ));
    InMux I__4331 (
            .O(N__31456),
            .I(\c0.n17350 ));
    InMux I__4330 (
            .O(N__31453),
            .I(\c0.n17351 ));
    InMux I__4329 (
            .O(N__31450),
            .I(\c0.n17352 ));
    SRMux I__4328 (
            .O(N__31447),
            .I(N__31444));
    LocalMux I__4327 (
            .O(N__31444),
            .I(N__31441));
    Span4Mux_v I__4326 (
            .O(N__31441),
            .I(N__31437));
    InMux I__4325 (
            .O(N__31440),
            .I(N__31434));
    Odrv4 I__4324 (
            .O(N__31437),
            .I(\c0.n19052 ));
    LocalMux I__4323 (
            .O(N__31434),
            .I(\c0.n19052 ));
    CascadeMux I__4322 (
            .O(N__31429),
            .I(N__31425));
    CascadeMux I__4321 (
            .O(N__31428),
            .I(N__31422));
    InMux I__4320 (
            .O(N__31425),
            .I(N__31419));
    InMux I__4319 (
            .O(N__31422),
            .I(N__31416));
    LocalMux I__4318 (
            .O(N__31419),
            .I(N__31413));
    LocalMux I__4317 (
            .O(N__31416),
            .I(\c0.n6_adj_3338 ));
    Odrv4 I__4316 (
            .O(N__31413),
            .I(\c0.n6_adj_3338 ));
    CEMux I__4315 (
            .O(N__31408),
            .I(N__31405));
    LocalMux I__4314 (
            .O(N__31405),
            .I(N__31402));
    Span4Mux_v I__4313 (
            .O(N__31402),
            .I(N__31399));
    Odrv4 I__4312 (
            .O(N__31399),
            .I(\c0.n12326 ));
    CascadeMux I__4311 (
            .O(N__31396),
            .I(\c0.n12326_cascade_ ));
    SRMux I__4310 (
            .O(N__31393),
            .I(N__31390));
    LocalMux I__4309 (
            .O(N__31390),
            .I(N__31387));
    Span4Mux_h I__4308 (
            .O(N__31387),
            .I(N__31384));
    Odrv4 I__4307 (
            .O(N__31384),
            .I(\c0.n12758 ));
    CascadeMux I__4306 (
            .O(N__31381),
            .I(\c0.n4_adj_3263_cascade_ ));
    CascadeMux I__4305 (
            .O(N__31378),
            .I(\c0.n936_cascade_ ));
    InMux I__4304 (
            .O(N__31375),
            .I(N__31372));
    LocalMux I__4303 (
            .O(N__31372),
            .I(\c0.n21566 ));
    CascadeMux I__4302 (
            .O(N__31369),
            .I(n10_cascade_));
    InMux I__4301 (
            .O(N__31366),
            .I(N__31363));
    LocalMux I__4300 (
            .O(N__31363),
            .I(N__31359));
    InMux I__4299 (
            .O(N__31362),
            .I(N__31356));
    Odrv4 I__4298 (
            .O(N__31359),
            .I(r_Tx_Data_3));
    LocalMux I__4297 (
            .O(N__31356),
            .I(r_Tx_Data_3));
    InMux I__4296 (
            .O(N__31351),
            .I(N__31345));
    InMux I__4295 (
            .O(N__31350),
            .I(N__31345));
    LocalMux I__4294 (
            .O(N__31345),
            .I(data_out_frame_12_1));
    InMux I__4293 (
            .O(N__31342),
            .I(N__31339));
    LocalMux I__4292 (
            .O(N__31339),
            .I(\c0.n11_adj_3104 ));
    InMux I__4291 (
            .O(N__31336),
            .I(N__31333));
    LocalMux I__4290 (
            .O(N__31333),
            .I(N__31330));
    Span4Mux_v I__4289 (
            .O(N__31330),
            .I(N__31327));
    Odrv4 I__4288 (
            .O(N__31327),
            .I(n10_adj_3593));
    InMux I__4287 (
            .O(N__31324),
            .I(N__31320));
    InMux I__4286 (
            .O(N__31323),
            .I(N__31317));
    LocalMux I__4285 (
            .O(N__31320),
            .I(r_Tx_Data_2));
    LocalMux I__4284 (
            .O(N__31317),
            .I(r_Tx_Data_2));
    InMux I__4283 (
            .O(N__31312),
            .I(\c0.n17346 ));
    InMux I__4282 (
            .O(N__31309),
            .I(\c0.n17347 ));
    InMux I__4281 (
            .O(N__31306),
            .I(\c0.n17348 ));
    CascadeMux I__4280 (
            .O(N__31303),
            .I(N__31299));
    CascadeMux I__4279 (
            .O(N__31302),
            .I(N__31296));
    InMux I__4278 (
            .O(N__31299),
            .I(N__31290));
    InMux I__4277 (
            .O(N__31296),
            .I(N__31290));
    CascadeMux I__4276 (
            .O(N__31295),
            .I(N__31287));
    LocalMux I__4275 (
            .O(N__31290),
            .I(N__31284));
    InMux I__4274 (
            .O(N__31287),
            .I(N__31281));
    Span4Mux_h I__4273 (
            .O(N__31284),
            .I(N__31278));
    LocalMux I__4272 (
            .O(N__31281),
            .I(tx_active));
    Odrv4 I__4271 (
            .O(N__31278),
            .I(tx_active));
    InMux I__4270 (
            .O(N__31273),
            .I(N__31267));
    InMux I__4269 (
            .O(N__31272),
            .I(N__31267));
    LocalMux I__4268 (
            .O(N__31267),
            .I(\c0.n15842 ));
    InMux I__4267 (
            .O(N__31264),
            .I(N__31261));
    LocalMux I__4266 (
            .O(N__31261),
            .I(N__31258));
    Span4Mux_h I__4265 (
            .O(N__31258),
            .I(N__31255));
    Odrv4 I__4264 (
            .O(N__31255),
            .I(\c0.n11_adj_3404 ));
    InMux I__4263 (
            .O(N__31252),
            .I(N__31249));
    LocalMux I__4262 (
            .O(N__31249),
            .I(\c0.n7_adj_3333 ));
    InMux I__4261 (
            .O(N__31246),
            .I(N__31243));
    LocalMux I__4260 (
            .O(N__31243),
            .I(N__31239));
    InMux I__4259 (
            .O(N__31242),
            .I(N__31236));
    Span4Mux_v I__4258 (
            .O(N__31239),
            .I(N__31233));
    LocalMux I__4257 (
            .O(N__31236),
            .I(data_out_frame_9_1));
    Odrv4 I__4256 (
            .O(N__31233),
            .I(data_out_frame_9_1));
    InMux I__4255 (
            .O(N__31228),
            .I(N__31225));
    LocalMux I__4254 (
            .O(N__31225),
            .I(\c0.n21605 ));
    CascadeMux I__4253 (
            .O(N__31222),
            .I(N__31219));
    InMux I__4252 (
            .O(N__31219),
            .I(N__31215));
    InMux I__4251 (
            .O(N__31218),
            .I(N__31212));
    LocalMux I__4250 (
            .O(N__31215),
            .I(N__31209));
    LocalMux I__4249 (
            .O(N__31212),
            .I(data_out_frame_8_1));
    Odrv4 I__4248 (
            .O(N__31209),
            .I(data_out_frame_8_1));
    CascadeMux I__4247 (
            .O(N__31204),
            .I(\c0.n21608_cascade_ ));
    InMux I__4246 (
            .O(N__31201),
            .I(N__31194));
    InMux I__4245 (
            .O(N__31200),
            .I(N__31194));
    InMux I__4244 (
            .O(N__31199),
            .I(N__31191));
    LocalMux I__4243 (
            .O(N__31194),
            .I(\c0.r_Tx_Data_0 ));
    LocalMux I__4242 (
            .O(N__31191),
            .I(\c0.r_Tx_Data_0 ));
    InMux I__4241 (
            .O(N__31186),
            .I(N__31183));
    LocalMux I__4240 (
            .O(N__31183),
            .I(N__31180));
    Span4Mux_h I__4239 (
            .O(N__31180),
            .I(N__31177));
    Odrv4 I__4238 (
            .O(N__31177),
            .I(\c0.n21466 ));
    InMux I__4237 (
            .O(N__31174),
            .I(N__31171));
    LocalMux I__4236 (
            .O(N__31171),
            .I(N__31168));
    Span4Mux_v I__4235 (
            .O(N__31168),
            .I(N__31164));
    CascadeMux I__4234 (
            .O(N__31167),
            .I(N__31160));
    Span4Mux_v I__4233 (
            .O(N__31164),
            .I(N__31157));
    InMux I__4232 (
            .O(N__31163),
            .I(N__31154));
    InMux I__4231 (
            .O(N__31160),
            .I(N__31151));
    Odrv4 I__4230 (
            .O(N__31157),
            .I(encoder1_position_9));
    LocalMux I__4229 (
            .O(N__31154),
            .I(encoder1_position_9));
    LocalMux I__4228 (
            .O(N__31151),
            .I(encoder1_position_9));
    InMux I__4227 (
            .O(N__31144),
            .I(N__31141));
    LocalMux I__4226 (
            .O(N__31141),
            .I(N__31137));
    CascadeMux I__4225 (
            .O(N__31140),
            .I(N__31134));
    Span4Mux_v I__4224 (
            .O(N__31137),
            .I(N__31131));
    InMux I__4223 (
            .O(N__31134),
            .I(N__31128));
    Span4Mux_v I__4222 (
            .O(N__31131),
            .I(N__31122));
    LocalMux I__4221 (
            .O(N__31128),
            .I(N__31122));
    InMux I__4220 (
            .O(N__31127),
            .I(N__31119));
    Span4Mux_h I__4219 (
            .O(N__31122),
            .I(N__31116));
    LocalMux I__4218 (
            .O(N__31119),
            .I(encoder0_position_0));
    Odrv4 I__4217 (
            .O(N__31116),
            .I(encoder0_position_0));
    CascadeMux I__4216 (
            .O(N__31111),
            .I(N__31106));
    InMux I__4215 (
            .O(N__31110),
            .I(N__31103));
    InMux I__4214 (
            .O(N__31109),
            .I(N__31100));
    InMux I__4213 (
            .O(N__31106),
            .I(N__31097));
    LocalMux I__4212 (
            .O(N__31103),
            .I(encoder1_position_25));
    LocalMux I__4211 (
            .O(N__31100),
            .I(encoder1_position_25));
    LocalMux I__4210 (
            .O(N__31097),
            .I(encoder1_position_25));
    CascadeMux I__4209 (
            .O(N__31090),
            .I(N__31087));
    InMux I__4208 (
            .O(N__31087),
            .I(N__31083));
    InMux I__4207 (
            .O(N__31086),
            .I(N__31080));
    LocalMux I__4206 (
            .O(N__31083),
            .I(N__31076));
    LocalMux I__4205 (
            .O(N__31080),
            .I(N__31073));
    InMux I__4204 (
            .O(N__31079),
            .I(N__31070));
    Span4Mux_h I__4203 (
            .O(N__31076),
            .I(N__31067));
    Odrv4 I__4202 (
            .O(N__31073),
            .I(encoder1_position_2));
    LocalMux I__4201 (
            .O(N__31070),
            .I(encoder1_position_2));
    Odrv4 I__4200 (
            .O(N__31067),
            .I(encoder1_position_2));
    InMux I__4199 (
            .O(N__31060),
            .I(N__31057));
    LocalMux I__4198 (
            .O(N__31057),
            .I(N__31053));
    CascadeMux I__4197 (
            .O(N__31056),
            .I(N__31049));
    Span4Mux_v I__4196 (
            .O(N__31053),
            .I(N__31046));
    InMux I__4195 (
            .O(N__31052),
            .I(N__31043));
    InMux I__4194 (
            .O(N__31049),
            .I(N__31040));
    Odrv4 I__4193 (
            .O(N__31046),
            .I(encoder1_position_17));
    LocalMux I__4192 (
            .O(N__31043),
            .I(encoder1_position_17));
    LocalMux I__4191 (
            .O(N__31040),
            .I(encoder1_position_17));
    CascadeMux I__4190 (
            .O(N__31033),
            .I(N__31029));
    CascadeMux I__4189 (
            .O(N__31032),
            .I(N__31026));
    InMux I__4188 (
            .O(N__31029),
            .I(N__31021));
    InMux I__4187 (
            .O(N__31026),
            .I(N__31021));
    LocalMux I__4186 (
            .O(N__31021),
            .I(data_out_frame_13_2));
    InMux I__4185 (
            .O(N__31018),
            .I(N__31014));
    InMux I__4184 (
            .O(N__31017),
            .I(N__31011));
    LocalMux I__4183 (
            .O(N__31014),
            .I(data_out_frame_12_2));
    LocalMux I__4182 (
            .O(N__31011),
            .I(data_out_frame_12_2));
    InMux I__4181 (
            .O(N__31006),
            .I(N__31003));
    LocalMux I__4180 (
            .O(N__31003),
            .I(N__31000));
    Sp12to4 I__4179 (
            .O(N__31000),
            .I(N__30997));
    Odrv12 I__4178 (
            .O(N__30997),
            .I(\c0.n11_adj_3108 ));
    InMux I__4177 (
            .O(N__30994),
            .I(N__30990));
    InMux I__4176 (
            .O(N__30993),
            .I(N__30987));
    LocalMux I__4175 (
            .O(N__30990),
            .I(data_out_frame_10_1));
    LocalMux I__4174 (
            .O(N__30987),
            .I(data_out_frame_10_1));
    CascadeMux I__4173 (
            .O(N__30982),
            .I(N__30978));
    InMux I__4172 (
            .O(N__30981),
            .I(N__30973));
    InMux I__4171 (
            .O(N__30978),
            .I(N__30973));
    LocalMux I__4170 (
            .O(N__30973),
            .I(data_out_frame_11_1));
    InMux I__4169 (
            .O(N__30970),
            .I(N__30966));
    InMux I__4168 (
            .O(N__30969),
            .I(N__30963));
    LocalMux I__4167 (
            .O(N__30966),
            .I(N__30960));
    LocalMux I__4166 (
            .O(N__30963),
            .I(data_out_frame_13_5));
    Odrv4 I__4165 (
            .O(N__30960),
            .I(data_out_frame_13_5));
    InMux I__4164 (
            .O(N__30955),
            .I(N__30949));
    InMux I__4163 (
            .O(N__30954),
            .I(N__30944));
    InMux I__4162 (
            .O(N__30953),
            .I(N__30944));
    CascadeMux I__4161 (
            .O(N__30952),
            .I(N__30940));
    LocalMux I__4160 (
            .O(N__30949),
            .I(N__30935));
    LocalMux I__4159 (
            .O(N__30944),
            .I(N__30935));
    InMux I__4158 (
            .O(N__30943),
            .I(N__30932));
    InMux I__4157 (
            .O(N__30940),
            .I(N__30929));
    Span4Mux_h I__4156 (
            .O(N__30935),
            .I(N__30926));
    LocalMux I__4155 (
            .O(N__30932),
            .I(\c0.r_SM_Main_2_N_2547_0 ));
    LocalMux I__4154 (
            .O(N__30929),
            .I(\c0.r_SM_Main_2_N_2547_0 ));
    Odrv4 I__4153 (
            .O(N__30926),
            .I(\c0.r_SM_Main_2_N_2547_0 ));
    CascadeMux I__4152 (
            .O(N__30919),
            .I(N__30915));
    InMux I__4151 (
            .O(N__30918),
            .I(N__30912));
    InMux I__4150 (
            .O(N__30915),
            .I(N__30909));
    LocalMux I__4149 (
            .O(N__30912),
            .I(N__30905));
    LocalMux I__4148 (
            .O(N__30909),
            .I(N__30902));
    InMux I__4147 (
            .O(N__30908),
            .I(N__30899));
    Span4Mux_h I__4146 (
            .O(N__30905),
            .I(N__30894));
    Span4Mux_h I__4145 (
            .O(N__30902),
            .I(N__30894));
    LocalMux I__4144 (
            .O(N__30899),
            .I(encoder1_position_4));
    Odrv4 I__4143 (
            .O(N__30894),
            .I(encoder1_position_4));
    InMux I__4142 (
            .O(N__30889),
            .I(N__30886));
    LocalMux I__4141 (
            .O(N__30886),
            .I(N__30882));
    InMux I__4140 (
            .O(N__30885),
            .I(N__30879));
    Span4Mux_h I__4139 (
            .O(N__30882),
            .I(N__30876));
    LocalMux I__4138 (
            .O(N__30879),
            .I(data_out_frame_13_4));
    Odrv4 I__4137 (
            .O(N__30876),
            .I(data_out_frame_13_4));
    InMux I__4136 (
            .O(N__30871),
            .I(N__30862));
    InMux I__4135 (
            .O(N__30870),
            .I(N__30862));
    InMux I__4134 (
            .O(N__30869),
            .I(N__30862));
    LocalMux I__4133 (
            .O(N__30862),
            .I(encoder1_position_31));
    InMux I__4132 (
            .O(N__30859),
            .I(N__30856));
    LocalMux I__4131 (
            .O(N__30856),
            .I(n2320));
    InMux I__4130 (
            .O(N__30853),
            .I(N__30849));
    CascadeMux I__4129 (
            .O(N__30852),
            .I(N__30846));
    LocalMux I__4128 (
            .O(N__30849),
            .I(N__30843));
    InMux I__4127 (
            .O(N__30846),
            .I(N__30840));
    Span4Mux_v I__4126 (
            .O(N__30843),
            .I(N__30837));
    LocalMux I__4125 (
            .O(N__30840),
            .I(r_Tx_Data_5));
    Odrv4 I__4124 (
            .O(N__30837),
            .I(r_Tx_Data_5));
    InMux I__4123 (
            .O(N__30832),
            .I(N__30829));
    LocalMux I__4122 (
            .O(N__30829),
            .I(N__30825));
    InMux I__4121 (
            .O(N__30828),
            .I(N__30822));
    Span4Mux_h I__4120 (
            .O(N__30825),
            .I(N__30819));
    LocalMux I__4119 (
            .O(N__30822),
            .I(data_out_frame_9_4));
    Odrv4 I__4118 (
            .O(N__30819),
            .I(data_out_frame_9_4));
    InMux I__4117 (
            .O(N__30814),
            .I(N__30810));
    InMux I__4116 (
            .O(N__30813),
            .I(N__30807));
    LocalMux I__4115 (
            .O(N__30810),
            .I(data_out_frame_8_4));
    LocalMux I__4114 (
            .O(N__30807),
            .I(data_out_frame_8_4));
    InMux I__4113 (
            .O(N__30802),
            .I(N__30799));
    LocalMux I__4112 (
            .O(N__30799),
            .I(N__30796));
    Span4Mux_v I__4111 (
            .O(N__30796),
            .I(N__30793));
    Odrv4 I__4110 (
            .O(N__30793),
            .I(\c0.n21287 ));
    CascadeMux I__4109 (
            .O(N__30790),
            .I(N__30787));
    InMux I__4108 (
            .O(N__30787),
            .I(N__30783));
    InMux I__4107 (
            .O(N__30786),
            .I(N__30779));
    LocalMux I__4106 (
            .O(N__30783),
            .I(N__30776));
    InMux I__4105 (
            .O(N__30782),
            .I(N__30773));
    LocalMux I__4104 (
            .O(N__30779),
            .I(N__30768));
    Span4Mux_h I__4103 (
            .O(N__30776),
            .I(N__30768));
    LocalMux I__4102 (
            .O(N__30773),
            .I(encoder0_position_9));
    Odrv4 I__4101 (
            .O(N__30768),
            .I(encoder0_position_9));
    InMux I__4100 (
            .O(N__30763),
            .I(N__30759));
    CascadeMux I__4099 (
            .O(N__30762),
            .I(N__30756));
    LocalMux I__4098 (
            .O(N__30759),
            .I(N__30753));
    InMux I__4097 (
            .O(N__30756),
            .I(N__30749));
    Span4Mux_v I__4096 (
            .O(N__30753),
            .I(N__30746));
    InMux I__4095 (
            .O(N__30752),
            .I(N__30743));
    LocalMux I__4094 (
            .O(N__30749),
            .I(encoder1_position_24));
    Odrv4 I__4093 (
            .O(N__30746),
            .I(encoder1_position_24));
    LocalMux I__4092 (
            .O(N__30743),
            .I(encoder1_position_24));
    CascadeMux I__4091 (
            .O(N__30736),
            .I(N__30732));
    InMux I__4090 (
            .O(N__30735),
            .I(N__30729));
    InMux I__4089 (
            .O(N__30732),
            .I(N__30726));
    LocalMux I__4088 (
            .O(N__30729),
            .I(\c0.data_out_frame_0_4 ));
    LocalMux I__4087 (
            .O(N__30726),
            .I(\c0.data_out_frame_0_4 ));
    CascadeMux I__4086 (
            .O(N__30721),
            .I(N__30718));
    InMux I__4085 (
            .O(N__30718),
            .I(N__30715));
    LocalMux I__4084 (
            .O(N__30715),
            .I(N__30710));
    InMux I__4083 (
            .O(N__30714),
            .I(N__30707));
    InMux I__4082 (
            .O(N__30713),
            .I(N__30704));
    Span4Mux_h I__4081 (
            .O(N__30710),
            .I(N__30701));
    LocalMux I__4080 (
            .O(N__30707),
            .I(encoder0_position_8));
    LocalMux I__4079 (
            .O(N__30704),
            .I(encoder0_position_8));
    Odrv4 I__4078 (
            .O(N__30701),
            .I(encoder0_position_8));
    InMux I__4077 (
            .O(N__30694),
            .I(N__30691));
    LocalMux I__4076 (
            .O(N__30691),
            .I(n2319));
    InMux I__4075 (
            .O(N__30688),
            .I(\quad_counter1.n17340 ));
    InMux I__4074 (
            .O(N__30685),
            .I(N__30681));
    CascadeMux I__4073 (
            .O(N__30684),
            .I(N__30677));
    LocalMux I__4072 (
            .O(N__30681),
            .I(N__30674));
    InMux I__4071 (
            .O(N__30680),
            .I(N__30671));
    InMux I__4070 (
            .O(N__30677),
            .I(N__30668));
    Odrv12 I__4069 (
            .O(N__30674),
            .I(encoder1_position_27));
    LocalMux I__4068 (
            .O(N__30671),
            .I(encoder1_position_27));
    LocalMux I__4067 (
            .O(N__30668),
            .I(encoder1_position_27));
    InMux I__4066 (
            .O(N__30661),
            .I(N__30658));
    LocalMux I__4065 (
            .O(N__30658),
            .I(n2318));
    InMux I__4064 (
            .O(N__30655),
            .I(\quad_counter1.n17341 ));
    InMux I__4063 (
            .O(N__30652),
            .I(\quad_counter1.n17342 ));
    InMux I__4062 (
            .O(N__30649),
            .I(\quad_counter1.n17343 ));
    InMux I__4061 (
            .O(N__30646),
            .I(N__30643));
    LocalMux I__4060 (
            .O(N__30643),
            .I(N__30639));
    InMux I__4059 (
            .O(N__30642),
            .I(N__30635));
    Span4Mux_v I__4058 (
            .O(N__30639),
            .I(N__30632));
    InMux I__4057 (
            .O(N__30638),
            .I(N__30629));
    LocalMux I__4056 (
            .O(N__30635),
            .I(N__30626));
    Span4Mux_v I__4055 (
            .O(N__30632),
            .I(N__30619));
    LocalMux I__4054 (
            .O(N__30629),
            .I(N__30619));
    Span4Mux_v I__4053 (
            .O(N__30626),
            .I(N__30619));
    Odrv4 I__4052 (
            .O(N__30619),
            .I(encoder1_position_30));
    InMux I__4051 (
            .O(N__30616),
            .I(N__30613));
    LocalMux I__4050 (
            .O(N__30613),
            .I(N__30610));
    Span4Mux_h I__4049 (
            .O(N__30610),
            .I(N__30607));
    Odrv4 I__4048 (
            .O(N__30607),
            .I(n2315));
    InMux I__4047 (
            .O(N__30604),
            .I(\quad_counter1.n17344 ));
    CascadeMux I__4046 (
            .O(N__30601),
            .I(N__30594));
    CascadeMux I__4045 (
            .O(N__30600),
            .I(N__30590));
    CascadeMux I__4044 (
            .O(N__30599),
            .I(N__30586));
    CascadeMux I__4043 (
            .O(N__30598),
            .I(N__30582));
    InMux I__4042 (
            .O(N__30597),
            .I(N__30561));
    InMux I__4041 (
            .O(N__30594),
            .I(N__30544));
    InMux I__4040 (
            .O(N__30593),
            .I(N__30544));
    InMux I__4039 (
            .O(N__30590),
            .I(N__30544));
    InMux I__4038 (
            .O(N__30589),
            .I(N__30544));
    InMux I__4037 (
            .O(N__30586),
            .I(N__30544));
    InMux I__4036 (
            .O(N__30585),
            .I(N__30544));
    InMux I__4035 (
            .O(N__30582),
            .I(N__30544));
    InMux I__4034 (
            .O(N__30581),
            .I(N__30544));
    InMux I__4033 (
            .O(N__30580),
            .I(N__30535));
    InMux I__4032 (
            .O(N__30579),
            .I(N__30535));
    InMux I__4031 (
            .O(N__30578),
            .I(N__30535));
    InMux I__4030 (
            .O(N__30577),
            .I(N__30535));
    InMux I__4029 (
            .O(N__30576),
            .I(N__30526));
    InMux I__4028 (
            .O(N__30575),
            .I(N__30526));
    InMux I__4027 (
            .O(N__30574),
            .I(N__30526));
    InMux I__4026 (
            .O(N__30573),
            .I(N__30526));
    InMux I__4025 (
            .O(N__30572),
            .I(N__30517));
    InMux I__4024 (
            .O(N__30571),
            .I(N__30517));
    InMux I__4023 (
            .O(N__30570),
            .I(N__30517));
    InMux I__4022 (
            .O(N__30569),
            .I(N__30517));
    InMux I__4021 (
            .O(N__30568),
            .I(N__30508));
    InMux I__4020 (
            .O(N__30567),
            .I(N__30508));
    InMux I__4019 (
            .O(N__30566),
            .I(N__30508));
    InMux I__4018 (
            .O(N__30565),
            .I(N__30508));
    CascadeMux I__4017 (
            .O(N__30564),
            .I(N__30502));
    LocalMux I__4016 (
            .O(N__30561),
            .I(N__30493));
    LocalMux I__4015 (
            .O(N__30544),
            .I(N__30493));
    LocalMux I__4014 (
            .O(N__30535),
            .I(N__30484));
    LocalMux I__4013 (
            .O(N__30526),
            .I(N__30484));
    LocalMux I__4012 (
            .O(N__30517),
            .I(N__30484));
    LocalMux I__4011 (
            .O(N__30508),
            .I(N__30484));
    InMux I__4010 (
            .O(N__30507),
            .I(N__30475));
    InMux I__4009 (
            .O(N__30506),
            .I(N__30475));
    InMux I__4008 (
            .O(N__30505),
            .I(N__30475));
    InMux I__4007 (
            .O(N__30502),
            .I(N__30475));
    InMux I__4006 (
            .O(N__30501),
            .I(N__30466));
    InMux I__4005 (
            .O(N__30500),
            .I(N__30466));
    InMux I__4004 (
            .O(N__30499),
            .I(N__30466));
    InMux I__4003 (
            .O(N__30498),
            .I(N__30466));
    Odrv12 I__4002 (
            .O(N__30493),
            .I(\quad_counter1.n2301 ));
    Odrv4 I__4001 (
            .O(N__30484),
            .I(\quad_counter1.n2301 ));
    LocalMux I__4000 (
            .O(N__30475),
            .I(\quad_counter1.n2301 ));
    LocalMux I__3999 (
            .O(N__30466),
            .I(\quad_counter1.n2301 ));
    InMux I__3998 (
            .O(N__30457),
            .I(bfn_13_13_0_));
    InMux I__3997 (
            .O(N__30454),
            .I(N__30451));
    LocalMux I__3996 (
            .O(N__30451),
            .I(n2314));
    InMux I__3995 (
            .O(N__30448),
            .I(N__30445));
    LocalMux I__3994 (
            .O(N__30445),
            .I(N__30442));
    Odrv12 I__3993 (
            .O(N__30442),
            .I(n2345));
    InMux I__3992 (
            .O(N__30439),
            .I(N__30435));
    InMux I__3991 (
            .O(N__30438),
            .I(N__30432));
    LocalMux I__3990 (
            .O(N__30435),
            .I(data_out_frame_12_5));
    LocalMux I__3989 (
            .O(N__30432),
            .I(data_out_frame_12_5));
    InMux I__3988 (
            .O(N__30427),
            .I(N__30424));
    LocalMux I__3987 (
            .O(N__30424),
            .I(N__30421));
    Odrv4 I__3986 (
            .O(N__30421),
            .I(n2327));
    InMux I__3985 (
            .O(N__30418),
            .I(\quad_counter1.n17332 ));
    CascadeMux I__3984 (
            .O(N__30415),
            .I(N__30412));
    InMux I__3983 (
            .O(N__30412),
            .I(N__30408));
    InMux I__3982 (
            .O(N__30411),
            .I(N__30404));
    LocalMux I__3981 (
            .O(N__30408),
            .I(N__30401));
    InMux I__3980 (
            .O(N__30407),
            .I(N__30398));
    LocalMux I__3979 (
            .O(N__30404),
            .I(N__30393));
    Span4Mux_h I__3978 (
            .O(N__30401),
            .I(N__30393));
    LocalMux I__3977 (
            .O(N__30398),
            .I(encoder1_position_19));
    Odrv4 I__3976 (
            .O(N__30393),
            .I(encoder1_position_19));
    InMux I__3975 (
            .O(N__30388),
            .I(N__30385));
    LocalMux I__3974 (
            .O(N__30385),
            .I(N__30382));
    Span4Mux_v I__3973 (
            .O(N__30382),
            .I(N__30379));
    Odrv4 I__3972 (
            .O(N__30379),
            .I(n2326));
    InMux I__3971 (
            .O(N__30376),
            .I(\quad_counter1.n17333 ));
    InMux I__3970 (
            .O(N__30373),
            .I(N__30369));
    CascadeMux I__3969 (
            .O(N__30372),
            .I(N__30365));
    LocalMux I__3968 (
            .O(N__30369),
            .I(N__30362));
    InMux I__3967 (
            .O(N__30368),
            .I(N__30359));
    InMux I__3966 (
            .O(N__30365),
            .I(N__30356));
    Odrv4 I__3965 (
            .O(N__30362),
            .I(encoder1_position_20));
    LocalMux I__3964 (
            .O(N__30359),
            .I(encoder1_position_20));
    LocalMux I__3963 (
            .O(N__30356),
            .I(encoder1_position_20));
    InMux I__3962 (
            .O(N__30349),
            .I(N__30346));
    LocalMux I__3961 (
            .O(N__30346),
            .I(n2325));
    InMux I__3960 (
            .O(N__30343),
            .I(\quad_counter1.n17334 ));
    InMux I__3959 (
            .O(N__30340),
            .I(\quad_counter1.n17335 ));
    CascadeMux I__3958 (
            .O(N__30337),
            .I(N__30332));
    InMux I__3957 (
            .O(N__30336),
            .I(N__30329));
    InMux I__3956 (
            .O(N__30335),
            .I(N__30326));
    InMux I__3955 (
            .O(N__30332),
            .I(N__30323));
    LocalMux I__3954 (
            .O(N__30329),
            .I(encoder1_position_22));
    LocalMux I__3953 (
            .O(N__30326),
            .I(encoder1_position_22));
    LocalMux I__3952 (
            .O(N__30323),
            .I(encoder1_position_22));
    InMux I__3951 (
            .O(N__30316),
            .I(N__30313));
    LocalMux I__3950 (
            .O(N__30313),
            .I(n2323));
    InMux I__3949 (
            .O(N__30310),
            .I(\quad_counter1.n17336 ));
    InMux I__3948 (
            .O(N__30307),
            .I(bfn_13_12_0_));
    InMux I__3947 (
            .O(N__30304),
            .I(N__30301));
    LocalMux I__3946 (
            .O(N__30301),
            .I(n2321));
    InMux I__3945 (
            .O(N__30298),
            .I(\quad_counter1.n17338 ));
    InMux I__3944 (
            .O(N__30295),
            .I(\quad_counter1.n17339 ));
    InMux I__3943 (
            .O(N__30292),
            .I(N__30288));
    CascadeMux I__3942 (
            .O(N__30291),
            .I(N__30284));
    LocalMux I__3941 (
            .O(N__30288),
            .I(N__30281));
    InMux I__3940 (
            .O(N__30287),
            .I(N__30278));
    InMux I__3939 (
            .O(N__30284),
            .I(N__30275));
    Odrv12 I__3938 (
            .O(N__30281),
            .I(encoder1_position_10));
    LocalMux I__3937 (
            .O(N__30278),
            .I(encoder1_position_10));
    LocalMux I__3936 (
            .O(N__30275),
            .I(encoder1_position_10));
    InMux I__3935 (
            .O(N__30268),
            .I(N__30265));
    LocalMux I__3934 (
            .O(N__30265),
            .I(n2335));
    InMux I__3933 (
            .O(N__30262),
            .I(\quad_counter1.n17324 ));
    InMux I__3932 (
            .O(N__30259),
            .I(N__30256));
    LocalMux I__3931 (
            .O(N__30256),
            .I(N__30252));
    CascadeMux I__3930 (
            .O(N__30255),
            .I(N__30248));
    Span4Mux_v I__3929 (
            .O(N__30252),
            .I(N__30245));
    InMux I__3928 (
            .O(N__30251),
            .I(N__30242));
    InMux I__3927 (
            .O(N__30248),
            .I(N__30239));
    Odrv4 I__3926 (
            .O(N__30245),
            .I(encoder1_position_11));
    LocalMux I__3925 (
            .O(N__30242),
            .I(encoder1_position_11));
    LocalMux I__3924 (
            .O(N__30239),
            .I(encoder1_position_11));
    InMux I__3923 (
            .O(N__30232),
            .I(N__30229));
    LocalMux I__3922 (
            .O(N__30229),
            .I(n2334));
    InMux I__3921 (
            .O(N__30226),
            .I(\quad_counter1.n17325 ));
    InMux I__3920 (
            .O(N__30223),
            .I(\quad_counter1.n17326 ));
    InMux I__3919 (
            .O(N__30220),
            .I(N__30215));
    CascadeMux I__3918 (
            .O(N__30219),
            .I(N__30212));
    InMux I__3917 (
            .O(N__30218),
            .I(N__30209));
    LocalMux I__3916 (
            .O(N__30215),
            .I(N__30206));
    InMux I__3915 (
            .O(N__30212),
            .I(N__30203));
    LocalMux I__3914 (
            .O(N__30209),
            .I(encoder1_position_13));
    Odrv4 I__3913 (
            .O(N__30206),
            .I(encoder1_position_13));
    LocalMux I__3912 (
            .O(N__30203),
            .I(encoder1_position_13));
    InMux I__3911 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__3910 (
            .O(N__30193),
            .I(n2332));
    InMux I__3909 (
            .O(N__30190),
            .I(\quad_counter1.n17327 ));
    InMux I__3908 (
            .O(N__30187),
            .I(N__30182));
    CascadeMux I__3907 (
            .O(N__30186),
            .I(N__30179));
    InMux I__3906 (
            .O(N__30185),
            .I(N__30176));
    LocalMux I__3905 (
            .O(N__30182),
            .I(N__30173));
    InMux I__3904 (
            .O(N__30179),
            .I(N__30170));
    LocalMux I__3903 (
            .O(N__30176),
            .I(encoder1_position_14));
    Odrv4 I__3902 (
            .O(N__30173),
            .I(encoder1_position_14));
    LocalMux I__3901 (
            .O(N__30170),
            .I(encoder1_position_14));
    InMux I__3900 (
            .O(N__30163),
            .I(N__30160));
    LocalMux I__3899 (
            .O(N__30160),
            .I(n2331));
    InMux I__3898 (
            .O(N__30157),
            .I(\quad_counter1.n17328 ));
    InMux I__3897 (
            .O(N__30154),
            .I(N__30150));
    CascadeMux I__3896 (
            .O(N__30153),
            .I(N__30146));
    LocalMux I__3895 (
            .O(N__30150),
            .I(N__30143));
    InMux I__3894 (
            .O(N__30149),
            .I(N__30140));
    InMux I__3893 (
            .O(N__30146),
            .I(N__30137));
    Odrv12 I__3892 (
            .O(N__30143),
            .I(encoder1_position_15));
    LocalMux I__3891 (
            .O(N__30140),
            .I(encoder1_position_15));
    LocalMux I__3890 (
            .O(N__30137),
            .I(encoder1_position_15));
    InMux I__3889 (
            .O(N__30130),
            .I(N__30127));
    LocalMux I__3888 (
            .O(N__30127),
            .I(n2330));
    InMux I__3887 (
            .O(N__30124),
            .I(bfn_13_11_0_));
    InMux I__3886 (
            .O(N__30121),
            .I(N__30118));
    LocalMux I__3885 (
            .O(N__30118),
            .I(N__30113));
    CascadeMux I__3884 (
            .O(N__30117),
            .I(N__30110));
    InMux I__3883 (
            .O(N__30116),
            .I(N__30107));
    Span4Mux_h I__3882 (
            .O(N__30113),
            .I(N__30104));
    InMux I__3881 (
            .O(N__30110),
            .I(N__30101));
    LocalMux I__3880 (
            .O(N__30107),
            .I(encoder1_position_16));
    Odrv4 I__3879 (
            .O(N__30104),
            .I(encoder1_position_16));
    LocalMux I__3878 (
            .O(N__30101),
            .I(encoder1_position_16));
    InMux I__3877 (
            .O(N__30094),
            .I(N__30091));
    LocalMux I__3876 (
            .O(N__30091),
            .I(n2329));
    InMux I__3875 (
            .O(N__30088),
            .I(\quad_counter1.n17330 ));
    InMux I__3874 (
            .O(N__30085),
            .I(N__30082));
    LocalMux I__3873 (
            .O(N__30082),
            .I(n2328));
    InMux I__3872 (
            .O(N__30079),
            .I(\quad_counter1.n17331 ));
    InMux I__3871 (
            .O(N__30076),
            .I(\quad_counter1.n17315 ));
    InMux I__3870 (
            .O(N__30073),
            .I(N__30070));
    LocalMux I__3869 (
            .O(N__30070),
            .I(N__30067));
    Span4Mux_v I__3868 (
            .O(N__30067),
            .I(N__30064));
    Odrv4 I__3867 (
            .O(N__30064),
            .I(n2343));
    InMux I__3866 (
            .O(N__30061),
            .I(\quad_counter1.n17316 ));
    InMux I__3865 (
            .O(N__30058),
            .I(\quad_counter1.n17317 ));
    InMux I__3864 (
            .O(N__30055),
            .I(N__30052));
    LocalMux I__3863 (
            .O(N__30052),
            .I(N__30049));
    Span4Mux_h I__3862 (
            .O(N__30049),
            .I(N__30046));
    Odrv4 I__3861 (
            .O(N__30046),
            .I(n2341));
    InMux I__3860 (
            .O(N__30043),
            .I(\quad_counter1.n17318 ));
    InMux I__3859 (
            .O(N__30040),
            .I(\quad_counter1.n17319 ));
    CascadeMux I__3858 (
            .O(N__30037),
            .I(N__30034));
    InMux I__3857 (
            .O(N__30034),
            .I(N__30030));
    InMux I__3856 (
            .O(N__30033),
            .I(N__30026));
    LocalMux I__3855 (
            .O(N__30030),
            .I(N__30023));
    InMux I__3854 (
            .O(N__30029),
            .I(N__30020));
    LocalMux I__3853 (
            .O(N__30026),
            .I(N__30017));
    Span4Mux_h I__3852 (
            .O(N__30023),
            .I(N__30014));
    LocalMux I__3851 (
            .O(N__30020),
            .I(encoder1_position_6));
    Odrv12 I__3850 (
            .O(N__30017),
            .I(encoder1_position_6));
    Odrv4 I__3849 (
            .O(N__30014),
            .I(encoder1_position_6));
    InMux I__3848 (
            .O(N__30007),
            .I(N__30004));
    LocalMux I__3847 (
            .O(N__30004),
            .I(N__30001));
    Span4Mux_v I__3846 (
            .O(N__30001),
            .I(N__29998));
    Odrv4 I__3845 (
            .O(N__29998),
            .I(n2339));
    InMux I__3844 (
            .O(N__29995),
            .I(\quad_counter1.n17320 ));
    CascadeMux I__3843 (
            .O(N__29992),
            .I(N__29988));
    InMux I__3842 (
            .O(N__29991),
            .I(N__29985));
    InMux I__3841 (
            .O(N__29988),
            .I(N__29982));
    LocalMux I__3840 (
            .O(N__29985),
            .I(N__29979));
    LocalMux I__3839 (
            .O(N__29982),
            .I(N__29975));
    Span4Mux_v I__3838 (
            .O(N__29979),
            .I(N__29972));
    InMux I__3837 (
            .O(N__29978),
            .I(N__29969));
    Span4Mux_h I__3836 (
            .O(N__29975),
            .I(N__29966));
    Odrv4 I__3835 (
            .O(N__29972),
            .I(encoder1_position_7));
    LocalMux I__3834 (
            .O(N__29969),
            .I(encoder1_position_7));
    Odrv4 I__3833 (
            .O(N__29966),
            .I(encoder1_position_7));
    InMux I__3832 (
            .O(N__29959),
            .I(N__29956));
    LocalMux I__3831 (
            .O(N__29956),
            .I(N__29953));
    Span4Mux_h I__3830 (
            .O(N__29953),
            .I(N__29950));
    Odrv4 I__3829 (
            .O(N__29950),
            .I(n2338));
    InMux I__3828 (
            .O(N__29947),
            .I(bfn_13_10_0_));
    InMux I__3827 (
            .O(N__29944),
            .I(N__29941));
    LocalMux I__3826 (
            .O(N__29941),
            .I(N__29938));
    Span4Mux_h I__3825 (
            .O(N__29938),
            .I(N__29935));
    Odrv4 I__3824 (
            .O(N__29935),
            .I(n2337));
    InMux I__3823 (
            .O(N__29932),
            .I(\quad_counter1.n17322 ));
    InMux I__3822 (
            .O(N__29929),
            .I(N__29926));
    LocalMux I__3821 (
            .O(N__29926),
            .I(n2336));
    InMux I__3820 (
            .O(N__29923),
            .I(\quad_counter1.n17323 ));
    InMux I__3819 (
            .O(N__29920),
            .I(N__29917));
    LocalMux I__3818 (
            .O(N__29917),
            .I(\quad_counter1.A_delayed ));
    InMux I__3817 (
            .O(N__29914),
            .I(N__29910));
    InMux I__3816 (
            .O(N__29913),
            .I(N__29907));
    LocalMux I__3815 (
            .O(N__29910),
            .I(N__29904));
    LocalMux I__3814 (
            .O(N__29907),
            .I(N__29900));
    Span4Mux_h I__3813 (
            .O(N__29904),
            .I(N__29897));
    InMux I__3812 (
            .O(N__29903),
            .I(N__29894));
    Span4Mux_h I__3811 (
            .O(N__29900),
            .I(N__29891));
    Odrv4 I__3810 (
            .O(N__29897),
            .I(B_filtered_adj_3582));
    LocalMux I__3809 (
            .O(N__29894),
            .I(B_filtered_adj_3582));
    Odrv4 I__3808 (
            .O(N__29891),
            .I(B_filtered_adj_3582));
    InMux I__3807 (
            .O(N__29884),
            .I(N__29879));
    InMux I__3806 (
            .O(N__29883),
            .I(N__29874));
    InMux I__3805 (
            .O(N__29882),
            .I(N__29874));
    LocalMux I__3804 (
            .O(N__29879),
            .I(\quad_counter1.B_delayed ));
    LocalMux I__3803 (
            .O(N__29874),
            .I(\quad_counter1.B_delayed ));
    CascadeMux I__3802 (
            .O(N__29869),
            .I(N__29863));
    InMux I__3801 (
            .O(N__29868),
            .I(N__29858));
    InMux I__3800 (
            .O(N__29867),
            .I(N__29858));
    InMux I__3799 (
            .O(N__29866),
            .I(N__29852));
    InMux I__3798 (
            .O(N__29863),
            .I(N__29852));
    LocalMux I__3797 (
            .O(N__29858),
            .I(N__29849));
    InMux I__3796 (
            .O(N__29857),
            .I(N__29846));
    LocalMux I__3795 (
            .O(N__29852),
            .I(N__29843));
    Span4Mux_h I__3794 (
            .O(N__29849),
            .I(N__29840));
    LocalMux I__3793 (
            .O(N__29846),
            .I(A_filtered_adj_3581));
    Odrv4 I__3792 (
            .O(N__29843),
            .I(A_filtered_adj_3581));
    Odrv4 I__3791 (
            .O(N__29840),
            .I(A_filtered_adj_3581));
    InMux I__3790 (
            .O(N__29833),
            .I(N__29830));
    LocalMux I__3789 (
            .O(N__29830),
            .I(\quad_counter1.count_direction ));
    InMux I__3788 (
            .O(N__29827),
            .I(\quad_counter1.n17314 ));
    InMux I__3787 (
            .O(N__29824),
            .I(N__29821));
    LocalMux I__3786 (
            .O(N__29821),
            .I(N__29818));
    Span4Mux_v I__3785 (
            .O(N__29818),
            .I(N__29813));
    InMux I__3784 (
            .O(N__29817),
            .I(N__29810));
    InMux I__3783 (
            .O(N__29816),
            .I(N__29807));
    Span4Mux_h I__3782 (
            .O(N__29813),
            .I(N__29804));
    LocalMux I__3781 (
            .O(N__29810),
            .I(\c0.FRAME_MATCHER_state_27 ));
    LocalMux I__3780 (
            .O(N__29807),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv4 I__3779 (
            .O(N__29804),
            .I(\c0.FRAME_MATCHER_state_27 ));
    InMux I__3778 (
            .O(N__29797),
            .I(N__29793));
    InMux I__3777 (
            .O(N__29796),
            .I(N__29789));
    LocalMux I__3776 (
            .O(N__29793),
            .I(N__29786));
    InMux I__3775 (
            .O(N__29792),
            .I(N__29783));
    LocalMux I__3774 (
            .O(N__29789),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv4 I__3773 (
            .O(N__29786),
            .I(\c0.FRAME_MATCHER_state_19 ));
    LocalMux I__3772 (
            .O(N__29783),
            .I(\c0.FRAME_MATCHER_state_19 ));
    InMux I__3771 (
            .O(N__29776),
            .I(N__29772));
    InMux I__3770 (
            .O(N__29775),
            .I(N__29768));
    LocalMux I__3769 (
            .O(N__29772),
            .I(N__29765));
    InMux I__3768 (
            .O(N__29771),
            .I(N__29762));
    LocalMux I__3767 (
            .O(N__29768),
            .I(N__29759));
    Span4Mux_h I__3766 (
            .O(N__29765),
            .I(N__29756));
    LocalMux I__3765 (
            .O(N__29762),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__3764 (
            .O(N__29759),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__3763 (
            .O(N__29756),
            .I(\c0.FRAME_MATCHER_state_24 ));
    CascadeMux I__3762 (
            .O(N__29749),
            .I(N__29746));
    InMux I__3761 (
            .O(N__29746),
            .I(N__29743));
    LocalMux I__3760 (
            .O(N__29743),
            .I(N__29740));
    Odrv4 I__3759 (
            .O(N__29740),
            .I(\c0.n17_adj_3486 ));
    InMux I__3758 (
            .O(N__29737),
            .I(N__29730));
    InMux I__3757 (
            .O(N__29736),
            .I(N__29730));
    InMux I__3756 (
            .O(N__29735),
            .I(N__29726));
    LocalMux I__3755 (
            .O(N__29730),
            .I(N__29723));
    InMux I__3754 (
            .O(N__29729),
            .I(N__29720));
    LocalMux I__3753 (
            .O(N__29726),
            .I(N__29717));
    Span4Mux_v I__3752 (
            .O(N__29723),
            .I(N__29714));
    LocalMux I__3751 (
            .O(N__29720),
            .I(\c0.FRAME_MATCHER_state_7 ));
    Odrv4 I__3750 (
            .O(N__29717),
            .I(\c0.FRAME_MATCHER_state_7 ));
    Odrv4 I__3749 (
            .O(N__29714),
            .I(\c0.FRAME_MATCHER_state_7 ));
    SRMux I__3748 (
            .O(N__29707),
            .I(N__29704));
    LocalMux I__3747 (
            .O(N__29704),
            .I(N__29701));
    Span4Mux_h I__3746 (
            .O(N__29701),
            .I(N__29698));
    Odrv4 I__3745 (
            .O(N__29698),
            .I(\c0.n18677 ));
    CascadeMux I__3744 (
            .O(N__29695),
            .I(N__29691));
    CascadeMux I__3743 (
            .O(N__29694),
            .I(N__29688));
    InMux I__3742 (
            .O(N__29691),
            .I(N__29684));
    InMux I__3741 (
            .O(N__29688),
            .I(N__29681));
    InMux I__3740 (
            .O(N__29687),
            .I(N__29678));
    LocalMux I__3739 (
            .O(N__29684),
            .I(N__29675));
    LocalMux I__3738 (
            .O(N__29681),
            .I(N__29672));
    LocalMux I__3737 (
            .O(N__29678),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv12 I__3736 (
            .O(N__29675),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__3735 (
            .O(N__29672),
            .I(\c0.FRAME_MATCHER_state_30 ));
    SRMux I__3734 (
            .O(N__29665),
            .I(N__29662));
    LocalMux I__3733 (
            .O(N__29662),
            .I(N__29659));
    Span4Mux_v I__3732 (
            .O(N__29659),
            .I(N__29656));
    Odrv4 I__3731 (
            .O(N__29656),
            .I(\c0.n18601 ));
    CascadeMux I__3730 (
            .O(N__29653),
            .I(\c0.n6_adj_3143_cascade_ ));
    InMux I__3729 (
            .O(N__29650),
            .I(N__29647));
    LocalMux I__3728 (
            .O(N__29647),
            .I(N__29644));
    Span4Mux_v I__3727 (
            .O(N__29644),
            .I(N__29641));
    Sp12to4 I__3726 (
            .O(N__29641),
            .I(N__29638));
    Odrv12 I__3725 (
            .O(N__29638),
            .I(\c0.n4_adj_3227 ));
    CascadeMux I__3724 (
            .O(N__29635),
            .I(N__29632));
    InMux I__3723 (
            .O(N__29632),
            .I(N__29629));
    LocalMux I__3722 (
            .O(N__29629),
            .I(\c0.n19045 ));
    InMux I__3721 (
            .O(N__29626),
            .I(N__29619));
    InMux I__3720 (
            .O(N__29625),
            .I(N__29619));
    InMux I__3719 (
            .O(N__29624),
            .I(N__29615));
    LocalMux I__3718 (
            .O(N__29619),
            .I(N__29612));
    InMux I__3717 (
            .O(N__29618),
            .I(N__29609));
    LocalMux I__3716 (
            .O(N__29615),
            .I(N__29604));
    Span4Mux_v I__3715 (
            .O(N__29612),
            .I(N__29604));
    LocalMux I__3714 (
            .O(N__29609),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__3713 (
            .O(N__29604),
            .I(\c0.FRAME_MATCHER_state_25 ));
    InMux I__3712 (
            .O(N__29599),
            .I(N__29595));
    InMux I__3711 (
            .O(N__29598),
            .I(N__29592));
    LocalMux I__3710 (
            .O(N__29595),
            .I(N__29585));
    LocalMux I__3709 (
            .O(N__29592),
            .I(N__29585));
    InMux I__3708 (
            .O(N__29591),
            .I(N__29582));
    InMux I__3707 (
            .O(N__29590),
            .I(N__29579));
    Span4Mux_h I__3706 (
            .O(N__29585),
            .I(N__29576));
    LocalMux I__3705 (
            .O(N__29582),
            .I(\c0.FRAME_MATCHER_state_28 ));
    LocalMux I__3704 (
            .O(N__29579),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__3703 (
            .O(N__29576),
            .I(\c0.FRAME_MATCHER_state_28 ));
    InMux I__3702 (
            .O(N__29569),
            .I(N__29563));
    InMux I__3701 (
            .O(N__29568),
            .I(N__29563));
    LocalMux I__3700 (
            .O(N__29563),
            .I(\c0.n10_adj_3438 ));
    InMux I__3699 (
            .O(N__29560),
            .I(N__29557));
    LocalMux I__3698 (
            .O(N__29557),
            .I(\c0.n19050 ));
    CascadeMux I__3697 (
            .O(N__29554),
            .I(N__29550));
    InMux I__3696 (
            .O(N__29553),
            .I(N__29545));
    InMux I__3695 (
            .O(N__29550),
            .I(N__29540));
    InMux I__3694 (
            .O(N__29549),
            .I(N__29540));
    InMux I__3693 (
            .O(N__29548),
            .I(N__29537));
    LocalMux I__3692 (
            .O(N__29545),
            .I(N__29532));
    LocalMux I__3691 (
            .O(N__29540),
            .I(N__29532));
    LocalMux I__3690 (
            .O(N__29537),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv12 I__3689 (
            .O(N__29532),
            .I(\c0.FRAME_MATCHER_state_6 ));
    InMux I__3688 (
            .O(N__29527),
            .I(N__29524));
    LocalMux I__3687 (
            .O(N__29524),
            .I(N__29520));
    InMux I__3686 (
            .O(N__29523),
            .I(N__29517));
    Span4Mux_h I__3685 (
            .O(N__29520),
            .I(N__29514));
    LocalMux I__3684 (
            .O(N__29517),
            .I(\c0.n63 ));
    Odrv4 I__3683 (
            .O(N__29514),
            .I(\c0.n63 ));
    InMux I__3682 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__3681 (
            .O(N__29506),
            .I(N__29503));
    Odrv12 I__3680 (
            .O(N__29503),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__3679 (
            .O(N__29500),
            .I(N__29497));
    InMux I__3678 (
            .O(N__29497),
            .I(N__29492));
    InMux I__3677 (
            .O(N__29496),
            .I(N__29489));
    InMux I__3676 (
            .O(N__29495),
            .I(N__29486));
    LocalMux I__3675 (
            .O(N__29492),
            .I(N__29483));
    LocalMux I__3674 (
            .O(N__29489),
            .I(\c0.FRAME_MATCHER_state_16 ));
    LocalMux I__3673 (
            .O(N__29486),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__3672 (
            .O(N__29483),
            .I(\c0.FRAME_MATCHER_state_16 ));
    SRMux I__3671 (
            .O(N__29476),
            .I(N__29473));
    LocalMux I__3670 (
            .O(N__29473),
            .I(\c0.n18659 ));
    InMux I__3669 (
            .O(N__29470),
            .I(N__29466));
    InMux I__3668 (
            .O(N__29469),
            .I(N__29463));
    LocalMux I__3667 (
            .O(N__29466),
            .I(N__29460));
    LocalMux I__3666 (
            .O(N__29463),
            .I(N__29457));
    Odrv12 I__3665 (
            .O(N__29460),
            .I(\c0.n19146 ));
    Odrv4 I__3664 (
            .O(N__29457),
            .I(\c0.n19146 ));
    InMux I__3663 (
            .O(N__29452),
            .I(N__29447));
    InMux I__3662 (
            .O(N__29451),
            .I(N__29442));
    InMux I__3661 (
            .O(N__29450),
            .I(N__29442));
    LocalMux I__3660 (
            .O(N__29447),
            .I(\c0.FRAME_MATCHER_state_3 ));
    LocalMux I__3659 (
            .O(N__29442),
            .I(\c0.FRAME_MATCHER_state_3 ));
    SRMux I__3658 (
            .O(N__29437),
            .I(N__29434));
    LocalMux I__3657 (
            .O(N__29434),
            .I(N__29431));
    Span4Mux_h I__3656 (
            .O(N__29431),
            .I(N__29428));
    Odrv4 I__3655 (
            .O(N__29428),
            .I(\c0.n18633 ));
    InMux I__3654 (
            .O(N__29425),
            .I(N__29420));
    InMux I__3653 (
            .O(N__29424),
            .I(N__29417));
    InMux I__3652 (
            .O(N__29423),
            .I(N__29414));
    LocalMux I__3651 (
            .O(N__29420),
            .I(N__29411));
    LocalMux I__3650 (
            .O(N__29417),
            .I(\c0.FRAME_MATCHER_state_14 ));
    LocalMux I__3649 (
            .O(N__29414),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__3648 (
            .O(N__29411),
            .I(\c0.FRAME_MATCHER_state_14 ));
    InMux I__3647 (
            .O(N__29404),
            .I(N__29401));
    LocalMux I__3646 (
            .O(N__29401),
            .I(N__29398));
    Span4Mux_v I__3645 (
            .O(N__29398),
            .I(N__29393));
    InMux I__3644 (
            .O(N__29397),
            .I(N__29390));
    InMux I__3643 (
            .O(N__29396),
            .I(N__29387));
    Span4Mux_h I__3642 (
            .O(N__29393),
            .I(N__29384));
    LocalMux I__3641 (
            .O(N__29390),
            .I(\c0.FRAME_MATCHER_state_9 ));
    LocalMux I__3640 (
            .O(N__29387),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__3639 (
            .O(N__29384),
            .I(\c0.FRAME_MATCHER_state_9 ));
    InMux I__3638 (
            .O(N__29377),
            .I(N__29374));
    LocalMux I__3637 (
            .O(N__29374),
            .I(\c0.n10_adj_3488 ));
    CascadeMux I__3636 (
            .O(N__29371),
            .I(\c0.n15850_cascade_ ));
    CascadeMux I__3635 (
            .O(N__29368),
            .I(\c0.n11427_cascade_ ));
    InMux I__3634 (
            .O(N__29365),
            .I(N__29362));
    LocalMux I__3633 (
            .O(N__29362),
            .I(N__29359));
    Odrv4 I__3632 (
            .O(N__29359),
            .I(\c0.n16_adj_3484 ));
    InMux I__3631 (
            .O(N__29356),
            .I(N__29351));
    InMux I__3630 (
            .O(N__29355),
            .I(N__29348));
    InMux I__3629 (
            .O(N__29354),
            .I(N__29345));
    LocalMux I__3628 (
            .O(N__29351),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__3627 (
            .O(N__29348),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__3626 (
            .O(N__29345),
            .I(\c0.FRAME_MATCHER_state_31 ));
    CascadeMux I__3625 (
            .O(N__29338),
            .I(\c0.n19045_cascade_ ));
    InMux I__3624 (
            .O(N__29335),
            .I(N__29332));
    LocalMux I__3623 (
            .O(N__29332),
            .I(\c0.n4_adj_3046 ));
    CascadeMux I__3622 (
            .O(N__29329),
            .I(N__29325));
    InMux I__3621 (
            .O(N__29328),
            .I(N__29321));
    InMux I__3620 (
            .O(N__29325),
            .I(N__29316));
    InMux I__3619 (
            .O(N__29324),
            .I(N__29316));
    LocalMux I__3618 (
            .O(N__29321),
            .I(N__29313));
    LocalMux I__3617 (
            .O(N__29316),
            .I(N__29310));
    Odrv4 I__3616 (
            .O(N__29313),
            .I(\c0.n15920 ));
    Odrv4 I__3615 (
            .O(N__29310),
            .I(\c0.n15920 ));
    CascadeMux I__3614 (
            .O(N__29305),
            .I(N__29299));
    InMux I__3613 (
            .O(N__29304),
            .I(N__29295));
    InMux I__3612 (
            .O(N__29303),
            .I(N__29292));
    InMux I__3611 (
            .O(N__29302),
            .I(N__29285));
    InMux I__3610 (
            .O(N__29299),
            .I(N__29285));
    InMux I__3609 (
            .O(N__29298),
            .I(N__29285));
    LocalMux I__3608 (
            .O(N__29295),
            .I(N__29273));
    LocalMux I__3607 (
            .O(N__29292),
            .I(N__29273));
    LocalMux I__3606 (
            .O(N__29285),
            .I(N__29273));
    InMux I__3605 (
            .O(N__29284),
            .I(N__29264));
    InMux I__3604 (
            .O(N__29283),
            .I(N__29264));
    InMux I__3603 (
            .O(N__29282),
            .I(N__29261));
    InMux I__3602 (
            .O(N__29281),
            .I(N__29256));
    InMux I__3601 (
            .O(N__29280),
            .I(N__29256));
    Span4Mux_v I__3600 (
            .O(N__29273),
            .I(N__29253));
    InMux I__3599 (
            .O(N__29272),
            .I(N__29244));
    InMux I__3598 (
            .O(N__29271),
            .I(N__29244));
    InMux I__3597 (
            .O(N__29270),
            .I(N__29244));
    InMux I__3596 (
            .O(N__29269),
            .I(N__29244));
    LocalMux I__3595 (
            .O(N__29264),
            .I(r_SM_Main_1_adj_3592));
    LocalMux I__3594 (
            .O(N__29261),
            .I(r_SM_Main_1_adj_3592));
    LocalMux I__3593 (
            .O(N__29256),
            .I(r_SM_Main_1_adj_3592));
    Odrv4 I__3592 (
            .O(N__29253),
            .I(r_SM_Main_1_adj_3592));
    LocalMux I__3591 (
            .O(N__29244),
            .I(r_SM_Main_1_adj_3592));
    InMux I__3590 (
            .O(N__29233),
            .I(N__29230));
    LocalMux I__3589 (
            .O(N__29230),
            .I(N__29227));
    Odrv4 I__3588 (
            .O(N__29227),
            .I(n4_adj_3580));
    InMux I__3587 (
            .O(N__29224),
            .I(N__29221));
    LocalMux I__3586 (
            .O(N__29221),
            .I(N__29218));
    Odrv4 I__3585 (
            .O(N__29218),
            .I(n9_adj_3591));
    InMux I__3584 (
            .O(N__29215),
            .I(N__29211));
    InMux I__3583 (
            .O(N__29214),
            .I(N__29208));
    LocalMux I__3582 (
            .O(N__29211),
            .I(r_Tx_Data_4));
    LocalMux I__3581 (
            .O(N__29208),
            .I(r_Tx_Data_4));
    CEMux I__3580 (
            .O(N__29203),
            .I(N__29200));
    LocalMux I__3579 (
            .O(N__29200),
            .I(N__29196));
    CEMux I__3578 (
            .O(N__29199),
            .I(N__29193));
    Span4Mux_v I__3577 (
            .O(N__29196),
            .I(N__29190));
    LocalMux I__3576 (
            .O(N__29193),
            .I(N__29187));
    Span4Mux_h I__3575 (
            .O(N__29190),
            .I(N__29183));
    Sp12to4 I__3574 (
            .O(N__29187),
            .I(N__29180));
    InMux I__3573 (
            .O(N__29186),
            .I(N__29177));
    Odrv4 I__3572 (
            .O(N__29183),
            .I(\c0.n12512 ));
    Odrv12 I__3571 (
            .O(N__29180),
            .I(\c0.n12512 ));
    LocalMux I__3570 (
            .O(N__29177),
            .I(\c0.n12512 ));
    CascadeMux I__3569 (
            .O(N__29170),
            .I(N__29165));
    InMux I__3568 (
            .O(N__29169),
            .I(N__29149));
    InMux I__3567 (
            .O(N__29168),
            .I(N__29149));
    InMux I__3566 (
            .O(N__29165),
            .I(N__29149));
    InMux I__3565 (
            .O(N__29164),
            .I(N__29149));
    CascadeMux I__3564 (
            .O(N__29163),
            .I(N__29146));
    InMux I__3563 (
            .O(N__29162),
            .I(N__29139));
    InMux I__3562 (
            .O(N__29161),
            .I(N__29134));
    InMux I__3561 (
            .O(N__29160),
            .I(N__29134));
    InMux I__3560 (
            .O(N__29159),
            .I(N__29129));
    InMux I__3559 (
            .O(N__29158),
            .I(N__29129));
    LocalMux I__3558 (
            .O(N__29149),
            .I(N__29126));
    InMux I__3557 (
            .O(N__29146),
            .I(N__29121));
    InMux I__3556 (
            .O(N__29145),
            .I(N__29121));
    InMux I__3555 (
            .O(N__29144),
            .I(N__29118));
    InMux I__3554 (
            .O(N__29143),
            .I(N__29113));
    InMux I__3553 (
            .O(N__29142),
            .I(N__29113));
    LocalMux I__3552 (
            .O(N__29139),
            .I(N__29108));
    LocalMux I__3551 (
            .O(N__29134),
            .I(N__29108));
    LocalMux I__3550 (
            .O(N__29129),
            .I(N__29105));
    Span4Mux_v I__3549 (
            .O(N__29126),
            .I(N__29102));
    LocalMux I__3548 (
            .O(N__29121),
            .I(\c0.r_SM_Main_0 ));
    LocalMux I__3547 (
            .O(N__29118),
            .I(\c0.r_SM_Main_0 ));
    LocalMux I__3546 (
            .O(N__29113),
            .I(\c0.r_SM_Main_0 ));
    Odrv4 I__3545 (
            .O(N__29108),
            .I(\c0.r_SM_Main_0 ));
    Odrv4 I__3544 (
            .O(N__29105),
            .I(\c0.r_SM_Main_0 ));
    Odrv4 I__3543 (
            .O(N__29102),
            .I(\c0.r_SM_Main_0 ));
    InMux I__3542 (
            .O(N__29089),
            .I(N__29086));
    LocalMux I__3541 (
            .O(N__29086),
            .I(\c0.n19023 ));
    SRMux I__3540 (
            .O(N__29083),
            .I(N__29080));
    LocalMux I__3539 (
            .O(N__29080),
            .I(N__29077));
    Sp12to4 I__3538 (
            .O(N__29077),
            .I(N__29074));
    Odrv12 I__3537 (
            .O(N__29074),
            .I(\c0.n18609 ));
    InMux I__3536 (
            .O(N__29071),
            .I(N__29068));
    LocalMux I__3535 (
            .O(N__29068),
            .I(N__29065));
    Span4Mux_h I__3534 (
            .O(N__29065),
            .I(N__29062));
    Odrv4 I__3533 (
            .O(N__29062),
            .I(\c0.n21456 ));
    InMux I__3532 (
            .O(N__29059),
            .I(N__29052));
    InMux I__3531 (
            .O(N__29058),
            .I(N__29043));
    InMux I__3530 (
            .O(N__29057),
            .I(N__29043));
    InMux I__3529 (
            .O(N__29056),
            .I(N__29043));
    InMux I__3528 (
            .O(N__29055),
            .I(N__29043));
    LocalMux I__3527 (
            .O(N__29052),
            .I(\c0.r_Bit_Index_1 ));
    LocalMux I__3526 (
            .O(N__29043),
            .I(\c0.r_Bit_Index_1 ));
    InMux I__3525 (
            .O(N__29038),
            .I(N__29035));
    LocalMux I__3524 (
            .O(N__29035),
            .I(\c0.n21614 ));
    InMux I__3523 (
            .O(N__29032),
            .I(N__29029));
    LocalMux I__3522 (
            .O(N__29029),
            .I(N__29026));
    Odrv4 I__3521 (
            .O(N__29026),
            .I(\c0.n32 ));
    CascadeMux I__3520 (
            .O(N__29023),
            .I(\c0.n2_adj_3556_cascade_ ));
    InMux I__3519 (
            .O(N__29020),
            .I(N__29017));
    LocalMux I__3518 (
            .O(N__29017),
            .I(\c0.n7_adj_3557 ));
    InMux I__3517 (
            .O(N__29014),
            .I(N__29011));
    LocalMux I__3516 (
            .O(N__29011),
            .I(\c0.n21329 ));
    CascadeMux I__3515 (
            .O(N__29008),
            .I(\c0.n19001_cascade_ ));
    InMux I__3514 (
            .O(N__29005),
            .I(N__29002));
    LocalMux I__3513 (
            .O(N__29002),
            .I(N__28999));
    Span4Mux_v I__3512 (
            .O(N__28999),
            .I(N__28996));
    Odrv4 I__3511 (
            .O(N__28996),
            .I(\c0.n30_adj_3559 ));
    CascadeMux I__3510 (
            .O(N__28993),
            .I(N__28989));
    InMux I__3509 (
            .O(N__28992),
            .I(N__28985));
    InMux I__3508 (
            .O(N__28989),
            .I(N__28980));
    InMux I__3507 (
            .O(N__28988),
            .I(N__28980));
    LocalMux I__3506 (
            .O(N__28985),
            .I(\c0.n12498 ));
    LocalMux I__3505 (
            .O(N__28980),
            .I(\c0.n12498 ));
    InMux I__3504 (
            .O(N__28975),
            .I(N__28972));
    LocalMux I__3503 (
            .O(N__28972),
            .I(\c0.n21577 ));
    CascadeMux I__3502 (
            .O(N__28969),
            .I(n21578_cascade_));
    InMux I__3501 (
            .O(N__28966),
            .I(N__28963));
    LocalMux I__3500 (
            .O(N__28963),
            .I(n21656));
    InMux I__3499 (
            .O(N__28960),
            .I(N__28956));
    InMux I__3498 (
            .O(N__28959),
            .I(N__28953));
    LocalMux I__3497 (
            .O(N__28956),
            .I(N__28950));
    LocalMux I__3496 (
            .O(N__28953),
            .I(data_out_frame_13_7));
    Odrv4 I__3495 (
            .O(N__28950),
            .I(data_out_frame_13_7));
    InMux I__3494 (
            .O(N__28945),
            .I(N__28942));
    LocalMux I__3493 (
            .O(N__28942),
            .I(\c0.n21467 ));
    InMux I__3492 (
            .O(N__28939),
            .I(N__28936));
    LocalMux I__3491 (
            .O(N__28936),
            .I(N__28933));
    Span4Mux_h I__3490 (
            .O(N__28933),
            .I(N__28930));
    Odrv4 I__3489 (
            .O(N__28930),
            .I(\c0.tx.n21330 ));
    InMux I__3488 (
            .O(N__28927),
            .I(N__28924));
    LocalMux I__3487 (
            .O(N__28924),
            .I(n9_adj_3588));
    InMux I__3486 (
            .O(N__28921),
            .I(N__28915));
    InMux I__3485 (
            .O(N__28920),
            .I(N__28915));
    LocalMux I__3484 (
            .O(N__28915),
            .I(r_Tx_Data_6));
    CascadeMux I__3483 (
            .O(N__28912),
            .I(\c0.n9753_cascade_ ));
    InMux I__3482 (
            .O(N__28909),
            .I(N__28905));
    InMux I__3481 (
            .O(N__28908),
            .I(N__28902));
    LocalMux I__3480 (
            .O(N__28905),
            .I(N__28899));
    LocalMux I__3479 (
            .O(N__28902),
            .I(data_out_frame_12_3));
    Odrv4 I__3478 (
            .O(N__28899),
            .I(data_out_frame_12_3));
    CascadeMux I__3477 (
            .O(N__28894),
            .I(N__28891));
    InMux I__3476 (
            .O(N__28891),
            .I(N__28885));
    InMux I__3475 (
            .O(N__28890),
            .I(N__28885));
    LocalMux I__3474 (
            .O(N__28885),
            .I(data_out_frame_13_3));
    InMux I__3473 (
            .O(N__28882),
            .I(N__28878));
    InMux I__3472 (
            .O(N__28881),
            .I(N__28875));
    LocalMux I__3471 (
            .O(N__28878),
            .I(data_out_frame_12_7));
    LocalMux I__3470 (
            .O(N__28875),
            .I(data_out_frame_12_7));
    CascadeMux I__3469 (
            .O(N__28870),
            .I(N__28866));
    InMux I__3468 (
            .O(N__28869),
            .I(N__28863));
    InMux I__3467 (
            .O(N__28866),
            .I(N__28860));
    LocalMux I__3466 (
            .O(N__28863),
            .I(data_out_frame_11_3));
    LocalMux I__3465 (
            .O(N__28860),
            .I(data_out_frame_11_3));
    InMux I__3464 (
            .O(N__28855),
            .I(N__28849));
    InMux I__3463 (
            .O(N__28854),
            .I(N__28849));
    LocalMux I__3462 (
            .O(N__28849),
            .I(data_out_frame_10_3));
    InMux I__3461 (
            .O(N__28846),
            .I(N__28843));
    LocalMux I__3460 (
            .O(N__28843),
            .I(N__28839));
    CascadeMux I__3459 (
            .O(N__28842),
            .I(N__28835));
    Span4Mux_h I__3458 (
            .O(N__28839),
            .I(N__28832));
    InMux I__3457 (
            .O(N__28838),
            .I(N__28829));
    InMux I__3456 (
            .O(N__28835),
            .I(N__28826));
    Span4Mux_v I__3455 (
            .O(N__28832),
            .I(N__28819));
    LocalMux I__3454 (
            .O(N__28829),
            .I(N__28819));
    LocalMux I__3453 (
            .O(N__28826),
            .I(N__28819));
    Odrv4 I__3452 (
            .O(N__28819),
            .I(encoder0_position_12));
    InMux I__3451 (
            .O(N__28816),
            .I(N__28812));
    InMux I__3450 (
            .O(N__28815),
            .I(N__28809));
    LocalMux I__3449 (
            .O(N__28812),
            .I(data_out_frame_13_6));
    LocalMux I__3448 (
            .O(N__28809),
            .I(data_out_frame_13_6));
    InMux I__3447 (
            .O(N__28804),
            .I(N__28801));
    LocalMux I__3446 (
            .O(N__28801),
            .I(\c0.n21301 ));
    InMux I__3445 (
            .O(N__28798),
            .I(N__28795));
    LocalMux I__3444 (
            .O(N__28795),
            .I(N__28792));
    Odrv4 I__3443 (
            .O(N__28792),
            .I(\c0.n21653 ));
    InMux I__3442 (
            .O(N__28789),
            .I(N__28786));
    LocalMux I__3441 (
            .O(N__28786),
            .I(N__28783));
    Span4Mux_h I__3440 (
            .O(N__28783),
            .I(N__28780));
    Odrv4 I__3439 (
            .O(N__28780),
            .I(\c0.n21305 ));
    InMux I__3438 (
            .O(N__28777),
            .I(N__28774));
    LocalMux I__3437 (
            .O(N__28774),
            .I(\c0.n21570 ));
    CascadeMux I__3436 (
            .O(N__28771),
            .I(\c0.n21307_cascade_ ));
    InMux I__3435 (
            .O(N__28768),
            .I(N__28764));
    InMux I__3434 (
            .O(N__28767),
            .I(N__28761));
    LocalMux I__3433 (
            .O(N__28764),
            .I(N__28758));
    LocalMux I__3432 (
            .O(N__28761),
            .I(data_out_frame_11_4));
    Odrv4 I__3431 (
            .O(N__28758),
            .I(data_out_frame_11_4));
    CascadeMux I__3430 (
            .O(N__28753),
            .I(N__28750));
    InMux I__3429 (
            .O(N__28750),
            .I(N__28747));
    LocalMux I__3428 (
            .O(N__28747),
            .I(N__28744));
    Odrv4 I__3427 (
            .O(N__28744),
            .I(\c0.n5_adj_3033 ));
    InMux I__3426 (
            .O(N__28741),
            .I(N__28737));
    InMux I__3425 (
            .O(N__28740),
            .I(N__28734));
    LocalMux I__3424 (
            .O(N__28737),
            .I(N__28731));
    LocalMux I__3423 (
            .O(N__28734),
            .I(data_out_frame_12_6));
    Odrv4 I__3422 (
            .O(N__28731),
            .I(data_out_frame_12_6));
    InMux I__3421 (
            .O(N__28726),
            .I(N__28722));
    InMux I__3420 (
            .O(N__28725),
            .I(N__28718));
    LocalMux I__3419 (
            .O(N__28722),
            .I(N__28715));
    InMux I__3418 (
            .O(N__28721),
            .I(N__28712));
    LocalMux I__3417 (
            .O(N__28718),
            .I(encoder0_position_17));
    Odrv4 I__3416 (
            .O(N__28715),
            .I(encoder0_position_17));
    LocalMux I__3415 (
            .O(N__28712),
            .I(encoder0_position_17));
    InMux I__3414 (
            .O(N__28705),
            .I(N__28701));
    InMux I__3413 (
            .O(N__28704),
            .I(N__28698));
    LocalMux I__3412 (
            .O(N__28701),
            .I(data_out_frame_7_1));
    LocalMux I__3411 (
            .O(N__28698),
            .I(data_out_frame_7_1));
    InMux I__3410 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__3409 (
            .O(N__28690),
            .I(\c0.n6_adj_3324 ));
    InMux I__3408 (
            .O(N__28687),
            .I(N__28684));
    LocalMux I__3407 (
            .O(N__28684),
            .I(N__28681));
    Odrv4 I__3406 (
            .O(N__28681),
            .I(n2250));
    InMux I__3405 (
            .O(N__28678),
            .I(N__28675));
    LocalMux I__3404 (
            .O(N__28675),
            .I(N__28670));
    CascadeMux I__3403 (
            .O(N__28674),
            .I(N__28667));
    InMux I__3402 (
            .O(N__28673),
            .I(N__28664));
    Span4Mux_v I__3401 (
            .O(N__28670),
            .I(N__28661));
    InMux I__3400 (
            .O(N__28667),
            .I(N__28658));
    LocalMux I__3399 (
            .O(N__28664),
            .I(encoder0_position_13));
    Odrv4 I__3398 (
            .O(N__28661),
            .I(encoder0_position_13));
    LocalMux I__3397 (
            .O(N__28658),
            .I(encoder0_position_13));
    CascadeMux I__3396 (
            .O(N__28651),
            .I(N__28648));
    InMux I__3395 (
            .O(N__28648),
            .I(N__28645));
    LocalMux I__3394 (
            .O(N__28645),
            .I(N__28641));
    InMux I__3393 (
            .O(N__28644),
            .I(N__28638));
    Span4Mux_h I__3392 (
            .O(N__28641),
            .I(N__28635));
    LocalMux I__3391 (
            .O(N__28638),
            .I(data_out_frame_11_6));
    Odrv4 I__3390 (
            .O(N__28635),
            .I(data_out_frame_11_6));
    InMux I__3389 (
            .O(N__28630),
            .I(N__28627));
    LocalMux I__3388 (
            .O(N__28627),
            .I(N__28624));
    Span4Mux_v I__3387 (
            .O(N__28624),
            .I(N__28621));
    Odrv4 I__3386 (
            .O(N__28621),
            .I(n2271));
    InMux I__3385 (
            .O(N__28618),
            .I(N__28615));
    LocalMux I__3384 (
            .O(N__28615),
            .I(\c0.n21650 ));
    CascadeMux I__3383 (
            .O(N__28612),
            .I(\c0.n21564_cascade_ ));
    InMux I__3382 (
            .O(N__28609),
            .I(N__28606));
    LocalMux I__3381 (
            .O(N__28606),
            .I(N__28603));
    Span4Mux_h I__3380 (
            .O(N__28603),
            .I(N__28600));
    Odrv4 I__3379 (
            .O(N__28600),
            .I(n2270));
    CascadeMux I__3378 (
            .O(N__28597),
            .I(N__28593));
    InMux I__3377 (
            .O(N__28596),
            .I(N__28590));
    InMux I__3376 (
            .O(N__28593),
            .I(N__28587));
    LocalMux I__3375 (
            .O(N__28590),
            .I(\quad_counter1.a_delay_counter_11 ));
    LocalMux I__3374 (
            .O(N__28587),
            .I(\quad_counter1.a_delay_counter_11 ));
    InMux I__3373 (
            .O(N__28582),
            .I(\quad_counter1.n17262 ));
    InMux I__3372 (
            .O(N__28579),
            .I(N__28575));
    InMux I__3371 (
            .O(N__28578),
            .I(N__28572));
    LocalMux I__3370 (
            .O(N__28575),
            .I(\quad_counter1.a_delay_counter_12 ));
    LocalMux I__3369 (
            .O(N__28572),
            .I(\quad_counter1.a_delay_counter_12 ));
    InMux I__3368 (
            .O(N__28567),
            .I(\quad_counter1.n17263 ));
    InMux I__3367 (
            .O(N__28564),
            .I(N__28560));
    InMux I__3366 (
            .O(N__28563),
            .I(N__28557));
    LocalMux I__3365 (
            .O(N__28560),
            .I(\quad_counter1.a_delay_counter_13 ));
    LocalMux I__3364 (
            .O(N__28557),
            .I(\quad_counter1.a_delay_counter_13 ));
    InMux I__3363 (
            .O(N__28552),
            .I(\quad_counter1.n17264 ));
    InMux I__3362 (
            .O(N__28549),
            .I(N__28545));
    InMux I__3361 (
            .O(N__28548),
            .I(N__28542));
    LocalMux I__3360 (
            .O(N__28545),
            .I(\quad_counter1.a_delay_counter_14 ));
    LocalMux I__3359 (
            .O(N__28542),
            .I(\quad_counter1.a_delay_counter_14 ));
    InMux I__3358 (
            .O(N__28537),
            .I(\quad_counter1.n17265 ));
    InMux I__3357 (
            .O(N__28534),
            .I(\quad_counter1.n17266 ));
    InMux I__3356 (
            .O(N__28531),
            .I(N__28527));
    InMux I__3355 (
            .O(N__28530),
            .I(N__28524));
    LocalMux I__3354 (
            .O(N__28527),
            .I(\quad_counter1.a_delay_counter_15 ));
    LocalMux I__3353 (
            .O(N__28524),
            .I(\quad_counter1.a_delay_counter_15 ));
    CEMux I__3352 (
            .O(N__28519),
            .I(N__28516));
    LocalMux I__3351 (
            .O(N__28516),
            .I(N__28512));
    CEMux I__3350 (
            .O(N__28515),
            .I(N__28509));
    Span4Mux_h I__3349 (
            .O(N__28512),
            .I(N__28505));
    LocalMux I__3348 (
            .O(N__28509),
            .I(N__28502));
    InMux I__3347 (
            .O(N__28508),
            .I(N__28499));
    Odrv4 I__3346 (
            .O(N__28505),
            .I(n12477));
    Odrv4 I__3345 (
            .O(N__28502),
            .I(n12477));
    LocalMux I__3344 (
            .O(N__28499),
            .I(n12477));
    SRMux I__3343 (
            .O(N__28492),
            .I(N__28488));
    SRMux I__3342 (
            .O(N__28491),
            .I(N__28485));
    LocalMux I__3341 (
            .O(N__28488),
            .I(N__28482));
    LocalMux I__3340 (
            .O(N__28485),
            .I(N__28479));
    Odrv12 I__3339 (
            .O(N__28482),
            .I(a_delay_counter_15__N_2916_adj_3589));
    Odrv4 I__3338 (
            .O(N__28479),
            .I(a_delay_counter_15__N_2916_adj_3589));
    InMux I__3337 (
            .O(N__28474),
            .I(N__28470));
    InMux I__3336 (
            .O(N__28473),
            .I(N__28467));
    LocalMux I__3335 (
            .O(N__28470),
            .I(N__28464));
    LocalMux I__3334 (
            .O(N__28467),
            .I(data_out_frame_9_2));
    Odrv4 I__3333 (
            .O(N__28464),
            .I(data_out_frame_9_2));
    InMux I__3332 (
            .O(N__28459),
            .I(N__28455));
    InMux I__3331 (
            .O(N__28458),
            .I(N__28452));
    LocalMux I__3330 (
            .O(N__28455),
            .I(data_out_frame_8_2));
    LocalMux I__3329 (
            .O(N__28452),
            .I(data_out_frame_8_2));
    InMux I__3328 (
            .O(N__28447),
            .I(\quad_counter1.n17253 ));
    InMux I__3327 (
            .O(N__28444),
            .I(N__28440));
    InMux I__3326 (
            .O(N__28443),
            .I(N__28437));
    LocalMux I__3325 (
            .O(N__28440),
            .I(\quad_counter1.a_delay_counter_3 ));
    LocalMux I__3324 (
            .O(N__28437),
            .I(\quad_counter1.a_delay_counter_3 ));
    InMux I__3323 (
            .O(N__28432),
            .I(\quad_counter1.n17254 ));
    InMux I__3322 (
            .O(N__28429),
            .I(N__28425));
    InMux I__3321 (
            .O(N__28428),
            .I(N__28422));
    LocalMux I__3320 (
            .O(N__28425),
            .I(\quad_counter1.a_delay_counter_4 ));
    LocalMux I__3319 (
            .O(N__28422),
            .I(\quad_counter1.a_delay_counter_4 ));
    InMux I__3318 (
            .O(N__28417),
            .I(\quad_counter1.n17255 ));
    InMux I__3317 (
            .O(N__28414),
            .I(N__28410));
    InMux I__3316 (
            .O(N__28413),
            .I(N__28407));
    LocalMux I__3315 (
            .O(N__28410),
            .I(\quad_counter1.a_delay_counter_5 ));
    LocalMux I__3314 (
            .O(N__28407),
            .I(\quad_counter1.a_delay_counter_5 ));
    InMux I__3313 (
            .O(N__28402),
            .I(\quad_counter1.n17256 ));
    InMux I__3312 (
            .O(N__28399),
            .I(N__28395));
    InMux I__3311 (
            .O(N__28398),
            .I(N__28392));
    LocalMux I__3310 (
            .O(N__28395),
            .I(\quad_counter1.a_delay_counter_6 ));
    LocalMux I__3309 (
            .O(N__28392),
            .I(\quad_counter1.a_delay_counter_6 ));
    InMux I__3308 (
            .O(N__28387),
            .I(\quad_counter1.n17257 ));
    InMux I__3307 (
            .O(N__28384),
            .I(N__28380));
    InMux I__3306 (
            .O(N__28383),
            .I(N__28377));
    LocalMux I__3305 (
            .O(N__28380),
            .I(\quad_counter1.a_delay_counter_7 ));
    LocalMux I__3304 (
            .O(N__28377),
            .I(\quad_counter1.a_delay_counter_7 ));
    InMux I__3303 (
            .O(N__28372),
            .I(\quad_counter1.n17258 ));
    CascadeMux I__3302 (
            .O(N__28369),
            .I(N__28365));
    InMux I__3301 (
            .O(N__28368),
            .I(N__28362));
    InMux I__3300 (
            .O(N__28365),
            .I(N__28359));
    LocalMux I__3299 (
            .O(N__28362),
            .I(\quad_counter1.a_delay_counter_8 ));
    LocalMux I__3298 (
            .O(N__28359),
            .I(\quad_counter1.a_delay_counter_8 ));
    InMux I__3297 (
            .O(N__28354),
            .I(bfn_12_9_0_));
    InMux I__3296 (
            .O(N__28351),
            .I(N__28347));
    InMux I__3295 (
            .O(N__28350),
            .I(N__28344));
    LocalMux I__3294 (
            .O(N__28347),
            .I(N__28341));
    LocalMux I__3293 (
            .O(N__28344),
            .I(\quad_counter1.a_delay_counter_9 ));
    Odrv4 I__3292 (
            .O(N__28341),
            .I(\quad_counter1.a_delay_counter_9 ));
    InMux I__3291 (
            .O(N__28336),
            .I(\quad_counter1.n17260 ));
    InMux I__3290 (
            .O(N__28333),
            .I(N__28329));
    InMux I__3289 (
            .O(N__28332),
            .I(N__28326));
    LocalMux I__3288 (
            .O(N__28329),
            .I(\quad_counter1.a_delay_counter_10 ));
    LocalMux I__3287 (
            .O(N__28326),
            .I(\quad_counter1.a_delay_counter_10 ));
    InMux I__3286 (
            .O(N__28321),
            .I(\quad_counter1.n17261 ));
    InMux I__3285 (
            .O(N__28318),
            .I(N__28314));
    InMux I__3284 (
            .O(N__28317),
            .I(N__28311));
    LocalMux I__3283 (
            .O(N__28314),
            .I(\quad_counter1.b_delay_counter_13 ));
    LocalMux I__3282 (
            .O(N__28311),
            .I(\quad_counter1.b_delay_counter_13 ));
    InMux I__3281 (
            .O(N__28306),
            .I(\quad_counter1.n17249 ));
    InMux I__3280 (
            .O(N__28303),
            .I(N__28299));
    InMux I__3279 (
            .O(N__28302),
            .I(N__28296));
    LocalMux I__3278 (
            .O(N__28299),
            .I(\quad_counter1.b_delay_counter_14 ));
    LocalMux I__3277 (
            .O(N__28296),
            .I(\quad_counter1.b_delay_counter_14 ));
    InMux I__3276 (
            .O(N__28291),
            .I(\quad_counter1.n17250 ));
    InMux I__3275 (
            .O(N__28288),
            .I(\quad_counter1.n17251 ));
    InMux I__3274 (
            .O(N__28285),
            .I(N__28281));
    InMux I__3273 (
            .O(N__28284),
            .I(N__28278));
    LocalMux I__3272 (
            .O(N__28281),
            .I(\quad_counter1.b_delay_counter_15 ));
    LocalMux I__3271 (
            .O(N__28278),
            .I(\quad_counter1.b_delay_counter_15 ));
    CEMux I__3270 (
            .O(N__28273),
            .I(N__28270));
    LocalMux I__3269 (
            .O(N__28270),
            .I(N__28267));
    Span4Mux_v I__3268 (
            .O(N__28267),
            .I(N__28263));
    CEMux I__3267 (
            .O(N__28266),
            .I(N__28260));
    Span4Mux_s2_v I__3266 (
            .O(N__28263),
            .I(N__28255));
    LocalMux I__3265 (
            .O(N__28260),
            .I(N__28255));
    Span4Mux_v I__3264 (
            .O(N__28255),
            .I(N__28252));
    Span4Mux_s2_v I__3263 (
            .O(N__28252),
            .I(N__28249));
    Odrv4 I__3262 (
            .O(N__28249),
            .I(n12417));
    SRMux I__3261 (
            .O(N__28246),
            .I(N__28241));
    InMux I__3260 (
            .O(N__28245),
            .I(N__28238));
    SRMux I__3259 (
            .O(N__28244),
            .I(N__28235));
    LocalMux I__3258 (
            .O(N__28241),
            .I(N__28232));
    LocalMux I__3257 (
            .O(N__28238),
            .I(N__28228));
    LocalMux I__3256 (
            .O(N__28235),
            .I(N__28223));
    Span4Mux_v I__3255 (
            .O(N__28232),
            .I(N__28223));
    InMux I__3254 (
            .O(N__28231),
            .I(N__28220));
    Odrv4 I__3253 (
            .O(N__28228),
            .I(b_delay_counter_15__N_2933));
    Odrv4 I__3252 (
            .O(N__28223),
            .I(b_delay_counter_15__N_2933));
    LocalMux I__3251 (
            .O(N__28220),
            .I(b_delay_counter_15__N_2933));
    InMux I__3250 (
            .O(N__28213),
            .I(N__28207));
    InMux I__3249 (
            .O(N__28212),
            .I(N__28207));
    LocalMux I__3248 (
            .O(N__28207),
            .I(N__28202));
    InMux I__3247 (
            .O(N__28206),
            .I(N__28199));
    InMux I__3246 (
            .O(N__28205),
            .I(N__28196));
    Span4Mux_v I__3245 (
            .O(N__28202),
            .I(N__28191));
    LocalMux I__3244 (
            .O(N__28199),
            .I(N__28191));
    LocalMux I__3243 (
            .O(N__28196),
            .I(N__28188));
    IoSpan4Mux I__3242 (
            .O(N__28191),
            .I(N__28185));
    Span12Mux_h I__3241 (
            .O(N__28188),
            .I(N__28182));
    IoSpan4Mux I__3240 (
            .O(N__28185),
            .I(N__28179));
    Odrv12 I__3239 (
            .O(N__28182),
            .I(PIN_12_c));
    Odrv4 I__3238 (
            .O(N__28179),
            .I(PIN_12_c));
    CascadeMux I__3237 (
            .O(N__28174),
            .I(N__28171));
    InMux I__3236 (
            .O(N__28171),
            .I(N__28164));
    InMux I__3235 (
            .O(N__28170),
            .I(N__28164));
    InMux I__3234 (
            .O(N__28169),
            .I(N__28161));
    LocalMux I__3233 (
            .O(N__28164),
            .I(N__28156));
    LocalMux I__3232 (
            .O(N__28161),
            .I(N__28156));
    Span4Mux_h I__3231 (
            .O(N__28156),
            .I(N__28153));
    Odrv4 I__3230 (
            .O(N__28153),
            .I(quadA_delayed_adj_3584));
    CascadeMux I__3229 (
            .O(N__28150),
            .I(a_delay_counter_15__N_2916_adj_3589_cascade_));
    InMux I__3228 (
            .O(N__28147),
            .I(N__28144));
    LocalMux I__3227 (
            .O(N__28144),
            .I(\quad_counter1.n20 ));
    InMux I__3226 (
            .O(N__28141),
            .I(N__28136));
    InMux I__3225 (
            .O(N__28140),
            .I(N__28131));
    InMux I__3224 (
            .O(N__28139),
            .I(N__28131));
    LocalMux I__3223 (
            .O(N__28136),
            .I(a_delay_counter_0_adj_3583));
    LocalMux I__3222 (
            .O(N__28131),
            .I(a_delay_counter_0_adj_3583));
    InMux I__3221 (
            .O(N__28126),
            .I(N__28123));
    LocalMux I__3220 (
            .O(N__28123),
            .I(n39_adj_3587));
    InMux I__3219 (
            .O(N__28120),
            .I(bfn_12_8_0_));
    InMux I__3218 (
            .O(N__28117),
            .I(N__28113));
    InMux I__3217 (
            .O(N__28116),
            .I(N__28110));
    LocalMux I__3216 (
            .O(N__28113),
            .I(\quad_counter1.a_delay_counter_1 ));
    LocalMux I__3215 (
            .O(N__28110),
            .I(\quad_counter1.a_delay_counter_1 ));
    InMux I__3214 (
            .O(N__28105),
            .I(\quad_counter1.n17252 ));
    InMux I__3213 (
            .O(N__28102),
            .I(N__28098));
    InMux I__3212 (
            .O(N__28101),
            .I(N__28095));
    LocalMux I__3211 (
            .O(N__28098),
            .I(\quad_counter1.a_delay_counter_2 ));
    LocalMux I__3210 (
            .O(N__28095),
            .I(\quad_counter1.a_delay_counter_2 ));
    InMux I__3209 (
            .O(N__28090),
            .I(N__28086));
    InMux I__3208 (
            .O(N__28089),
            .I(N__28083));
    LocalMux I__3207 (
            .O(N__28086),
            .I(\quad_counter1.b_delay_counter_5 ));
    LocalMux I__3206 (
            .O(N__28083),
            .I(\quad_counter1.b_delay_counter_5 ));
    InMux I__3205 (
            .O(N__28078),
            .I(\quad_counter1.n17241 ));
    CascadeMux I__3204 (
            .O(N__28075),
            .I(N__28071));
    InMux I__3203 (
            .O(N__28074),
            .I(N__28068));
    InMux I__3202 (
            .O(N__28071),
            .I(N__28065));
    LocalMux I__3201 (
            .O(N__28068),
            .I(\quad_counter1.b_delay_counter_6 ));
    LocalMux I__3200 (
            .O(N__28065),
            .I(\quad_counter1.b_delay_counter_6 ));
    InMux I__3199 (
            .O(N__28060),
            .I(\quad_counter1.n17242 ));
    InMux I__3198 (
            .O(N__28057),
            .I(N__28053));
    InMux I__3197 (
            .O(N__28056),
            .I(N__28050));
    LocalMux I__3196 (
            .O(N__28053),
            .I(\quad_counter1.b_delay_counter_7 ));
    LocalMux I__3195 (
            .O(N__28050),
            .I(\quad_counter1.b_delay_counter_7 ));
    InMux I__3194 (
            .O(N__28045),
            .I(\quad_counter1.n17243 ));
    InMux I__3193 (
            .O(N__28042),
            .I(N__28038));
    InMux I__3192 (
            .O(N__28041),
            .I(N__28035));
    LocalMux I__3191 (
            .O(N__28038),
            .I(\quad_counter1.b_delay_counter_8 ));
    LocalMux I__3190 (
            .O(N__28035),
            .I(\quad_counter1.b_delay_counter_8 ));
    InMux I__3189 (
            .O(N__28030),
            .I(bfn_12_6_0_));
    InMux I__3188 (
            .O(N__28027),
            .I(N__28023));
    InMux I__3187 (
            .O(N__28026),
            .I(N__28020));
    LocalMux I__3186 (
            .O(N__28023),
            .I(\quad_counter1.b_delay_counter_9 ));
    LocalMux I__3185 (
            .O(N__28020),
            .I(\quad_counter1.b_delay_counter_9 ));
    InMux I__3184 (
            .O(N__28015),
            .I(\quad_counter1.n17245 ));
    InMux I__3183 (
            .O(N__28012),
            .I(N__28008));
    InMux I__3182 (
            .O(N__28011),
            .I(N__28005));
    LocalMux I__3181 (
            .O(N__28008),
            .I(\quad_counter1.b_delay_counter_10 ));
    LocalMux I__3180 (
            .O(N__28005),
            .I(\quad_counter1.b_delay_counter_10 ));
    InMux I__3179 (
            .O(N__28000),
            .I(\quad_counter1.n17246 ));
    InMux I__3178 (
            .O(N__27997),
            .I(N__27993));
    InMux I__3177 (
            .O(N__27996),
            .I(N__27990));
    LocalMux I__3176 (
            .O(N__27993),
            .I(\quad_counter1.b_delay_counter_11 ));
    LocalMux I__3175 (
            .O(N__27990),
            .I(\quad_counter1.b_delay_counter_11 ));
    InMux I__3174 (
            .O(N__27985),
            .I(\quad_counter1.n17247 ));
    CascadeMux I__3173 (
            .O(N__27982),
            .I(N__27978));
    InMux I__3172 (
            .O(N__27981),
            .I(N__27975));
    InMux I__3171 (
            .O(N__27978),
            .I(N__27972));
    LocalMux I__3170 (
            .O(N__27975),
            .I(\quad_counter1.b_delay_counter_12 ));
    LocalMux I__3169 (
            .O(N__27972),
            .I(\quad_counter1.b_delay_counter_12 ));
    InMux I__3168 (
            .O(N__27967),
            .I(\quad_counter1.n17248 ));
    SRMux I__3167 (
            .O(N__27964),
            .I(N__27961));
    LocalMux I__3166 (
            .O(N__27961),
            .I(N__27958));
    Span4Mux_h I__3165 (
            .O(N__27958),
            .I(N__27955));
    Odrv4 I__3164 (
            .O(N__27955),
            .I(\c0.n18651 ));
    SRMux I__3163 (
            .O(N__27952),
            .I(N__27949));
    LocalMux I__3162 (
            .O(N__27949),
            .I(N__27946));
    Span4Mux_h I__3161 (
            .O(N__27946),
            .I(N__27943));
    Odrv4 I__3160 (
            .O(N__27943),
            .I(\c0.n18625 ));
    SRMux I__3159 (
            .O(N__27940),
            .I(N__27937));
    LocalMux I__3158 (
            .O(N__27937),
            .I(N__27934));
    Span4Mux_h I__3157 (
            .O(N__27934),
            .I(N__27931));
    Odrv4 I__3156 (
            .O(N__27931),
            .I(\c0.n18641 ));
    InMux I__3155 (
            .O(N__27928),
            .I(N__27923));
    InMux I__3154 (
            .O(N__27927),
            .I(N__27918));
    InMux I__3153 (
            .O(N__27926),
            .I(N__27918));
    LocalMux I__3152 (
            .O(N__27923),
            .I(b_delay_counter_0));
    LocalMux I__3151 (
            .O(N__27918),
            .I(b_delay_counter_0));
    InMux I__3150 (
            .O(N__27913),
            .I(N__27910));
    LocalMux I__3149 (
            .O(N__27910),
            .I(n187));
    InMux I__3148 (
            .O(N__27907),
            .I(bfn_12_5_0_));
    CascadeMux I__3147 (
            .O(N__27904),
            .I(N__27900));
    InMux I__3146 (
            .O(N__27903),
            .I(N__27897));
    InMux I__3145 (
            .O(N__27900),
            .I(N__27894));
    LocalMux I__3144 (
            .O(N__27897),
            .I(\quad_counter1.b_delay_counter_1 ));
    LocalMux I__3143 (
            .O(N__27894),
            .I(\quad_counter1.b_delay_counter_1 ));
    InMux I__3142 (
            .O(N__27889),
            .I(\quad_counter1.n17237 ));
    CascadeMux I__3141 (
            .O(N__27886),
            .I(N__27882));
    InMux I__3140 (
            .O(N__27885),
            .I(N__27879));
    InMux I__3139 (
            .O(N__27882),
            .I(N__27876));
    LocalMux I__3138 (
            .O(N__27879),
            .I(\quad_counter1.b_delay_counter_2 ));
    LocalMux I__3137 (
            .O(N__27876),
            .I(\quad_counter1.b_delay_counter_2 ));
    InMux I__3136 (
            .O(N__27871),
            .I(\quad_counter1.n17238 ));
    InMux I__3135 (
            .O(N__27868),
            .I(N__27864));
    InMux I__3134 (
            .O(N__27867),
            .I(N__27861));
    LocalMux I__3133 (
            .O(N__27864),
            .I(\quad_counter1.b_delay_counter_3 ));
    LocalMux I__3132 (
            .O(N__27861),
            .I(\quad_counter1.b_delay_counter_3 ));
    InMux I__3131 (
            .O(N__27856),
            .I(\quad_counter1.n17239 ));
    InMux I__3130 (
            .O(N__27853),
            .I(N__27849));
    InMux I__3129 (
            .O(N__27852),
            .I(N__27846));
    LocalMux I__3128 (
            .O(N__27849),
            .I(\quad_counter1.b_delay_counter_4 ));
    LocalMux I__3127 (
            .O(N__27846),
            .I(\quad_counter1.b_delay_counter_4 ));
    InMux I__3126 (
            .O(N__27841),
            .I(\quad_counter1.n17240 ));
    SRMux I__3125 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__3124 (
            .O(N__27835),
            .I(N__27832));
    Span4Mux_v I__3123 (
            .O(N__27832),
            .I(N__27829));
    Odrv4 I__3122 (
            .O(N__27829),
            .I(\c0.n18637 ));
    InMux I__3121 (
            .O(N__27826),
            .I(N__27817));
    InMux I__3120 (
            .O(N__27825),
            .I(N__27817));
    InMux I__3119 (
            .O(N__27824),
            .I(N__27817));
    LocalMux I__3118 (
            .O(N__27817),
            .I(\c0.FRAME_MATCHER_state_22 ));
    SRMux I__3117 (
            .O(N__27814),
            .I(N__27811));
    LocalMux I__3116 (
            .O(N__27811),
            .I(N__27808));
    Odrv4 I__3115 (
            .O(N__27808),
            .I(\c0.n18635 ));
    InMux I__3114 (
            .O(N__27805),
            .I(N__27799));
    InMux I__3113 (
            .O(N__27804),
            .I(N__27799));
    LocalMux I__3112 (
            .O(N__27799),
            .I(N__27795));
    InMux I__3111 (
            .O(N__27798),
            .I(N__27792));
    Span4Mux_v I__3110 (
            .O(N__27795),
            .I(N__27789));
    LocalMux I__3109 (
            .O(N__27792),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv4 I__3108 (
            .O(N__27789),
            .I(\c0.FRAME_MATCHER_state_26 ));
    SRMux I__3107 (
            .O(N__27784),
            .I(N__27781));
    LocalMux I__3106 (
            .O(N__27781),
            .I(N__27778));
    Span4Mux_h I__3105 (
            .O(N__27778),
            .I(N__27775));
    Odrv4 I__3104 (
            .O(N__27775),
            .I(\c0.n18623 ));
    InMux I__3103 (
            .O(N__27772),
            .I(N__27767));
    InMux I__3102 (
            .O(N__27771),
            .I(N__27764));
    InMux I__3101 (
            .O(N__27770),
            .I(N__27761));
    LocalMux I__3100 (
            .O(N__27767),
            .I(N__27756));
    LocalMux I__3099 (
            .O(N__27764),
            .I(N__27756));
    LocalMux I__3098 (
            .O(N__27761),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv4 I__3097 (
            .O(N__27756),
            .I(\c0.FRAME_MATCHER_state_13 ));
    SRMux I__3096 (
            .O(N__27751),
            .I(N__27748));
    LocalMux I__3095 (
            .O(N__27748),
            .I(N__27745));
    Span4Mux_h I__3094 (
            .O(N__27745),
            .I(N__27742));
    Odrv4 I__3093 (
            .O(N__27742),
            .I(\c0.n18665 ));
    InMux I__3092 (
            .O(N__27739),
            .I(N__27734));
    InMux I__3091 (
            .O(N__27738),
            .I(N__27731));
    InMux I__3090 (
            .O(N__27737),
            .I(N__27728));
    LocalMux I__3089 (
            .O(N__27734),
            .I(N__27723));
    LocalMux I__3088 (
            .O(N__27731),
            .I(N__27723));
    LocalMux I__3087 (
            .O(N__27728),
            .I(\c0.FRAME_MATCHER_state_23 ));
    Odrv12 I__3086 (
            .O(N__27723),
            .I(\c0.FRAME_MATCHER_state_23 ));
    InMux I__3085 (
            .O(N__27718),
            .I(N__27714));
    CascadeMux I__3084 (
            .O(N__27717),
            .I(N__27711));
    LocalMux I__3083 (
            .O(N__27714),
            .I(N__27707));
    InMux I__3082 (
            .O(N__27711),
            .I(N__27702));
    InMux I__3081 (
            .O(N__27710),
            .I(N__27702));
    Odrv4 I__3080 (
            .O(N__27707),
            .I(\c0.FRAME_MATCHER_state_20 ));
    LocalMux I__3079 (
            .O(N__27702),
            .I(\c0.FRAME_MATCHER_state_20 ));
    InMux I__3078 (
            .O(N__27697),
            .I(N__27694));
    LocalMux I__3077 (
            .O(N__27694),
            .I(\c0.tx.n4 ));
    CascadeMux I__3076 (
            .O(N__27691),
            .I(\c0.tx.n21179_cascade_ ));
    InMux I__3075 (
            .O(N__27688),
            .I(N__27682));
    InMux I__3074 (
            .O(N__27687),
            .I(N__27682));
    LocalMux I__3073 (
            .O(N__27682),
            .I(N__27675));
    InMux I__3072 (
            .O(N__27681),
            .I(N__27672));
    InMux I__3071 (
            .O(N__27680),
            .I(N__27665));
    InMux I__3070 (
            .O(N__27679),
            .I(N__27665));
    InMux I__3069 (
            .O(N__27678),
            .I(N__27665));
    Span4Mux_h I__3068 (
            .O(N__27675),
            .I(N__27662));
    LocalMux I__3067 (
            .O(N__27672),
            .I(\c0.r_Clock_Count_8 ));
    LocalMux I__3066 (
            .O(N__27665),
            .I(\c0.r_Clock_Count_8 ));
    Odrv4 I__3065 (
            .O(N__27662),
            .I(\c0.r_Clock_Count_8 ));
    SRMux I__3064 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__3063 (
            .O(N__27652),
            .I(N__27648));
    SRMux I__3062 (
            .O(N__27651),
            .I(N__27645));
    Span4Mux_h I__3061 (
            .O(N__27648),
            .I(N__27642));
    LocalMux I__3060 (
            .O(N__27645),
            .I(N__27639));
    Odrv4 I__3059 (
            .O(N__27642),
            .I(\c0.tx.n12759 ));
    Odrv4 I__3058 (
            .O(N__27639),
            .I(\c0.tx.n12759 ));
    InMux I__3057 (
            .O(N__27634),
            .I(N__27629));
    InMux I__3056 (
            .O(N__27633),
            .I(N__27626));
    InMux I__3055 (
            .O(N__27632),
            .I(N__27623));
    LocalMux I__3054 (
            .O(N__27629),
            .I(N__27620));
    LocalMux I__3053 (
            .O(N__27626),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__3052 (
            .O(N__27623),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv12 I__3051 (
            .O(N__27620),
            .I(\c0.FRAME_MATCHER_state_15 ));
    CascadeMux I__3050 (
            .O(N__27613),
            .I(N__27608));
    InMux I__3049 (
            .O(N__27612),
            .I(N__27605));
    InMux I__3048 (
            .O(N__27611),
            .I(N__27602));
    InMux I__3047 (
            .O(N__27608),
            .I(N__27599));
    LocalMux I__3046 (
            .O(N__27605),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__3045 (
            .O(N__27602),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__3044 (
            .O(N__27599),
            .I(\c0.FRAME_MATCHER_state_10 ));
    InMux I__3043 (
            .O(N__27592),
            .I(N__27583));
    InMux I__3042 (
            .O(N__27591),
            .I(N__27583));
    InMux I__3041 (
            .O(N__27590),
            .I(N__27583));
    LocalMux I__3040 (
            .O(N__27583),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__3039 (
            .O(N__27580),
            .I(N__27577));
    LocalMux I__3038 (
            .O(N__27577),
            .I(N__27574));
    Span4Mux_h I__3037 (
            .O(N__27574),
            .I(N__27571));
    Odrv4 I__3036 (
            .O(N__27571),
            .I(\c0.n18669 ));
    SRMux I__3035 (
            .O(N__27568),
            .I(N__27565));
    LocalMux I__3034 (
            .O(N__27565),
            .I(N__27562));
    Odrv4 I__3033 (
            .O(N__27562),
            .I(\c0.n18679 ));
    CascadeMux I__3032 (
            .O(N__27559),
            .I(\c0.n21506_cascade_ ));
    InMux I__3031 (
            .O(N__27556),
            .I(N__27552));
    InMux I__3030 (
            .O(N__27555),
            .I(N__27549));
    LocalMux I__3029 (
            .O(N__27552),
            .I(\c0.n55 ));
    LocalMux I__3028 (
            .O(N__27549),
            .I(\c0.n55 ));
    CascadeMux I__3027 (
            .O(N__27544),
            .I(N__27539));
    InMux I__3026 (
            .O(N__27543),
            .I(N__27536));
    InMux I__3025 (
            .O(N__27542),
            .I(N__27531));
    InMux I__3024 (
            .O(N__27539),
            .I(N__27531));
    LocalMux I__3023 (
            .O(N__27536),
            .I(\c0.r_Bit_Index_2 ));
    LocalMux I__3022 (
            .O(N__27531),
            .I(\c0.r_Bit_Index_2 ));
    CascadeMux I__3021 (
            .O(N__27526),
            .I(\c0.n21414_cascade_ ));
    InMux I__3020 (
            .O(N__27523),
            .I(N__27520));
    LocalMux I__3019 (
            .O(N__27520),
            .I(\c0.n11 ));
    InMux I__3018 (
            .O(N__27517),
            .I(N__27511));
    InMux I__3017 (
            .O(N__27516),
            .I(N__27508));
    InMux I__3016 (
            .O(N__27515),
            .I(N__27503));
    InMux I__3015 (
            .O(N__27514),
            .I(N__27503));
    LocalMux I__3014 (
            .O(N__27511),
            .I(\c0.n15938 ));
    LocalMux I__3013 (
            .O(N__27508),
            .I(\c0.n15938 ));
    LocalMux I__3012 (
            .O(N__27503),
            .I(\c0.n15938 ));
    InMux I__3011 (
            .O(N__27496),
            .I(N__27493));
    LocalMux I__3010 (
            .O(N__27493),
            .I(\c0.tx.n8 ));
    CascadeMux I__3009 (
            .O(N__27490),
            .I(\c0.n55_cascade_ ));
    CascadeMux I__3008 (
            .O(N__27487),
            .I(\c0.n14301_cascade_ ));
    InMux I__3007 (
            .O(N__27484),
            .I(N__27481));
    LocalMux I__3006 (
            .O(N__27481),
            .I(\c0.n15942 ));
    InMux I__3005 (
            .O(N__27478),
            .I(N__27475));
    LocalMux I__3004 (
            .O(N__27475),
            .I(n6866));
    InMux I__3003 (
            .O(N__27472),
            .I(N__27468));
    InMux I__3002 (
            .O(N__27471),
            .I(N__27465));
    LocalMux I__3001 (
            .O(N__27468),
            .I(data_out_frame_10_4));
    LocalMux I__3000 (
            .O(N__27465),
            .I(data_out_frame_10_4));
    InMux I__2999 (
            .O(N__27460),
            .I(N__27457));
    LocalMux I__2998 (
            .O(N__27457),
            .I(\c0.n21288 ));
    InMux I__2997 (
            .O(N__27454),
            .I(N__27451));
    LocalMux I__2996 (
            .O(N__27451),
            .I(N__27448));
    Span4Mux_v I__2995 (
            .O(N__27448),
            .I(N__27445));
    Odrv4 I__2994 (
            .O(N__27445),
            .I(n2273));
    CascadeMux I__2993 (
            .O(N__27442),
            .I(N__27439));
    InMux I__2992 (
            .O(N__27439),
            .I(N__27436));
    LocalMux I__2991 (
            .O(N__27436),
            .I(N__27432));
    InMux I__2990 (
            .O(N__27435),
            .I(N__27428));
    Span4Mux_h I__2989 (
            .O(N__27432),
            .I(N__27425));
    InMux I__2988 (
            .O(N__27431),
            .I(N__27422));
    LocalMux I__2987 (
            .O(N__27428),
            .I(N__27417));
    Span4Mux_v I__2986 (
            .O(N__27425),
            .I(N__27417));
    LocalMux I__2985 (
            .O(N__27422),
            .I(encoder0_position_6));
    Odrv4 I__2984 (
            .O(N__27417),
            .I(encoder0_position_6));
    InMux I__2983 (
            .O(N__27412),
            .I(N__27409));
    LocalMux I__2982 (
            .O(N__27409),
            .I(\c0.n21517 ));
    CascadeMux I__2981 (
            .O(N__27406),
            .I(\c0.n21626_cascade_ ));
    CascadeMux I__2980 (
            .O(N__27403),
            .I(N__27399));
    InMux I__2979 (
            .O(N__27402),
            .I(N__27395));
    InMux I__2978 (
            .O(N__27399),
            .I(N__27392));
    InMux I__2977 (
            .O(N__27398),
            .I(N__27389));
    LocalMux I__2976 (
            .O(N__27395),
            .I(N__27386));
    LocalMux I__2975 (
            .O(N__27392),
            .I(N__27383));
    LocalMux I__2974 (
            .O(N__27389),
            .I(encoder0_position_7));
    Odrv4 I__2973 (
            .O(N__27386),
            .I(encoder0_position_7));
    Odrv4 I__2972 (
            .O(N__27383),
            .I(encoder0_position_7));
    InMux I__2971 (
            .O(N__27376),
            .I(N__27370));
    InMux I__2970 (
            .O(N__27375),
            .I(N__27370));
    LocalMux I__2969 (
            .O(N__27370),
            .I(data_out_frame_9_7));
    CascadeMux I__2968 (
            .O(N__27367),
            .I(N__27364));
    InMux I__2967 (
            .O(N__27364),
            .I(N__27361));
    LocalMux I__2966 (
            .O(N__27361),
            .I(\c0.n11_adj_3472 ));
    InMux I__2965 (
            .O(N__27358),
            .I(N__27355));
    LocalMux I__2964 (
            .O(N__27355),
            .I(\c0.n11_adj_3479 ));
    CascadeMux I__2963 (
            .O(N__27352),
            .I(\c0.n11_adj_3444_cascade_ ));
    CascadeMux I__2962 (
            .O(N__27349),
            .I(\c0.n21289_cascade_ ));
    InMux I__2961 (
            .O(N__27346),
            .I(N__27342));
    InMux I__2960 (
            .O(N__27345),
            .I(N__27339));
    LocalMux I__2959 (
            .O(N__27342),
            .I(N__27336));
    LocalMux I__2958 (
            .O(N__27339),
            .I(data_out_frame_6_1));
    Odrv4 I__2957 (
            .O(N__27336),
            .I(data_out_frame_6_1));
    InMux I__2956 (
            .O(N__27331),
            .I(N__27328));
    LocalMux I__2955 (
            .O(N__27328),
            .I(N__27323));
    CascadeMux I__2954 (
            .O(N__27327),
            .I(N__27320));
    InMux I__2953 (
            .O(N__27326),
            .I(N__27317));
    Span4Mux_v I__2952 (
            .O(N__27323),
            .I(N__27314));
    InMux I__2951 (
            .O(N__27320),
            .I(N__27311));
    LocalMux I__2950 (
            .O(N__27317),
            .I(encoder0_position_1));
    Odrv4 I__2949 (
            .O(N__27314),
            .I(encoder0_position_1));
    LocalMux I__2948 (
            .O(N__27311),
            .I(encoder0_position_1));
    InMux I__2947 (
            .O(N__27304),
            .I(N__27301));
    LocalMux I__2946 (
            .O(N__27301),
            .I(n2251));
    InMux I__2945 (
            .O(N__27298),
            .I(N__27294));
    CascadeMux I__2944 (
            .O(N__27297),
            .I(N__27290));
    LocalMux I__2943 (
            .O(N__27294),
            .I(N__27287));
    InMux I__2942 (
            .O(N__27293),
            .I(N__27284));
    InMux I__2941 (
            .O(N__27290),
            .I(N__27281));
    Odrv4 I__2940 (
            .O(N__27287),
            .I(encoder0_position_28));
    LocalMux I__2939 (
            .O(N__27284),
            .I(encoder0_position_28));
    LocalMux I__2938 (
            .O(N__27281),
            .I(encoder0_position_28));
    InMux I__2937 (
            .O(N__27274),
            .I(N__27270));
    CascadeMux I__2936 (
            .O(N__27273),
            .I(N__27266));
    LocalMux I__2935 (
            .O(N__27270),
            .I(N__27263));
    InMux I__2934 (
            .O(N__27269),
            .I(N__27260));
    InMux I__2933 (
            .O(N__27266),
            .I(N__27257));
    Odrv4 I__2932 (
            .O(N__27263),
            .I(encoder0_position_16));
    LocalMux I__2931 (
            .O(N__27260),
            .I(encoder0_position_16));
    LocalMux I__2930 (
            .O(N__27257),
            .I(encoder0_position_16));
    InMux I__2929 (
            .O(N__27250),
            .I(N__27246));
    CascadeMux I__2928 (
            .O(N__27249),
            .I(N__27242));
    LocalMux I__2927 (
            .O(N__27246),
            .I(N__27239));
    InMux I__2926 (
            .O(N__27245),
            .I(N__27236));
    InMux I__2925 (
            .O(N__27242),
            .I(N__27233));
    Odrv12 I__2924 (
            .O(N__27239),
            .I(encoder0_position_14));
    LocalMux I__2923 (
            .O(N__27236),
            .I(encoder0_position_14));
    LocalMux I__2922 (
            .O(N__27233),
            .I(encoder0_position_14));
    CascadeMux I__2921 (
            .O(N__27226),
            .I(N__27222));
    InMux I__2920 (
            .O(N__27225),
            .I(N__27219));
    InMux I__2919 (
            .O(N__27222),
            .I(N__27216));
    LocalMux I__2918 (
            .O(N__27219),
            .I(data_out_frame_8_6));
    LocalMux I__2917 (
            .O(N__27216),
            .I(data_out_frame_8_6));
    CascadeMux I__2916 (
            .O(N__27211),
            .I(N__27208));
    InMux I__2915 (
            .O(N__27208),
            .I(N__27204));
    InMux I__2914 (
            .O(N__27207),
            .I(N__27200));
    LocalMux I__2913 (
            .O(N__27204),
            .I(N__27197));
    InMux I__2912 (
            .O(N__27203),
            .I(N__27194));
    LocalMux I__2911 (
            .O(N__27200),
            .I(N__27189));
    Span4Mux_h I__2910 (
            .O(N__27197),
            .I(N__27189));
    LocalMux I__2909 (
            .O(N__27194),
            .I(encoder0_position_4));
    Odrv4 I__2908 (
            .O(N__27189),
            .I(encoder0_position_4));
    InMux I__2907 (
            .O(N__27184),
            .I(N__27181));
    LocalMux I__2906 (
            .O(N__27181),
            .I(\c0.n21632 ));
    InMux I__2905 (
            .O(N__27178),
            .I(N__27175));
    LocalMux I__2904 (
            .O(N__27175),
            .I(N__27172));
    Odrv4 I__2903 (
            .O(N__27172),
            .I(\c0.n21299 ));
    InMux I__2902 (
            .O(N__27169),
            .I(N__27165));
    InMux I__2901 (
            .O(N__27168),
            .I(N__27162));
    LocalMux I__2900 (
            .O(N__27165),
            .I(N__27159));
    LocalMux I__2899 (
            .O(N__27162),
            .I(data_out_frame_8_7));
    Odrv4 I__2898 (
            .O(N__27159),
            .I(data_out_frame_8_7));
    InMux I__2897 (
            .O(N__27154),
            .I(N__27150));
    CascadeMux I__2896 (
            .O(N__27153),
            .I(N__27146));
    LocalMux I__2895 (
            .O(N__27150),
            .I(N__27143));
    InMux I__2894 (
            .O(N__27149),
            .I(N__27140));
    InMux I__2893 (
            .O(N__27146),
            .I(N__27137));
    Odrv4 I__2892 (
            .O(N__27143),
            .I(encoder0_position_25));
    LocalMux I__2891 (
            .O(N__27140),
            .I(encoder0_position_25));
    LocalMux I__2890 (
            .O(N__27137),
            .I(encoder0_position_25));
    CascadeMux I__2889 (
            .O(N__27130),
            .I(N__27125));
    InMux I__2888 (
            .O(N__27129),
            .I(N__27122));
    InMux I__2887 (
            .O(N__27128),
            .I(N__27119));
    InMux I__2886 (
            .O(N__27125),
            .I(N__27116));
    LocalMux I__2885 (
            .O(N__27122),
            .I(encoder0_position_10));
    LocalMux I__2884 (
            .O(N__27119),
            .I(encoder0_position_10));
    LocalMux I__2883 (
            .O(N__27116),
            .I(encoder0_position_10));
    InMux I__2882 (
            .O(N__27109),
            .I(N__27104));
    CascadeMux I__2881 (
            .O(N__27108),
            .I(N__27101));
    InMux I__2880 (
            .O(N__27107),
            .I(N__27098));
    LocalMux I__2879 (
            .O(N__27104),
            .I(N__27095));
    InMux I__2878 (
            .O(N__27101),
            .I(N__27092));
    LocalMux I__2877 (
            .O(N__27098),
            .I(encoder0_position_20));
    Odrv4 I__2876 (
            .O(N__27095),
            .I(encoder0_position_20));
    LocalMux I__2875 (
            .O(N__27092),
            .I(encoder0_position_20));
    InMux I__2874 (
            .O(N__27085),
            .I(N__27082));
    LocalMux I__2873 (
            .O(N__27082),
            .I(N__27078));
    InMux I__2872 (
            .O(N__27081),
            .I(N__27075));
    Span4Mux_h I__2871 (
            .O(N__27078),
            .I(N__27072));
    LocalMux I__2870 (
            .O(N__27075),
            .I(data_out_frame_7_4));
    Odrv4 I__2869 (
            .O(N__27072),
            .I(data_out_frame_7_4));
    InMux I__2868 (
            .O(N__27067),
            .I(N__27064));
    LocalMux I__2867 (
            .O(N__27064),
            .I(n2253));
    InMux I__2866 (
            .O(N__27061),
            .I(N__27058));
    LocalMux I__2865 (
            .O(N__27058),
            .I(n2249));
    CascadeMux I__2864 (
            .O(N__27055),
            .I(N__27052));
    InMux I__2863 (
            .O(N__27052),
            .I(N__27048));
    CascadeMux I__2862 (
            .O(N__27051),
            .I(N__27044));
    LocalMux I__2861 (
            .O(N__27048),
            .I(N__27041));
    InMux I__2860 (
            .O(N__27047),
            .I(N__27038));
    InMux I__2859 (
            .O(N__27044),
            .I(N__27035));
    Odrv4 I__2858 (
            .O(N__27041),
            .I(encoder0_position_30));
    LocalMux I__2857 (
            .O(N__27038),
            .I(encoder0_position_30));
    LocalMux I__2856 (
            .O(N__27035),
            .I(encoder0_position_30));
    InMux I__2855 (
            .O(N__27028),
            .I(N__27025));
    LocalMux I__2854 (
            .O(N__27025),
            .I(n2267));
    InMux I__2853 (
            .O(N__27022),
            .I(N__27019));
    LocalMux I__2852 (
            .O(N__27019),
            .I(n2266));
    InMux I__2851 (
            .O(N__27016),
            .I(N__27013));
    LocalMux I__2850 (
            .O(N__27013),
            .I(n2265));
    InMux I__2849 (
            .O(N__27010),
            .I(N__27007));
    LocalMux I__2848 (
            .O(N__27007),
            .I(n2264));
    InMux I__2847 (
            .O(N__27004),
            .I(N__27000));
    CascadeMux I__2846 (
            .O(N__27003),
            .I(N__26997));
    LocalMux I__2845 (
            .O(N__27000),
            .I(N__26993));
    InMux I__2844 (
            .O(N__26997),
            .I(N__26990));
    InMux I__2843 (
            .O(N__26996),
            .I(N__26987));
    Span12Mux_v I__2842 (
            .O(N__26993),
            .I(N__26984));
    LocalMux I__2841 (
            .O(N__26990),
            .I(N__26981));
    LocalMux I__2840 (
            .O(N__26987),
            .I(encoder0_position_15));
    Odrv12 I__2839 (
            .O(N__26984),
            .I(encoder0_position_15));
    Odrv4 I__2838 (
            .O(N__26981),
            .I(encoder0_position_15));
    InMux I__2837 (
            .O(N__26974),
            .I(N__26971));
    LocalMux I__2836 (
            .O(N__26971),
            .I(n2263));
    InMux I__2835 (
            .O(N__26968),
            .I(N__26965));
    LocalMux I__2834 (
            .O(N__26965),
            .I(n2262));
    InMux I__2833 (
            .O(N__26962),
            .I(N__26959));
    LocalMux I__2832 (
            .O(N__26959),
            .I(N__26955));
    InMux I__2831 (
            .O(N__26958),
            .I(N__26952));
    Span4Mux_h I__2830 (
            .O(N__26955),
            .I(N__26949));
    LocalMux I__2829 (
            .O(N__26952),
            .I(data_out_frame_6_4));
    Odrv4 I__2828 (
            .O(N__26949),
            .I(data_out_frame_6_4));
    CascadeMux I__2827 (
            .O(N__26944),
            .I(\quad_counter1.n16_cascade_ ));
    CascadeMux I__2826 (
            .O(N__26941),
            .I(\quad_counter1.n24_adj_3578_cascade_ ));
    InMux I__2825 (
            .O(N__26938),
            .I(N__26932));
    InMux I__2824 (
            .O(N__26937),
            .I(N__26932));
    LocalMux I__2823 (
            .O(N__26932),
            .I(n11351));
    CascadeMux I__2822 (
            .O(N__26929),
            .I(N__26924));
    InMux I__2821 (
            .O(N__26928),
            .I(N__26919));
    InMux I__2820 (
            .O(N__26927),
            .I(N__26919));
    InMux I__2819 (
            .O(N__26924),
            .I(N__26916));
    LocalMux I__2818 (
            .O(N__26919),
            .I(N__26911));
    LocalMux I__2817 (
            .O(N__26916),
            .I(N__26911));
    Odrv4 I__2816 (
            .O(N__26911),
            .I(B_filtered));
    InMux I__2815 (
            .O(N__26908),
            .I(N__26905));
    LocalMux I__2814 (
            .O(N__26905),
            .I(N__26900));
    InMux I__2813 (
            .O(N__26904),
            .I(N__26895));
    InMux I__2812 (
            .O(N__26903),
            .I(N__26895));
    Odrv4 I__2811 (
            .O(N__26900),
            .I(\quad_counter0.B_delayed ));
    LocalMux I__2810 (
            .O(N__26895),
            .I(\quad_counter0.B_delayed ));
    InMux I__2809 (
            .O(N__26890),
            .I(N__26887));
    LocalMux I__2808 (
            .O(N__26887),
            .I(\quad_counter1.n6 ));
    InMux I__2807 (
            .O(N__26884),
            .I(N__26875));
    InMux I__2806 (
            .O(N__26883),
            .I(N__26875));
    InMux I__2805 (
            .O(N__26882),
            .I(N__26870));
    InMux I__2804 (
            .O(N__26881),
            .I(N__26870));
    InMux I__2803 (
            .O(N__26880),
            .I(N__26867));
    LocalMux I__2802 (
            .O(N__26875),
            .I(N__26864));
    LocalMux I__2801 (
            .O(N__26870),
            .I(N__26861));
    LocalMux I__2800 (
            .O(N__26867),
            .I(A_filtered));
    Odrv4 I__2799 (
            .O(N__26864),
            .I(A_filtered));
    Odrv4 I__2798 (
            .O(N__26861),
            .I(A_filtered));
    InMux I__2797 (
            .O(N__26854),
            .I(N__26851));
    LocalMux I__2796 (
            .O(N__26851),
            .I(\quad_counter0.A_delayed ));
    InMux I__2795 (
            .O(N__26848),
            .I(N__26845));
    LocalMux I__2794 (
            .O(N__26845),
            .I(\quad_counter1.n22 ));
    InMux I__2793 (
            .O(N__26842),
            .I(N__26839));
    LocalMux I__2792 (
            .O(N__26839),
            .I(n2269));
    InMux I__2791 (
            .O(N__26836),
            .I(N__26833));
    LocalMux I__2790 (
            .O(N__26833),
            .I(n2268));
    CascadeMux I__2789 (
            .O(N__26830),
            .I(n11343_cascade_));
    CascadeMux I__2788 (
            .O(N__26827),
            .I(n12417_cascade_));
    InMux I__2787 (
            .O(N__26824),
            .I(N__26821));
    LocalMux I__2786 (
            .O(N__26821),
            .I(\quad_counter1.n28_adj_3574 ));
    InMux I__2785 (
            .O(N__26818),
            .I(N__26810));
    InMux I__2784 (
            .O(N__26817),
            .I(N__26810));
    InMux I__2783 (
            .O(N__26816),
            .I(N__26805));
    InMux I__2782 (
            .O(N__26815),
            .I(N__26805));
    LocalMux I__2781 (
            .O(N__26810),
            .I(N__26800));
    LocalMux I__2780 (
            .O(N__26805),
            .I(N__26800));
    Span4Mux_v I__2779 (
            .O(N__26800),
            .I(N__26797));
    Sp12to4 I__2778 (
            .O(N__26797),
            .I(N__26794));
    Odrv12 I__2777 (
            .O(N__26794),
            .I(PIN_13_c));
    CascadeMux I__2776 (
            .O(N__26791),
            .I(N__26788));
    InMux I__2775 (
            .O(N__26788),
            .I(N__26785));
    LocalMux I__2774 (
            .O(N__26785),
            .I(n11343));
    InMux I__2773 (
            .O(N__26782),
            .I(N__26775));
    InMux I__2772 (
            .O(N__26781),
            .I(N__26775));
    InMux I__2771 (
            .O(N__26780),
            .I(N__26772));
    LocalMux I__2770 (
            .O(N__26775),
            .I(quadB_delayed_adj_3585));
    LocalMux I__2769 (
            .O(N__26772),
            .I(quadB_delayed_adj_3585));
    InMux I__2768 (
            .O(N__26767),
            .I(N__26764));
    LocalMux I__2767 (
            .O(N__26764),
            .I(\quad_counter1.n26_adj_3575 ));
    InMux I__2766 (
            .O(N__26761),
            .I(N__26758));
    LocalMux I__2765 (
            .O(N__26758),
            .I(\quad_counter1.n27_adj_3576 ));
    SRMux I__2764 (
            .O(N__26755),
            .I(N__26752));
    LocalMux I__2763 (
            .O(N__26752),
            .I(N__26749));
    Odrv4 I__2762 (
            .O(N__26749),
            .I(\c0.n18671 ));
    SRMux I__2761 (
            .O(N__26746),
            .I(N__26743));
    LocalMux I__2760 (
            .O(N__26743),
            .I(N__26740));
    Span4Mux_h I__2759 (
            .O(N__26740),
            .I(N__26737));
    Odrv4 I__2758 (
            .O(N__26737),
            .I(\c0.n18617 ));
    CascadeMux I__2757 (
            .O(N__26734),
            .I(\quad_counter1.n25_adj_3577_cascade_ ));
    CascadeMux I__2756 (
            .O(N__26731),
            .I(N__26727));
    InMux I__2755 (
            .O(N__26730),
            .I(N__26724));
    InMux I__2754 (
            .O(N__26727),
            .I(N__26721));
    LocalMux I__2753 (
            .O(N__26724),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__2752 (
            .O(N__26721),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__2751 (
            .O(N__26716),
            .I(\c0.tx.n17274 ));
    InMux I__2750 (
            .O(N__26713),
            .I(N__26709));
    InMux I__2749 (
            .O(N__26712),
            .I(N__26706));
    LocalMux I__2748 (
            .O(N__26709),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__2747 (
            .O(N__26706),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__2746 (
            .O(N__26701),
            .I(\c0.tx.n17275 ));
    InMux I__2745 (
            .O(N__26698),
            .I(N__26694));
    InMux I__2744 (
            .O(N__26697),
            .I(N__26691));
    LocalMux I__2743 (
            .O(N__26694),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__2742 (
            .O(N__26691),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__2741 (
            .O(N__26686),
            .I(\c0.tx.n17276 ));
    InMux I__2740 (
            .O(N__26683),
            .I(N__26679));
    InMux I__2739 (
            .O(N__26682),
            .I(N__26676));
    LocalMux I__2738 (
            .O(N__26679),
            .I(\c0.tx.r_Clock_Count_4 ));
    LocalMux I__2737 (
            .O(N__26676),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__2736 (
            .O(N__26671),
            .I(\c0.tx.n17277 ));
    InMux I__2735 (
            .O(N__26668),
            .I(N__26664));
    InMux I__2734 (
            .O(N__26667),
            .I(N__26661));
    LocalMux I__2733 (
            .O(N__26664),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__2732 (
            .O(N__26661),
            .I(\c0.tx.r_Clock_Count_5 ));
    InMux I__2731 (
            .O(N__26656),
            .I(\c0.tx.n17278 ));
    InMux I__2730 (
            .O(N__26653),
            .I(N__26649));
    InMux I__2729 (
            .O(N__26652),
            .I(N__26646));
    LocalMux I__2728 (
            .O(N__26649),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__2727 (
            .O(N__26646),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__2726 (
            .O(N__26641),
            .I(\c0.tx.n17279 ));
    InMux I__2725 (
            .O(N__26638),
            .I(N__26634));
    InMux I__2724 (
            .O(N__26637),
            .I(N__26631));
    LocalMux I__2723 (
            .O(N__26634),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__2722 (
            .O(N__26631),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__2721 (
            .O(N__26626),
            .I(\c0.tx.n17280 ));
    InMux I__2720 (
            .O(N__26623),
            .I(bfn_10_19_0_));
    CascadeMux I__2719 (
            .O(N__26620),
            .I(N__26617));
    InMux I__2718 (
            .O(N__26617),
            .I(N__26596));
    InMux I__2717 (
            .O(N__26616),
            .I(N__26596));
    InMux I__2716 (
            .O(N__26615),
            .I(N__26596));
    InMux I__2715 (
            .O(N__26614),
            .I(N__26591));
    InMux I__2714 (
            .O(N__26613),
            .I(N__26588));
    InMux I__2713 (
            .O(N__26612),
            .I(N__26581));
    InMux I__2712 (
            .O(N__26611),
            .I(N__26581));
    InMux I__2711 (
            .O(N__26610),
            .I(N__26581));
    InMux I__2710 (
            .O(N__26609),
            .I(N__26578));
    InMux I__2709 (
            .O(N__26608),
            .I(N__26565));
    InMux I__2708 (
            .O(N__26607),
            .I(N__26565));
    InMux I__2707 (
            .O(N__26606),
            .I(N__26565));
    InMux I__2706 (
            .O(N__26605),
            .I(N__26565));
    InMux I__2705 (
            .O(N__26604),
            .I(N__26565));
    InMux I__2704 (
            .O(N__26603),
            .I(N__26565));
    LocalMux I__2703 (
            .O(N__26596),
            .I(N__26562));
    InMux I__2702 (
            .O(N__26595),
            .I(N__26559));
    InMux I__2701 (
            .O(N__26594),
            .I(N__26556));
    LocalMux I__2700 (
            .O(N__26591),
            .I(N__26551));
    LocalMux I__2699 (
            .O(N__26588),
            .I(N__26551));
    LocalMux I__2698 (
            .O(N__26581),
            .I(N__26548));
    LocalMux I__2697 (
            .O(N__26578),
            .I(N__26543));
    LocalMux I__2696 (
            .O(N__26565),
            .I(N__26543));
    Span4Mux_h I__2695 (
            .O(N__26562),
            .I(N__26536));
    LocalMux I__2694 (
            .O(N__26559),
            .I(N__26536));
    LocalMux I__2693 (
            .O(N__26556),
            .I(N__26533));
    Sp12to4 I__2692 (
            .O(N__26551),
            .I(N__26530));
    Span4Mux_v I__2691 (
            .O(N__26548),
            .I(N__26527));
    Sp12to4 I__2690 (
            .O(N__26543),
            .I(N__26524));
    InMux I__2689 (
            .O(N__26542),
            .I(N__26519));
    InMux I__2688 (
            .O(N__26541),
            .I(N__26519));
    Span4Mux_h I__2687 (
            .O(N__26536),
            .I(N__26516));
    Span4Mux_v I__2686 (
            .O(N__26533),
            .I(N__26513));
    Span12Mux_v I__2685 (
            .O(N__26530),
            .I(N__26504));
    Sp12to4 I__2684 (
            .O(N__26527),
            .I(N__26504));
    Span12Mux_v I__2683 (
            .O(N__26524),
            .I(N__26504));
    LocalMux I__2682 (
            .O(N__26519),
            .I(N__26504));
    Span4Mux_v I__2681 (
            .O(N__26516),
            .I(N__26499));
    Span4Mux_h I__2680 (
            .O(N__26513),
            .I(N__26499));
    Odrv12 I__2679 (
            .O(N__26504),
            .I(PIN_8_c));
    Odrv4 I__2678 (
            .O(N__26499),
            .I(PIN_8_c));
    CascadeMux I__2677 (
            .O(N__26494),
            .I(N__26479));
    InMux I__2676 (
            .O(N__26493),
            .I(N__26475));
    InMux I__2675 (
            .O(N__26492),
            .I(N__26466));
    InMux I__2674 (
            .O(N__26491),
            .I(N__26466));
    InMux I__2673 (
            .O(N__26490),
            .I(N__26453));
    InMux I__2672 (
            .O(N__26489),
            .I(N__26453));
    InMux I__2671 (
            .O(N__26488),
            .I(N__26453));
    InMux I__2670 (
            .O(N__26487),
            .I(N__26453));
    InMux I__2669 (
            .O(N__26486),
            .I(N__26453));
    InMux I__2668 (
            .O(N__26485),
            .I(N__26453));
    InMux I__2667 (
            .O(N__26484),
            .I(N__26446));
    InMux I__2666 (
            .O(N__26483),
            .I(N__26446));
    InMux I__2665 (
            .O(N__26482),
            .I(N__26446));
    InMux I__2664 (
            .O(N__26479),
            .I(N__26443));
    InMux I__2663 (
            .O(N__26478),
            .I(N__26440));
    LocalMux I__2662 (
            .O(N__26475),
            .I(N__26437));
    InMux I__2661 (
            .O(N__26474),
            .I(N__26430));
    InMux I__2660 (
            .O(N__26473),
            .I(N__26430));
    InMux I__2659 (
            .O(N__26472),
            .I(N__26430));
    InMux I__2658 (
            .O(N__26471),
            .I(N__26427));
    LocalMux I__2657 (
            .O(N__26466),
            .I(N__26424));
    LocalMux I__2656 (
            .O(N__26453),
            .I(N__26419));
    LocalMux I__2655 (
            .O(N__26446),
            .I(N__26419));
    LocalMux I__2654 (
            .O(N__26443),
            .I(N__26416));
    LocalMux I__2653 (
            .O(N__26440),
            .I(N__26411));
    Span4Mux_h I__2652 (
            .O(N__26437),
            .I(N__26411));
    LocalMux I__2651 (
            .O(N__26430),
            .I(N__26408));
    LocalMux I__2650 (
            .O(N__26427),
            .I(N__26405));
    Span4Mux_v I__2649 (
            .O(N__26424),
            .I(N__26400));
    Span4Mux_v I__2648 (
            .O(N__26419),
            .I(N__26400));
    Span12Mux_h I__2647 (
            .O(N__26416),
            .I(N__26397));
    Span4Mux_v I__2646 (
            .O(N__26411),
            .I(N__26392));
    Span4Mux_h I__2645 (
            .O(N__26408),
            .I(N__26392));
    Odrv4 I__2644 (
            .O(N__26405),
            .I(quadB_delayed));
    Odrv4 I__2643 (
            .O(N__26400),
            .I(quadB_delayed));
    Odrv12 I__2642 (
            .O(N__26397),
            .I(quadB_delayed));
    Odrv4 I__2641 (
            .O(N__26392),
            .I(quadB_delayed));
    InMux I__2640 (
            .O(N__26383),
            .I(N__26380));
    LocalMux I__2639 (
            .O(N__26380),
            .I(N__26377));
    Odrv4 I__2638 (
            .O(N__26377),
            .I(\quad_counter0.n13187 ));
    InMux I__2637 (
            .O(N__26374),
            .I(N__26370));
    InMux I__2636 (
            .O(N__26373),
            .I(N__26367));
    LocalMux I__2635 (
            .O(N__26370),
            .I(N__26361));
    LocalMux I__2634 (
            .O(N__26367),
            .I(N__26361));
    CascadeMux I__2633 (
            .O(N__26366),
            .I(N__26358));
    Span4Mux_h I__2632 (
            .O(N__26361),
            .I(N__26355));
    InMux I__2631 (
            .O(N__26358),
            .I(N__26352));
    Odrv4 I__2630 (
            .O(N__26355),
            .I(\quad_counter0.b_delay_counter_2 ));
    LocalMux I__2629 (
            .O(N__26352),
            .I(\quad_counter0.b_delay_counter_2 ));
    CascadeMux I__2628 (
            .O(N__26347),
            .I(\c0.n21331_cascade_ ));
    CascadeMux I__2627 (
            .O(N__26344),
            .I(\c0.n17354_cascade_ ));
    InMux I__2626 (
            .O(N__26341),
            .I(N__26338));
    LocalMux I__2625 (
            .O(N__26338),
            .I(\c0.n21521 ));
    CascadeMux I__2624 (
            .O(N__26335),
            .I(\c0.tx.n6_cascade_ ));
    CascadeMux I__2623 (
            .O(N__26332),
            .I(\c0.n15938_cascade_ ));
    InMux I__2622 (
            .O(N__26329),
            .I(N__26326));
    LocalMux I__2621 (
            .O(N__26326),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__2620 (
            .O(N__26323),
            .I(bfn_10_18_0_));
    InMux I__2619 (
            .O(N__26320),
            .I(N__26317));
    LocalMux I__2618 (
            .O(N__26317),
            .I(\quad_counter0.n13269 ));
    InMux I__2617 (
            .O(N__26314),
            .I(N__26309));
    InMux I__2616 (
            .O(N__26313),
            .I(N__26306));
    InMux I__2615 (
            .O(N__26312),
            .I(N__26303));
    LocalMux I__2614 (
            .O(N__26309),
            .I(N__26300));
    LocalMux I__2613 (
            .O(N__26306),
            .I(N__26295));
    LocalMux I__2612 (
            .O(N__26303),
            .I(N__26295));
    Odrv12 I__2611 (
            .O(N__26300),
            .I(\quad_counter0.b_delay_counter_15 ));
    Odrv4 I__2610 (
            .O(N__26295),
            .I(\quad_counter0.b_delay_counter_15 ));
    InMux I__2609 (
            .O(N__26290),
            .I(N__26287));
    LocalMux I__2608 (
            .O(N__26287),
            .I(N__26284));
    Odrv4 I__2607 (
            .O(N__26284),
            .I(\quad_counter0.n26_adj_2991 ));
    InMux I__2606 (
            .O(N__26281),
            .I(N__26278));
    LocalMux I__2605 (
            .O(N__26278),
            .I(N__26275));
    Odrv4 I__2604 (
            .O(N__26275),
            .I(\quad_counter0.n27_adj_2992 ));
    CascadeMux I__2603 (
            .O(N__26272),
            .I(N__26269));
    InMux I__2602 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__2601 (
            .O(N__26266),
            .I(\quad_counter0.n28_adj_2990 ));
    InMux I__2600 (
            .O(N__26263),
            .I(N__26260));
    LocalMux I__2599 (
            .O(N__26260),
            .I(\quad_counter0.n25_adj_2993 ));
    InMux I__2598 (
            .O(N__26257),
            .I(N__26254));
    LocalMux I__2597 (
            .O(N__26254),
            .I(N__26251));
    Span12Mux_v I__2596 (
            .O(N__26251),
            .I(N__26248));
    Odrv12 I__2595 (
            .O(N__26248),
            .I(n11347));
    CascadeMux I__2594 (
            .O(N__26245),
            .I(n11347_cascade_));
    CascadeMux I__2593 (
            .O(N__26242),
            .I(N__26224));
    CascadeMux I__2592 (
            .O(N__26241),
            .I(N__26221));
    CascadeMux I__2591 (
            .O(N__26240),
            .I(N__26218));
    CascadeMux I__2590 (
            .O(N__26239),
            .I(N__26215));
    CascadeMux I__2589 (
            .O(N__26238),
            .I(N__26212));
    CascadeMux I__2588 (
            .O(N__26237),
            .I(N__26209));
    CascadeMux I__2587 (
            .O(N__26236),
            .I(N__26206));
    CascadeMux I__2586 (
            .O(N__26235),
            .I(N__26203));
    CascadeMux I__2585 (
            .O(N__26234),
            .I(N__26200));
    CascadeMux I__2584 (
            .O(N__26233),
            .I(N__26197));
    CascadeMux I__2583 (
            .O(N__26232),
            .I(N__26194));
    CascadeMux I__2582 (
            .O(N__26231),
            .I(N__26191));
    CascadeMux I__2581 (
            .O(N__26230),
            .I(N__26188));
    CascadeMux I__2580 (
            .O(N__26229),
            .I(N__26185));
    CascadeMux I__2579 (
            .O(N__26228),
            .I(N__26182));
    CascadeMux I__2578 (
            .O(N__26227),
            .I(N__26179));
    InMux I__2577 (
            .O(N__26224),
            .I(N__26170));
    InMux I__2576 (
            .O(N__26221),
            .I(N__26170));
    InMux I__2575 (
            .O(N__26218),
            .I(N__26170));
    InMux I__2574 (
            .O(N__26215),
            .I(N__26170));
    InMux I__2573 (
            .O(N__26212),
            .I(N__26161));
    InMux I__2572 (
            .O(N__26209),
            .I(N__26161));
    InMux I__2571 (
            .O(N__26206),
            .I(N__26161));
    InMux I__2570 (
            .O(N__26203),
            .I(N__26161));
    InMux I__2569 (
            .O(N__26200),
            .I(N__26152));
    InMux I__2568 (
            .O(N__26197),
            .I(N__26152));
    InMux I__2567 (
            .O(N__26194),
            .I(N__26152));
    InMux I__2566 (
            .O(N__26191),
            .I(N__26152));
    InMux I__2565 (
            .O(N__26188),
            .I(N__26143));
    InMux I__2564 (
            .O(N__26185),
            .I(N__26143));
    InMux I__2563 (
            .O(N__26182),
            .I(N__26143));
    InMux I__2562 (
            .O(N__26179),
            .I(N__26143));
    LocalMux I__2561 (
            .O(N__26170),
            .I(\quad_counter0.n21603 ));
    LocalMux I__2560 (
            .O(N__26161),
            .I(\quad_counter0.n21603 ));
    LocalMux I__2559 (
            .O(N__26152),
            .I(\quad_counter0.n21603 ));
    LocalMux I__2558 (
            .O(N__26143),
            .I(\quad_counter0.n21603 ));
    InMux I__2557 (
            .O(N__26134),
            .I(N__26128));
    InMux I__2556 (
            .O(N__26133),
            .I(N__26128));
    LocalMux I__2555 (
            .O(N__26128),
            .I(data_out_frame_10_6));
    InMux I__2554 (
            .O(N__26125),
            .I(N__26122));
    LocalMux I__2553 (
            .O(N__26122),
            .I(\c0.n21629 ));
    InMux I__2552 (
            .O(N__26119),
            .I(N__26116));
    LocalMux I__2551 (
            .O(N__26116),
            .I(N__26113));
    Span4Mux_v I__2550 (
            .O(N__26113),
            .I(N__26110));
    Odrv4 I__2549 (
            .O(N__26110),
            .I(n2275));
    InMux I__2548 (
            .O(N__26107),
            .I(N__26104));
    LocalMux I__2547 (
            .O(N__26104),
            .I(N__26101));
    Odrv12 I__2546 (
            .O(N__26101),
            .I(n2272));
    InMux I__2545 (
            .O(N__26098),
            .I(N__26095));
    LocalMux I__2544 (
            .O(N__26095),
            .I(N__26092));
    Odrv12 I__2543 (
            .O(N__26092),
            .I(n2274));
    InMux I__2542 (
            .O(N__26089),
            .I(N__26086));
    LocalMux I__2541 (
            .O(N__26086),
            .I(n2248));
    InMux I__2540 (
            .O(N__26083),
            .I(N__26080));
    LocalMux I__2539 (
            .O(N__26080),
            .I(N__26077));
    Odrv4 I__2538 (
            .O(N__26077),
            .I(\c0.n5_adj_3471 ));
    CascadeMux I__2537 (
            .O(N__26074),
            .I(N__26070));
    CascadeMux I__2536 (
            .O(N__26073),
            .I(N__26066));
    InMux I__2535 (
            .O(N__26070),
            .I(N__26063));
    InMux I__2534 (
            .O(N__26069),
            .I(N__26060));
    InMux I__2533 (
            .O(N__26066),
            .I(N__26057));
    LocalMux I__2532 (
            .O(N__26063),
            .I(N__26054));
    LocalMux I__2531 (
            .O(N__26060),
            .I(encoder0_position_5));
    LocalMux I__2530 (
            .O(N__26057),
            .I(encoder0_position_5));
    Odrv12 I__2529 (
            .O(N__26054),
            .I(encoder0_position_5));
    InMux I__2528 (
            .O(N__26047),
            .I(N__26041));
    InMux I__2527 (
            .O(N__26046),
            .I(N__26041));
    LocalMux I__2526 (
            .O(N__26041),
            .I(data_out_frame_9_6));
    InMux I__2525 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__2524 (
            .O(N__26035),
            .I(\quad_counter0.n13254 ));
    InMux I__2523 (
            .O(N__26032),
            .I(N__26027));
    InMux I__2522 (
            .O(N__26031),
            .I(N__26024));
    InMux I__2521 (
            .O(N__26030),
            .I(N__26021));
    LocalMux I__2520 (
            .O(N__26027),
            .I(N__26018));
    LocalMux I__2519 (
            .O(N__26024),
            .I(\quad_counter0.b_delay_counter_10 ));
    LocalMux I__2518 (
            .O(N__26021),
            .I(\quad_counter0.b_delay_counter_10 ));
    Odrv4 I__2517 (
            .O(N__26018),
            .I(\quad_counter0.b_delay_counter_10 ));
    InMux I__2516 (
            .O(N__26011),
            .I(N__26008));
    LocalMux I__2515 (
            .O(N__26008),
            .I(n2255));
    InMux I__2514 (
            .O(N__26005),
            .I(\quad_counter0.n17306 ));
    InMux I__2513 (
            .O(N__26002),
            .I(N__25999));
    LocalMux I__2512 (
            .O(N__25999),
            .I(n2254));
    InMux I__2511 (
            .O(N__25996),
            .I(\quad_counter0.n17307 ));
    InMux I__2510 (
            .O(N__25993),
            .I(\quad_counter0.n17308 ));
    InMux I__2509 (
            .O(N__25990),
            .I(\quad_counter0.n17309 ));
    InMux I__2508 (
            .O(N__25987),
            .I(\quad_counter0.n17310 ));
    InMux I__2507 (
            .O(N__25984),
            .I(\quad_counter0.n17311 ));
    InMux I__2506 (
            .O(N__25981),
            .I(\quad_counter0.n17312 ));
    InMux I__2505 (
            .O(N__25978),
            .I(N__25974));
    CascadeMux I__2504 (
            .O(N__25977),
            .I(N__25960));
    LocalMux I__2503 (
            .O(N__25974),
            .I(N__25951));
    InMux I__2502 (
            .O(N__25973),
            .I(N__25942));
    InMux I__2501 (
            .O(N__25972),
            .I(N__25942));
    InMux I__2500 (
            .O(N__25971),
            .I(N__25942));
    InMux I__2499 (
            .O(N__25970),
            .I(N__25942));
    InMux I__2498 (
            .O(N__25969),
            .I(N__25933));
    InMux I__2497 (
            .O(N__25968),
            .I(N__25933));
    InMux I__2496 (
            .O(N__25967),
            .I(N__25933));
    InMux I__2495 (
            .O(N__25966),
            .I(N__25933));
    InMux I__2494 (
            .O(N__25965),
            .I(N__25922));
    InMux I__2493 (
            .O(N__25964),
            .I(N__25922));
    InMux I__2492 (
            .O(N__25963),
            .I(N__25922));
    InMux I__2491 (
            .O(N__25960),
            .I(N__25922));
    InMux I__2490 (
            .O(N__25959),
            .I(N__25922));
    InMux I__2489 (
            .O(N__25958),
            .I(N__25915));
    InMux I__2488 (
            .O(N__25957),
            .I(N__25915));
    InMux I__2487 (
            .O(N__25956),
            .I(N__25915));
    CascadeMux I__2486 (
            .O(N__25955),
            .I(N__25902));
    CascadeMux I__2485 (
            .O(N__25954),
            .I(N__25897));
    Span4Mux_v I__2484 (
            .O(N__25951),
            .I(N__25884));
    LocalMux I__2483 (
            .O(N__25942),
            .I(N__25884));
    LocalMux I__2482 (
            .O(N__25933),
            .I(N__25884));
    LocalMux I__2481 (
            .O(N__25922),
            .I(N__25884));
    LocalMux I__2480 (
            .O(N__25915),
            .I(N__25884));
    InMux I__2479 (
            .O(N__25914),
            .I(N__25875));
    InMux I__2478 (
            .O(N__25913),
            .I(N__25875));
    InMux I__2477 (
            .O(N__25912),
            .I(N__25875));
    InMux I__2476 (
            .O(N__25911),
            .I(N__25875));
    InMux I__2475 (
            .O(N__25910),
            .I(N__25866));
    InMux I__2474 (
            .O(N__25909),
            .I(N__25866));
    InMux I__2473 (
            .O(N__25908),
            .I(N__25866));
    InMux I__2472 (
            .O(N__25907),
            .I(N__25866));
    InMux I__2471 (
            .O(N__25906),
            .I(N__25859));
    InMux I__2470 (
            .O(N__25905),
            .I(N__25859));
    InMux I__2469 (
            .O(N__25902),
            .I(N__25859));
    InMux I__2468 (
            .O(N__25901),
            .I(N__25848));
    InMux I__2467 (
            .O(N__25900),
            .I(N__25848));
    InMux I__2466 (
            .O(N__25897),
            .I(N__25848));
    InMux I__2465 (
            .O(N__25896),
            .I(N__25848));
    InMux I__2464 (
            .O(N__25895),
            .I(N__25848));
    Odrv4 I__2463 (
            .O(N__25884),
            .I(\quad_counter0.n2228 ));
    LocalMux I__2462 (
            .O(N__25875),
            .I(\quad_counter0.n2228 ));
    LocalMux I__2461 (
            .O(N__25866),
            .I(\quad_counter0.n2228 ));
    LocalMux I__2460 (
            .O(N__25859),
            .I(\quad_counter0.n2228 ));
    LocalMux I__2459 (
            .O(N__25848),
            .I(\quad_counter0.n2228 ));
    InMux I__2458 (
            .O(N__25837),
            .I(bfn_10_13_0_));
    InMux I__2457 (
            .O(N__25834),
            .I(\quad_counter0.n17298 ));
    InMux I__2456 (
            .O(N__25831),
            .I(\quad_counter0.n17299 ));
    InMux I__2455 (
            .O(N__25828),
            .I(N__25825));
    LocalMux I__2454 (
            .O(N__25825),
            .I(n2261));
    InMux I__2453 (
            .O(N__25822),
            .I(\quad_counter0.n17300 ));
    InMux I__2452 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__2451 (
            .O(N__25816),
            .I(n2260));
    InMux I__2450 (
            .O(N__25813),
            .I(\quad_counter0.n17301 ));
    InMux I__2449 (
            .O(N__25810),
            .I(N__25807));
    LocalMux I__2448 (
            .O(N__25807),
            .I(n2259));
    InMux I__2447 (
            .O(N__25804),
            .I(\quad_counter0.n17302 ));
    InMux I__2446 (
            .O(N__25801),
            .I(N__25798));
    LocalMux I__2445 (
            .O(N__25798),
            .I(n2258));
    InMux I__2444 (
            .O(N__25795),
            .I(\quad_counter0.n17303 ));
    CascadeMux I__2443 (
            .O(N__25792),
            .I(N__25787));
    InMux I__2442 (
            .O(N__25791),
            .I(N__25784));
    InMux I__2441 (
            .O(N__25790),
            .I(N__25781));
    InMux I__2440 (
            .O(N__25787),
            .I(N__25778));
    LocalMux I__2439 (
            .O(N__25784),
            .I(encoder0_position_22));
    LocalMux I__2438 (
            .O(N__25781),
            .I(encoder0_position_22));
    LocalMux I__2437 (
            .O(N__25778),
            .I(encoder0_position_22));
    InMux I__2436 (
            .O(N__25771),
            .I(N__25768));
    LocalMux I__2435 (
            .O(N__25768),
            .I(n2257));
    InMux I__2434 (
            .O(N__25765),
            .I(\quad_counter0.n17304 ));
    InMux I__2433 (
            .O(N__25762),
            .I(N__25759));
    LocalMux I__2432 (
            .O(N__25759),
            .I(n2256));
    InMux I__2431 (
            .O(N__25756),
            .I(bfn_10_12_0_));
    InMux I__2430 (
            .O(N__25753),
            .I(bfn_10_10_0_));
    InMux I__2429 (
            .O(N__25750),
            .I(\quad_counter0.n17290 ));
    InMux I__2428 (
            .O(N__25747),
            .I(\quad_counter0.n17291 ));
    InMux I__2427 (
            .O(N__25744),
            .I(\quad_counter0.n17292 ));
    InMux I__2426 (
            .O(N__25741),
            .I(\quad_counter0.n17293 ));
    InMux I__2425 (
            .O(N__25738),
            .I(\quad_counter0.n17294 ));
    InMux I__2424 (
            .O(N__25735),
            .I(\quad_counter0.n17295 ));
    InMux I__2423 (
            .O(N__25732),
            .I(\quad_counter0.n17296 ));
    InMux I__2422 (
            .O(N__25729),
            .I(bfn_10_11_0_));
    InMux I__2421 (
            .O(N__25726),
            .I(N__25723));
    LocalMux I__2420 (
            .O(N__25723),
            .I(\quad_counter0.count_direction ));
    InMux I__2419 (
            .O(N__25720),
            .I(N__25717));
    LocalMux I__2418 (
            .O(N__25717),
            .I(N__25714));
    Odrv12 I__2417 (
            .O(N__25714),
            .I(n2279));
    InMux I__2416 (
            .O(N__25711),
            .I(\quad_counter0.n17282 ));
    InMux I__2415 (
            .O(N__25708),
            .I(N__25705));
    LocalMux I__2414 (
            .O(N__25705),
            .I(n2278));
    InMux I__2413 (
            .O(N__25702),
            .I(\quad_counter0.n17283 ));
    InMux I__2412 (
            .O(N__25699),
            .I(N__25694));
    InMux I__2411 (
            .O(N__25698),
            .I(N__25691));
    InMux I__2410 (
            .O(N__25697),
            .I(N__25688));
    LocalMux I__2409 (
            .O(N__25694),
            .I(encoder0_position_2));
    LocalMux I__2408 (
            .O(N__25691),
            .I(encoder0_position_2));
    LocalMux I__2407 (
            .O(N__25688),
            .I(encoder0_position_2));
    InMux I__2406 (
            .O(N__25681),
            .I(N__25678));
    LocalMux I__2405 (
            .O(N__25678),
            .I(n2277));
    InMux I__2404 (
            .O(N__25675),
            .I(\quad_counter0.n17284 ));
    InMux I__2403 (
            .O(N__25672),
            .I(N__25668));
    CascadeMux I__2402 (
            .O(N__25671),
            .I(N__25665));
    LocalMux I__2401 (
            .O(N__25668),
            .I(N__25662));
    InMux I__2400 (
            .O(N__25665),
            .I(N__25658));
    Span4Mux_v I__2399 (
            .O(N__25662),
            .I(N__25655));
    InMux I__2398 (
            .O(N__25661),
            .I(N__25652));
    LocalMux I__2397 (
            .O(N__25658),
            .I(N__25649));
    Odrv4 I__2396 (
            .O(N__25655),
            .I(encoder0_position_3));
    LocalMux I__2395 (
            .O(N__25652),
            .I(encoder0_position_3));
    Odrv4 I__2394 (
            .O(N__25649),
            .I(encoder0_position_3));
    InMux I__2393 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__2392 (
            .O(N__25639),
            .I(n2276));
    InMux I__2391 (
            .O(N__25636),
            .I(\quad_counter0.n17285 ));
    InMux I__2390 (
            .O(N__25633),
            .I(\quad_counter0.n17286 ));
    InMux I__2389 (
            .O(N__25630),
            .I(\quad_counter0.n17287 ));
    InMux I__2388 (
            .O(N__25627),
            .I(\quad_counter0.n17288 ));
    CEMux I__2387 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__2386 (
            .O(N__25621),
            .I(N__25618));
    Span4Mux_v I__2385 (
            .O(N__25618),
            .I(N__25613));
    CEMux I__2384 (
            .O(N__25617),
            .I(N__25610));
    InMux I__2383 (
            .O(N__25616),
            .I(N__25607));
    Odrv4 I__2382 (
            .O(N__25613),
            .I(n12447));
    LocalMux I__2381 (
            .O(N__25610),
            .I(n12447));
    LocalMux I__2380 (
            .O(N__25607),
            .I(n12447));
    CascadeMux I__2379 (
            .O(N__25600),
            .I(N__25595));
    InMux I__2378 (
            .O(N__25599),
            .I(N__25585));
    InMux I__2377 (
            .O(N__25598),
            .I(N__25585));
    InMux I__2376 (
            .O(N__25595),
            .I(N__25585));
    InMux I__2375 (
            .O(N__25594),
            .I(N__25585));
    LocalMux I__2374 (
            .O(N__25585),
            .I(N__25582));
    Span4Mux_v I__2373 (
            .O(N__25582),
            .I(N__25579));
    Sp12to4 I__2372 (
            .O(N__25579),
            .I(N__25576));
    Span12Mux_h I__2371 (
            .O(N__25576),
            .I(N__25573));
    Span12Mux_v I__2370 (
            .O(N__25573),
            .I(N__25570));
    Odrv12 I__2369 (
            .O(N__25570),
            .I(PIN_7_c));
    InMux I__2368 (
            .O(N__25567),
            .I(N__25558));
    InMux I__2367 (
            .O(N__25566),
            .I(N__25558));
    InMux I__2366 (
            .O(N__25565),
            .I(N__25558));
    LocalMux I__2365 (
            .O(N__25558),
            .I(quadA_delayed));
    InMux I__2364 (
            .O(N__25555),
            .I(N__25551));
    InMux I__2363 (
            .O(N__25554),
            .I(N__25548));
    LocalMux I__2362 (
            .O(N__25551),
            .I(\quad_counter0.a_delay_counter_15 ));
    LocalMux I__2361 (
            .O(N__25548),
            .I(\quad_counter0.a_delay_counter_15 ));
    InMux I__2360 (
            .O(N__25543),
            .I(N__25539));
    InMux I__2359 (
            .O(N__25542),
            .I(N__25536));
    LocalMux I__2358 (
            .O(N__25539),
            .I(\quad_counter0.a_delay_counter_8 ));
    LocalMux I__2357 (
            .O(N__25536),
            .I(\quad_counter0.a_delay_counter_8 ));
    CascadeMux I__2356 (
            .O(N__25531),
            .I(N__25527));
    InMux I__2355 (
            .O(N__25530),
            .I(N__25524));
    InMux I__2354 (
            .O(N__25527),
            .I(N__25521));
    LocalMux I__2353 (
            .O(N__25524),
            .I(\quad_counter0.a_delay_counter_1 ));
    LocalMux I__2352 (
            .O(N__25521),
            .I(\quad_counter0.a_delay_counter_1 ));
    InMux I__2351 (
            .O(N__25516),
            .I(N__25512));
    InMux I__2350 (
            .O(N__25515),
            .I(N__25509));
    LocalMux I__2349 (
            .O(N__25512),
            .I(\quad_counter0.a_delay_counter_6 ));
    LocalMux I__2348 (
            .O(N__25509),
            .I(\quad_counter0.a_delay_counter_6 ));
    InMux I__2347 (
            .O(N__25504),
            .I(N__25500));
    InMux I__2346 (
            .O(N__25503),
            .I(N__25497));
    LocalMux I__2345 (
            .O(N__25500),
            .I(\quad_counter0.a_delay_counter_9 ));
    LocalMux I__2344 (
            .O(N__25497),
            .I(\quad_counter0.a_delay_counter_9 ));
    InMux I__2343 (
            .O(N__25492),
            .I(N__25488));
    InMux I__2342 (
            .O(N__25491),
            .I(N__25485));
    LocalMux I__2341 (
            .O(N__25488),
            .I(\quad_counter0.a_delay_counter_7 ));
    LocalMux I__2340 (
            .O(N__25485),
            .I(\quad_counter0.a_delay_counter_7 ));
    CascadeMux I__2339 (
            .O(N__25480),
            .I(\quad_counter0.n18_cascade_ ));
    CascadeMux I__2338 (
            .O(N__25477),
            .I(N__25474));
    InMux I__2337 (
            .O(N__25474),
            .I(N__25469));
    InMux I__2336 (
            .O(N__25473),
            .I(N__25466));
    InMux I__2335 (
            .O(N__25472),
            .I(N__25463));
    LocalMux I__2334 (
            .O(N__25469),
            .I(a_delay_counter_0));
    LocalMux I__2333 (
            .O(N__25466),
            .I(a_delay_counter_0));
    LocalMux I__2332 (
            .O(N__25463),
            .I(a_delay_counter_0));
    CascadeMux I__2331 (
            .O(N__25456),
            .I(\quad_counter0.n20_cascade_ ));
    InMux I__2330 (
            .O(N__25453),
            .I(N__25449));
    InMux I__2329 (
            .O(N__25452),
            .I(N__25446));
    LocalMux I__2328 (
            .O(N__25449),
            .I(\quad_counter0.a_delay_counter_2 ));
    LocalMux I__2327 (
            .O(N__25446),
            .I(\quad_counter0.a_delay_counter_2 ));
    InMux I__2326 (
            .O(N__25441),
            .I(N__25435));
    InMux I__2325 (
            .O(N__25440),
            .I(N__25435));
    LocalMux I__2324 (
            .O(N__25435),
            .I(n11349));
    InMux I__2323 (
            .O(N__25432),
            .I(N__25428));
    InMux I__2322 (
            .O(N__25431),
            .I(N__25425));
    LocalMux I__2321 (
            .O(N__25428),
            .I(\quad_counter0.a_delay_counter_5 ));
    LocalMux I__2320 (
            .O(N__25425),
            .I(\quad_counter0.a_delay_counter_5 ));
    InMux I__2319 (
            .O(N__25420),
            .I(N__25416));
    InMux I__2318 (
            .O(N__25419),
            .I(N__25413));
    LocalMux I__2317 (
            .O(N__25416),
            .I(\quad_counter0.a_delay_counter_10 ));
    LocalMux I__2316 (
            .O(N__25413),
            .I(\quad_counter0.a_delay_counter_10 ));
    CascadeMux I__2315 (
            .O(N__25408),
            .I(N__25404));
    InMux I__2314 (
            .O(N__25407),
            .I(N__25401));
    InMux I__2313 (
            .O(N__25404),
            .I(N__25398));
    LocalMux I__2312 (
            .O(N__25401),
            .I(\quad_counter0.a_delay_counter_12 ));
    LocalMux I__2311 (
            .O(N__25398),
            .I(\quad_counter0.a_delay_counter_12 ));
    InMux I__2310 (
            .O(N__25393),
            .I(N__25389));
    InMux I__2309 (
            .O(N__25392),
            .I(N__25386));
    LocalMux I__2308 (
            .O(N__25389),
            .I(\quad_counter0.a_delay_counter_3 ));
    LocalMux I__2307 (
            .O(N__25386),
            .I(\quad_counter0.a_delay_counter_3 ));
    InMux I__2306 (
            .O(N__25381),
            .I(N__25378));
    LocalMux I__2305 (
            .O(N__25378),
            .I(\quad_counter0.n20954 ));
    InMux I__2304 (
            .O(N__25375),
            .I(N__25371));
    InMux I__2303 (
            .O(N__25374),
            .I(N__25368));
    LocalMux I__2302 (
            .O(N__25371),
            .I(\quad_counter0.a_delay_counter_4 ));
    LocalMux I__2301 (
            .O(N__25368),
            .I(\quad_counter0.a_delay_counter_4 ));
    InMux I__2300 (
            .O(N__25363),
            .I(N__25359));
    InMux I__2299 (
            .O(N__25362),
            .I(N__25356));
    LocalMux I__2298 (
            .O(N__25359),
            .I(\quad_counter0.a_delay_counter_11 ));
    LocalMux I__2297 (
            .O(N__25356),
            .I(\quad_counter0.a_delay_counter_11 ));
    CascadeMux I__2296 (
            .O(N__25351),
            .I(N__25347));
    InMux I__2295 (
            .O(N__25350),
            .I(N__25344));
    InMux I__2294 (
            .O(N__25347),
            .I(N__25341));
    LocalMux I__2293 (
            .O(N__25344),
            .I(\quad_counter0.a_delay_counter_14 ));
    LocalMux I__2292 (
            .O(N__25341),
            .I(\quad_counter0.a_delay_counter_14 ));
    InMux I__2291 (
            .O(N__25336),
            .I(N__25332));
    InMux I__2290 (
            .O(N__25335),
            .I(N__25329));
    LocalMux I__2289 (
            .O(N__25332),
            .I(\quad_counter0.a_delay_counter_13 ));
    LocalMux I__2288 (
            .O(N__25329),
            .I(\quad_counter0.a_delay_counter_13 ));
    InMux I__2287 (
            .O(N__25324),
            .I(N__25321));
    LocalMux I__2286 (
            .O(N__25321),
            .I(\quad_counter0.n19 ));
    SRMux I__2285 (
            .O(N__25318),
            .I(N__25315));
    LocalMux I__2284 (
            .O(N__25315),
            .I(N__25312));
    Span4Mux_h I__2283 (
            .O(N__25312),
            .I(N__25309));
    Odrv4 I__2282 (
            .O(N__25309),
            .I(\c0.n18649 ));
    SRMux I__2281 (
            .O(N__25306),
            .I(N__25303));
    LocalMux I__2280 (
            .O(N__25303),
            .I(\c0.n18639 ));
    SRMux I__2279 (
            .O(N__25300),
            .I(N__25297));
    LocalMux I__2278 (
            .O(N__25297),
            .I(N__25294));
    Span4Mux_v I__2277 (
            .O(N__25294),
            .I(N__25291));
    Odrv4 I__2276 (
            .O(N__25291),
            .I(\c0.n18663 ));
    SRMux I__2275 (
            .O(N__25288),
            .I(N__25285));
    LocalMux I__2274 (
            .O(N__25285),
            .I(N__25281));
    SRMux I__2273 (
            .O(N__25284),
            .I(N__25278));
    Span4Mux_h I__2272 (
            .O(N__25281),
            .I(N__25272));
    LocalMux I__2271 (
            .O(N__25278),
            .I(N__25272));
    InMux I__2270 (
            .O(N__25277),
            .I(N__25269));
    Odrv4 I__2269 (
            .O(N__25272),
            .I(a_delay_counter_15__N_2916));
    LocalMux I__2268 (
            .O(N__25269),
            .I(a_delay_counter_15__N_2916));
    InMux I__2267 (
            .O(N__25264),
            .I(N__25261));
    LocalMux I__2266 (
            .O(N__25261),
            .I(\quad_counter0.n13266 ));
    InMux I__2265 (
            .O(N__25258),
            .I(N__25253));
    InMux I__2264 (
            .O(N__25257),
            .I(N__25250));
    InMux I__2263 (
            .O(N__25256),
            .I(N__25247));
    LocalMux I__2262 (
            .O(N__25253),
            .I(\quad_counter0.b_delay_counter_14 ));
    LocalMux I__2261 (
            .O(N__25250),
            .I(\quad_counter0.b_delay_counter_14 ));
    LocalMux I__2260 (
            .O(N__25247),
            .I(\quad_counter0.b_delay_counter_14 ));
    InMux I__2259 (
            .O(N__25240),
            .I(N__25237));
    LocalMux I__2258 (
            .O(N__25237),
            .I(\quad_counter0.n13248 ));
    InMux I__2257 (
            .O(N__25234),
            .I(N__25229));
    InMux I__2256 (
            .O(N__25233),
            .I(N__25226));
    InMux I__2255 (
            .O(N__25232),
            .I(N__25223));
    LocalMux I__2254 (
            .O(N__25229),
            .I(N__25220));
    LocalMux I__2253 (
            .O(N__25226),
            .I(\quad_counter0.b_delay_counter_8 ));
    LocalMux I__2252 (
            .O(N__25223),
            .I(\quad_counter0.b_delay_counter_8 ));
    Odrv4 I__2251 (
            .O(N__25220),
            .I(\quad_counter0.b_delay_counter_8 ));
    InMux I__2250 (
            .O(N__25213),
            .I(N__25210));
    LocalMux I__2249 (
            .O(N__25210),
            .I(N__25207));
    Odrv4 I__2248 (
            .O(N__25207),
            .I(\quad_counter0.n13203 ));
    InMux I__2247 (
            .O(N__25204),
            .I(N__25199));
    InMux I__2246 (
            .O(N__25203),
            .I(N__25196));
    CascadeMux I__2245 (
            .O(N__25202),
            .I(N__25193));
    LocalMux I__2244 (
            .O(N__25199),
            .I(N__25188));
    LocalMux I__2243 (
            .O(N__25196),
            .I(N__25188));
    InMux I__2242 (
            .O(N__25193),
            .I(N__25185));
    Odrv4 I__2241 (
            .O(N__25188),
            .I(\quad_counter0.b_delay_counter_6 ));
    LocalMux I__2240 (
            .O(N__25185),
            .I(\quad_counter0.b_delay_counter_6 ));
    InMux I__2239 (
            .O(N__25180),
            .I(N__25176));
    InMux I__2238 (
            .O(N__25179),
            .I(N__25173));
    LocalMux I__2237 (
            .O(N__25176),
            .I(N__25167));
    LocalMux I__2236 (
            .O(N__25173),
            .I(N__25167));
    InMux I__2235 (
            .O(N__25172),
            .I(N__25164));
    Odrv4 I__2234 (
            .O(N__25167),
            .I(\quad_counter0.b_delay_counter_0 ));
    LocalMux I__2233 (
            .O(N__25164),
            .I(\quad_counter0.b_delay_counter_0 ));
    InMux I__2232 (
            .O(N__25159),
            .I(N__25156));
    LocalMux I__2231 (
            .O(N__25156),
            .I(\quad_counter0.n13251 ));
    InMux I__2230 (
            .O(N__25153),
            .I(N__25148));
    InMux I__2229 (
            .O(N__25152),
            .I(N__25145));
    InMux I__2228 (
            .O(N__25151),
            .I(N__25142));
    LocalMux I__2227 (
            .O(N__25148),
            .I(\quad_counter0.b_delay_counter_9 ));
    LocalMux I__2226 (
            .O(N__25145),
            .I(\quad_counter0.b_delay_counter_9 ));
    LocalMux I__2225 (
            .O(N__25142),
            .I(\quad_counter0.b_delay_counter_9 ));
    InMux I__2224 (
            .O(N__25135),
            .I(N__25132));
    LocalMux I__2223 (
            .O(N__25132),
            .I(N__25129));
    Odrv4 I__2222 (
            .O(N__25129),
            .I(\quad_counter0.n13194 ));
    InMux I__2221 (
            .O(N__25126),
            .I(N__25122));
    InMux I__2220 (
            .O(N__25125),
            .I(N__25119));
    LocalMux I__2219 (
            .O(N__25122),
            .I(N__25113));
    LocalMux I__2218 (
            .O(N__25119),
            .I(N__25113));
    InMux I__2217 (
            .O(N__25118),
            .I(N__25110));
    Odrv4 I__2216 (
            .O(N__25113),
            .I(\quad_counter0.b_delay_counter_3 ));
    LocalMux I__2215 (
            .O(N__25110),
            .I(\quad_counter0.b_delay_counter_3 ));
    InMux I__2214 (
            .O(N__25105),
            .I(N__25102));
    LocalMux I__2213 (
            .O(N__25102),
            .I(N__25099));
    Odrv4 I__2212 (
            .O(N__25099),
            .I(\quad_counter0.n13200 ));
    InMux I__2211 (
            .O(N__25096),
            .I(N__25092));
    InMux I__2210 (
            .O(N__25095),
            .I(N__25089));
    LocalMux I__2209 (
            .O(N__25092),
            .I(N__25083));
    LocalMux I__2208 (
            .O(N__25089),
            .I(N__25083));
    InMux I__2207 (
            .O(N__25088),
            .I(N__25080));
    Odrv12 I__2206 (
            .O(N__25083),
            .I(\quad_counter0.b_delay_counter_5 ));
    LocalMux I__2205 (
            .O(N__25080),
            .I(\quad_counter0.b_delay_counter_5 ));
    InMux I__2204 (
            .O(N__25075),
            .I(\quad_counter0.n17216 ));
    InMux I__2203 (
            .O(N__25072),
            .I(N__25068));
    InMux I__2202 (
            .O(N__25071),
            .I(N__25065));
    LocalMux I__2201 (
            .O(N__25068),
            .I(N__25059));
    LocalMux I__2200 (
            .O(N__25065),
            .I(N__25059));
    InMux I__2199 (
            .O(N__25064),
            .I(N__25056));
    Span4Mux_v I__2198 (
            .O(N__25059),
            .I(N__25051));
    LocalMux I__2197 (
            .O(N__25056),
            .I(N__25051));
    Odrv4 I__2196 (
            .O(N__25051),
            .I(\quad_counter0.b_delay_counter_11 ));
    InMux I__2195 (
            .O(N__25048),
            .I(N__25045));
    LocalMux I__2194 (
            .O(N__25045),
            .I(N__25042));
    Odrv12 I__2193 (
            .O(N__25042),
            .I(\quad_counter0.n13257 ));
    InMux I__2192 (
            .O(N__25039),
            .I(\quad_counter0.n17217 ));
    InMux I__2191 (
            .O(N__25036),
            .I(\quad_counter0.n17218 ));
    InMux I__2190 (
            .O(N__25033),
            .I(N__25028));
    InMux I__2189 (
            .O(N__25032),
            .I(N__25025));
    CascadeMux I__2188 (
            .O(N__25031),
            .I(N__25022));
    LocalMux I__2187 (
            .O(N__25028),
            .I(N__25017));
    LocalMux I__2186 (
            .O(N__25025),
            .I(N__25017));
    InMux I__2185 (
            .O(N__25022),
            .I(N__25014));
    Odrv4 I__2184 (
            .O(N__25017),
            .I(\quad_counter0.b_delay_counter_13 ));
    LocalMux I__2183 (
            .O(N__25014),
            .I(\quad_counter0.b_delay_counter_13 ));
    InMux I__2182 (
            .O(N__25009),
            .I(N__25006));
    LocalMux I__2181 (
            .O(N__25006),
            .I(N__25003));
    Odrv4 I__2180 (
            .O(N__25003),
            .I(\quad_counter0.n13263 ));
    InMux I__2179 (
            .O(N__25000),
            .I(\quad_counter0.n17219 ));
    InMux I__2178 (
            .O(N__24997),
            .I(\quad_counter0.n17220 ));
    InMux I__2177 (
            .O(N__24994),
            .I(\quad_counter0.n17221 ));
    InMux I__2176 (
            .O(N__24991),
            .I(N__24988));
    LocalMux I__2175 (
            .O(N__24988),
            .I(\quad_counter0.n13260 ));
    InMux I__2174 (
            .O(N__24985),
            .I(N__24980));
    InMux I__2173 (
            .O(N__24984),
            .I(N__24977));
    InMux I__2172 (
            .O(N__24983),
            .I(N__24974));
    LocalMux I__2171 (
            .O(N__24980),
            .I(\quad_counter0.b_delay_counter_12 ));
    LocalMux I__2170 (
            .O(N__24977),
            .I(\quad_counter0.b_delay_counter_12 ));
    LocalMux I__2169 (
            .O(N__24974),
            .I(\quad_counter0.b_delay_counter_12 ));
    InMux I__2168 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__2167 (
            .O(N__24964),
            .I(N__24961));
    Odrv4 I__2166 (
            .O(N__24961),
            .I(\quad_counter0.n13444 ));
    InMux I__2165 (
            .O(N__24958),
            .I(N__24955));
    LocalMux I__2164 (
            .O(N__24955),
            .I(\quad_counter0.n13182 ));
    InMux I__2163 (
            .O(N__24952),
            .I(\quad_counter0.n17207 ));
    InMux I__2162 (
            .O(N__24949),
            .I(\quad_counter0.n17208 ));
    InMux I__2161 (
            .O(N__24946),
            .I(\quad_counter0.n17209 ));
    InMux I__2160 (
            .O(N__24943),
            .I(N__24939));
    InMux I__2159 (
            .O(N__24942),
            .I(N__24936));
    LocalMux I__2158 (
            .O(N__24939),
            .I(N__24933));
    LocalMux I__2157 (
            .O(N__24936),
            .I(N__24929));
    Span4Mux_v I__2156 (
            .O(N__24933),
            .I(N__24926));
    InMux I__2155 (
            .O(N__24932),
            .I(N__24923));
    Span4Mux_v I__2154 (
            .O(N__24929),
            .I(N__24916));
    Span4Mux_h I__2153 (
            .O(N__24926),
            .I(N__24916));
    LocalMux I__2152 (
            .O(N__24923),
            .I(N__24916));
    Odrv4 I__2151 (
            .O(N__24916),
            .I(\quad_counter0.b_delay_counter_4 ));
    InMux I__2150 (
            .O(N__24913),
            .I(N__24910));
    LocalMux I__2149 (
            .O(N__24910),
            .I(N__24907));
    Span4Mux_h I__2148 (
            .O(N__24907),
            .I(N__24904));
    Odrv4 I__2147 (
            .O(N__24904),
            .I(\quad_counter0.n13197 ));
    InMux I__2146 (
            .O(N__24901),
            .I(\quad_counter0.n17210 ));
    InMux I__2145 (
            .O(N__24898),
            .I(\quad_counter0.n17211 ));
    InMux I__2144 (
            .O(N__24895),
            .I(\quad_counter0.n17212 ));
    CascadeMux I__2143 (
            .O(N__24892),
            .I(N__24887));
    InMux I__2142 (
            .O(N__24891),
            .I(N__24884));
    InMux I__2141 (
            .O(N__24890),
            .I(N__24881));
    InMux I__2140 (
            .O(N__24887),
            .I(N__24878));
    LocalMux I__2139 (
            .O(N__24884),
            .I(\quad_counter0.b_delay_counter_7 ));
    LocalMux I__2138 (
            .O(N__24881),
            .I(\quad_counter0.b_delay_counter_7 ));
    LocalMux I__2137 (
            .O(N__24878),
            .I(\quad_counter0.b_delay_counter_7 ));
    InMux I__2136 (
            .O(N__24871),
            .I(N__24868));
    LocalMux I__2135 (
            .O(N__24868),
            .I(\quad_counter0.n13214 ));
    InMux I__2134 (
            .O(N__24865),
            .I(\quad_counter0.n17213 ));
    InMux I__2133 (
            .O(N__24862),
            .I(bfn_9_15_0_));
    InMux I__2132 (
            .O(N__24859),
            .I(\quad_counter0.n17215 ));
    InMux I__2131 (
            .O(N__24856),
            .I(N__24850));
    InMux I__2130 (
            .O(N__24855),
            .I(N__24850));
    LocalMux I__2129 (
            .O(N__24850),
            .I(data_out_frame_5_1));
    CascadeMux I__2128 (
            .O(N__24847),
            .I(N__24844));
    InMux I__2127 (
            .O(N__24844),
            .I(N__24838));
    InMux I__2126 (
            .O(N__24843),
            .I(N__24838));
    LocalMux I__2125 (
            .O(N__24838),
            .I(data_out_frame_7_6));
    InMux I__2124 (
            .O(N__24835),
            .I(bfn_9_14_0_));
    InMux I__2123 (
            .O(N__24832),
            .I(N__24827));
    InMux I__2122 (
            .O(N__24831),
            .I(N__24824));
    InMux I__2121 (
            .O(N__24830),
            .I(N__24821));
    LocalMux I__2120 (
            .O(N__24827),
            .I(\quad_counter0.b_delay_counter_1 ));
    LocalMux I__2119 (
            .O(N__24824),
            .I(\quad_counter0.b_delay_counter_1 ));
    LocalMux I__2118 (
            .O(N__24821),
            .I(\quad_counter0.b_delay_counter_1 ));
    InMux I__2117 (
            .O(N__24814),
            .I(N__24808));
    InMux I__2116 (
            .O(N__24813),
            .I(N__24808));
    LocalMux I__2115 (
            .O(N__24808),
            .I(data_out_frame_6_6));
    InMux I__2114 (
            .O(N__24805),
            .I(\quad_counter0.n17236 ));
    InMux I__2113 (
            .O(N__24802),
            .I(\quad_counter0.n17227 ));
    InMux I__2112 (
            .O(N__24799),
            .I(\quad_counter0.n17228 ));
    InMux I__2111 (
            .O(N__24796),
            .I(bfn_9_8_0_));
    InMux I__2110 (
            .O(N__24793),
            .I(\quad_counter0.n17230 ));
    InMux I__2109 (
            .O(N__24790),
            .I(\quad_counter0.n17231 ));
    InMux I__2108 (
            .O(N__24787),
            .I(\quad_counter0.n17232 ));
    InMux I__2107 (
            .O(N__24784),
            .I(\quad_counter0.n17233 ));
    InMux I__2106 (
            .O(N__24781),
            .I(\quad_counter0.n17234 ));
    InMux I__2105 (
            .O(N__24778),
            .I(\quad_counter0.n17235 ));
    SRMux I__2104 (
            .O(N__24775),
            .I(N__24772));
    LocalMux I__2103 (
            .O(N__24772),
            .I(\c0.n18661 ));
    InMux I__2102 (
            .O(N__24769),
            .I(N__24766));
    LocalMux I__2101 (
            .O(N__24766),
            .I(n39));
    InMux I__2100 (
            .O(N__24763),
            .I(bfn_9_7_0_));
    InMux I__2099 (
            .O(N__24760),
            .I(\quad_counter0.n17222 ));
    InMux I__2098 (
            .O(N__24757),
            .I(\quad_counter0.n17223 ));
    InMux I__2097 (
            .O(N__24754),
            .I(\quad_counter0.n17224 ));
    InMux I__2096 (
            .O(N__24751),
            .I(\quad_counter0.n17225 ));
    InMux I__2095 (
            .O(N__24748),
            .I(\quad_counter0.n17226 ));
    IoInMux I__2094 (
            .O(N__24745),
            .I(N__24742));
    LocalMux I__2093 (
            .O(N__24742),
            .I(N__24739));
    Odrv4 I__2092 (
            .O(N__24739),
            .I(tx_enable));
    IoInMux I__2091 (
            .O(N__24736),
            .I(N__24733));
    LocalMux I__2090 (
            .O(N__24733),
            .I(N__24729));
    InMux I__2089 (
            .O(N__24732),
            .I(N__24726));
    IoSpan4Mux I__2088 (
            .O(N__24729),
            .I(N__24723));
    LocalMux I__2087 (
            .O(N__24726),
            .I(N__24720));
    Span4Mux_s3_v I__2086 (
            .O(N__24723),
            .I(N__24717));
    Span4Mux_h I__2085 (
            .O(N__24720),
            .I(N__24714));
    Sp12to4 I__2084 (
            .O(N__24717),
            .I(N__24711));
    Span4Mux_v I__2083 (
            .O(N__24714),
            .I(N__24708));
    Span12Mux_s11_v I__2082 (
            .O(N__24711),
            .I(N__24703));
    Sp12to4 I__2081 (
            .O(N__24708),
            .I(N__24703));
    Span12Mux_v I__2080 (
            .O(N__24703),
            .I(N__24700));
    Odrv12 I__2079 (
            .O(N__24700),
            .I(LED_c));
    SRMux I__2078 (
            .O(N__24697),
            .I(N__24694));
    LocalMux I__2077 (
            .O(N__24694),
            .I(N__24691));
    Span4Mux_h I__2076 (
            .O(N__24691),
            .I(N__24688));
    Odrv4 I__2075 (
            .O(N__24688),
            .I(\c0.n18673 ));
    IoInMux I__2074 (
            .O(N__24685),
            .I(N__24682));
    LocalMux I__2073 (
            .O(N__24682),
            .I(N__24679));
    IoSpan4Mux I__2072 (
            .O(N__24679),
            .I(N__24676));
    IoSpan4Mux I__2071 (
            .O(N__24676),
            .I(N__24673));
    IoSpan4Mux I__2070 (
            .O(N__24673),
            .I(N__24670));
    Odrv4 I__2069 (
            .O(N__24670),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\quad_counter1.n17321 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\quad_counter1.n17329 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\quad_counter1.n17337 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\quad_counter1.n17345 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\quad_counter0.n17289 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(\quad_counter0.n17297 ),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\quad_counter0.n17305 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\quad_counter0.n17313 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\quad_counter1.n17244 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\quad_counter1.n17259 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\quad_counter0.n17214 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\quad_counter0.n17229 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\c0.tx.n17281 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\c0.n17180_THRU_CRY_2_THRU_CO ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\c0.n17181_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\c0.n17182_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\c0.n17183_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\c0.n17184_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\c0.n17185_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\c0.n17186_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\c0.n17187_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\c0.n17188_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\c0.n17189_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\c0.n17190_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\c0.n17191_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\c0.n17192_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\c0.n17193_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\c0.n17194_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\c0.n17195_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\c0.n17196_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\c0.n17197_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\c0.n17198_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\c0.n17199_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\c0.n17200_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(\c0.n17201_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(\c0.n17202_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_14_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_29_0_ (
            .carryinitin(\c0.n17203_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_29_0_));
    defparam IN_MUX_bfv_14_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_30_0_ (
            .carryinitin(\c0.n17204_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_30_0_));
    defparam IN_MUX_bfv_14_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_31_0_ (
            .carryinitin(\c0.n17205_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_31_0_));
    defparam IN_MUX_bfv_14_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_32_0_ (
            .carryinitin(\c0.n17206_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__24685),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_2_3_5 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_2_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34182),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_49_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_49_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_49_LC_5_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_R_49_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24732),
            .lcout(\c0.rx.r_Rx_Data_R ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71000),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i0_LC_6_9_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i0_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i0_LC_6_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i0_LC_6_9_1  (
            .in0(N__35721),
            .in1(N__31127),
            .in2(_gnd_net_),
            .in3(N__25720),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71023),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i4_LC_7_13_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i4_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i4_LC_7_13_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i4_LC_7_13_7  (
            .in0(N__26595),
            .in1(N__26478),
            .in2(_gnd_net_),
            .in3(N__24913),
            .lcout(\quad_counter0.b_delay_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71001),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_delayed_62_LC_7_16_5 .C_ON=1'b0;
    defparam \quad_counter0.quadB_delayed_62_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadB_delayed_62_LC_7_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.quadB_delayed_62_LC_7_16_5  (
            .in0(N__26594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadB_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70991),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i9_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_7_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_7_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__29397),
            .in2(_gnd_net_),
            .in3(N__40555),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70993),
            .ce(),
            .sr(N__24697));
    defparam \c0.i1_2_lut_adj_924_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_924_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_924_LC_7_20_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_924_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__29396),
            .in2(_gnd_net_),
            .in3(N__41472),
            .lcout(\c0.n18673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_249_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_249_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_249_LC_7_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_249_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__27632),
            .in2(_gnd_net_),
            .in3(N__41449),
            .lcout(\c0.n18661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i15_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_7_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_7_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__27633),
            .in2(_gnd_net_),
            .in3(N__40554),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71007),
            .ce(),
            .sr(N__24775));
    defparam \quad_counter0.a_delay_counter__i0_LC_9_6_6 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i0_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i0_LC_9_6_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \quad_counter0.a_delay_counter__i0_LC_9_6_6  (
            .in0(N__25277),
            .in1(N__24769),
            .in2(N__25477),
            .in3(N__25616),
            .lcout(a_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71100),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_85_2_lut_LC_9_7_0 .C_ON=1'b1;
    defparam \quad_counter0.add_85_2_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_85_2_lut_LC_9_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_85_2_lut_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__25473),
            .in2(_gnd_net_),
            .in3(N__24763),
            .lcout(n39),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\quad_counter0.n17222 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i1_LC_9_7_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i1_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i1_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i1_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__25530),
            .in2(_gnd_net_),
            .in3(N__24760),
            .lcout(\quad_counter0.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n17222 ),
            .carryout(\quad_counter0.n17223 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i2_LC_9_7_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i2_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i2_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__25453),
            .in2(_gnd_net_),
            .in3(N__24757),
            .lcout(\quad_counter0.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n17223 ),
            .carryout(\quad_counter0.n17224 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i3_LC_9_7_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i3_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i3_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i3_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__25393),
            .in2(_gnd_net_),
            .in3(N__24754),
            .lcout(\quad_counter0.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n17224 ),
            .carryout(\quad_counter0.n17225 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i4_LC_9_7_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i4_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i4_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i4_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__25375),
            .in2(_gnd_net_),
            .in3(N__24751),
            .lcout(\quad_counter0.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n17225 ),
            .carryout(\quad_counter0.n17226 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i5_LC_9_7_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i5_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i5_LC_9_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i5_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__25432),
            .in2(_gnd_net_),
            .in3(N__24748),
            .lcout(\quad_counter0.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n17226 ),
            .carryout(\quad_counter0.n17227 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i6_LC_9_7_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i6_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i6_LC_9_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i6_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__25516),
            .in2(_gnd_net_),
            .in3(N__24802),
            .lcout(\quad_counter0.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n17227 ),
            .carryout(\quad_counter0.n17228 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i7_LC_9_7_7 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i7_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i7_LC_9_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i7_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__25492),
            .in2(_gnd_net_),
            .in3(N__24799),
            .lcout(\quad_counter0.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n17228 ),
            .carryout(\quad_counter0.n17229 ),
            .clk(N__71086),
            .ce(N__25617),
            .sr(N__25284));
    defparam \quad_counter0.a_delay_counter__i8_LC_9_8_0 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i8_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i8_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i8_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__25543),
            .in2(_gnd_net_),
            .in3(N__24796),
            .lcout(\quad_counter0.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\quad_counter0.n17230 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i9_LC_9_8_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i9_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i9_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i9_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__25504),
            .in2(_gnd_net_),
            .in3(N__24793),
            .lcout(\quad_counter0.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n17230 ),
            .carryout(\quad_counter0.n17231 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i10_LC_9_8_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i10_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i10_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i10_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__25420),
            .in2(_gnd_net_),
            .in3(N__24790),
            .lcout(\quad_counter0.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n17231 ),
            .carryout(\quad_counter0.n17232 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i11_LC_9_8_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i11_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i11_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i11_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__25363),
            .in2(_gnd_net_),
            .in3(N__24787),
            .lcout(\quad_counter0.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n17232 ),
            .carryout(\quad_counter0.n17233 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i12_LC_9_8_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i12_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i12_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i12_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__25407),
            .in2(_gnd_net_),
            .in3(N__24784),
            .lcout(\quad_counter0.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n17233 ),
            .carryout(\quad_counter0.n17234 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i13_LC_9_8_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i13_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i13_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i13_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__25336),
            .in2(_gnd_net_),
            .in3(N__24781),
            .lcout(\quad_counter0.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n17234 ),
            .carryout(\quad_counter0.n17235 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i14_LC_9_8_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i14_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i14_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i14_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__25350),
            .in2(_gnd_net_),
            .in3(N__24778),
            .lcout(\quad_counter0.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n17235 ),
            .carryout(\quad_counter0.n17236 ),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.a_delay_counter__i15_LC_9_8_7 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i15_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i15_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i15_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__25555),
            .in2(_gnd_net_),
            .in3(N__24805),
            .lcout(\quad_counter0.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71072),
            .ce(N__25624),
            .sr(N__25288));
    defparam \quad_counter0.B_delayed_68_LC_9_9_0 .C_ON=1'b0;
    defparam \quad_counter0.B_delayed_68_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_delayed_68_LC_9_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.B_delayed_68_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26928),
            .lcout(\quad_counter0.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71058),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.B_65_LC_9_9_1 .C_ON=1'b0;
    defparam \quad_counter0.B_65_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_65_LC_9_9_1 .LUT_INIT=16'b1011101010101000;
    LogicCell40 \quad_counter0.B_65_LC_9_9_1  (
            .in0(N__26927),
            .in1(N__26257),
            .in2(N__26494),
            .in3(N__26614),
            .lcout(B_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71058),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1060_1_lut_2_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \quad_counter0.i1060_1_lut_2_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1060_1_lut_2_lut_LC_9_9_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \quad_counter0.i1060_1_lut_2_lut_LC_9_9_2  (
            .in0(N__26881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26903),
            .lcout(\quad_counter0.n2228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.A_filtered_I_0_2_lut_LC_9_9_6  (
            .in0(N__26882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26904),
            .lcout(\quad_counter0.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i2_LC_9_9_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i2_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i2_LC_9_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i2_LC_9_9_7  (
            .in0(N__35720),
            .in1(N__25698),
            .in2(_gnd_net_),
            .in3(N__25681),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71058),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__2__5364_LC_9_10_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__2__5364_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__2__5364_LC_9_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_9__2__5364_LC_9_10_1  (
            .in0(N__25699),
            .in1(N__28473),
            .in2(_gnd_net_),
            .in3(N__46918),
            .lcout(data_out_frame_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71045),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i21_LC_9_10_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i21_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i21_LC_9_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i21_LC_9_10_2  (
            .in0(N__35731),
            .in1(N__33458),
            .in2(_gnd_net_),
            .in3(N__25801),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71045),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i18_LC_9_11_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i18_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i18_LC_9_11_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i18_LC_9_11_0  (
            .in0(N__35712),
            .in1(N__35756),
            .in2(_gnd_net_),
            .in3(N__25828),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i19_LC_9_11_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i19_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i19_LC_9_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i19_LC_9_11_1  (
            .in0(N__33002),
            .in1(N__35716),
            .in2(_gnd_net_),
            .in3(N__25819),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i20_LC_9_11_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i20_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i20_LC_9_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i20_LC_9_11_2  (
            .in0(N__35713),
            .in1(N__27107),
            .in2(_gnd_net_),
            .in3(N__25810),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i11_LC_9_11_3 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i11_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i11_LC_9_11_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i11_LC_9_11_3  (
            .in0(N__26613),
            .in1(N__26493),
            .in2(_gnd_net_),
            .in3(N__25048),
            .lcout(\quad_counter0.b_delay_counter_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i22_LC_9_11_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i22_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i22_LC_9_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i22_LC_9_11_4  (
            .in0(N__35714),
            .in1(N__25790),
            .in2(_gnd_net_),
            .in3(N__25771),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i23_LC_9_11_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i23_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i23_LC_9_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter0.count_i0_i23_LC_9_11_5  (
            .in0(N__25762),
            .in1(N__33965),
            .in2(_gnd_net_),
            .in3(N__35717),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i24_LC_9_11_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i24_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i24_LC_9_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i24_LC_9_11_6  (
            .in0(N__35715),
            .in1(N__32885),
            .in2(_gnd_net_),
            .in3(N__26011),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i25_LC_9_11_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i25_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i25_LC_9_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter0.count_i0_i25_LC_9_11_7  (
            .in0(N__26002),
            .in1(N__27149),
            .in2(_gnd_net_),
            .in3(N__35718),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71034),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__6__5384_LC_9_12_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__6__5384_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__6__5384_LC_9_12_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_out_frame_6__6__5384_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__46824),
            .in2(N__27055),
            .in3(N__24814),
            .lcout(data_out_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71024),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__1__5397_LC_9_12_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__1__5397_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__1__5397_LC_9_12_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame_5__1__5397_LC_9_12_1  (
            .in0(N__41059),
            .in1(N__24856),
            .in2(N__46904),
            .in3(_gnd_net_),
            .lcout(data_out_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71024),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_9_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_9_12_2  (
            .in0(N__24843),
            .in1(N__24813),
            .in2(_gnd_net_),
            .in3(N__40915),
            .lcout(\c0.n5_adj_3471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__3__5363_LC_9_12_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__3__5363_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__3__5363_LC_9_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_9__3__5363_LC_9_12_4  (
            .in0(N__33204),
            .in1(N__25672),
            .in2(_gnd_net_),
            .in3(N__46826),
            .lcout(data_out_frame_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71024),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17971_3_lut_LC_9_12_5 .C_ON=1'b0;
    defparam \c0.i17971_3_lut_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17971_3_lut_LC_9_12_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i17971_3_lut_LC_9_12_5  (
            .in0(N__40914),
            .in1(N__24855),
            .in2(_gnd_net_),
            .in3(N__36965),
            .lcout(\c0.n21559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__6__5376_LC_9_12_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__6__5376_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__6__5376_LC_9_12_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame_7__6__5376_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__46825),
            .in2(N__24847),
            .in3(N__25791),
            .lcout(data_out_frame_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71024),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_9_13_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_9_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_9_13_0  (
            .in0(N__27085),
            .in1(N__26962),
            .in2(_gnd_net_),
            .in3(N__40935),
            .lcout(\c0.n5_adj_3033 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i13_LC_9_13_1 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i13_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i13_LC_9_13_1 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \quad_counter0.b_delay_counter__i13_LC_9_13_1  (
            .in0(N__26615),
            .in1(N__25009),
            .in2(_gnd_net_),
            .in3(N__26483),
            .lcout(\quad_counter0.b_delay_counter_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71014),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i1_LC_9_13_2 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i1_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i1_LC_9_13_2 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \quad_counter0.b_delay_counter__i1_LC_9_13_2  (
            .in0(N__26482),
            .in1(N__24958),
            .in2(_gnd_net_),
            .in3(N__26616),
            .lcout(\quad_counter0.b_delay_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71014),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_LC_9_13_4 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_LC_9_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_LC_9_13_4  (
            .in0(N__26032),
            .in1(N__25064),
            .in2(N__24892),
            .in3(N__24932),
            .lcout(\quad_counter0.n27_adj_2992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_LC_9_13_5 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_LC_9_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_LC_9_13_5  (
            .in0(N__24830),
            .in1(N__26312),
            .in2(N__25031),
            .in3(N__25234),
            .lcout(\quad_counter0.n26_adj_2991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i7_LC_9_13_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i7_LC_9_13_7 .LUT_INIT=16'b1010000000001010;
    LogicCell40 \quad_counter0.b_delay_counter__i7_LC_9_13_7  (
            .in0(N__24871),
            .in1(_gnd_net_),
            .in2(N__26620),
            .in3(N__26484),
            .lcout(\quad_counter0.b_delay_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71014),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_2_lut_LC_9_14_0 .C_ON=1'b1;
    defparam \quad_counter0.add_86_2_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_2_lut_LC_9_14_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_2_lut_LC_9_14_0  (
            .in0(N__25180),
            .in1(N__25179),
            .in2(N__26227),
            .in3(N__24835),
            .lcout(\quad_counter0.n13444 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\quad_counter0.n17207 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_3_lut_LC_9_14_1 .C_ON=1'b1;
    defparam \quad_counter0.add_86_3_lut_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_3_lut_LC_9_14_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_3_lut_LC_9_14_1  (
            .in0(N__24832),
            .in1(N__24831),
            .in2(N__26231),
            .in3(N__24952),
            .lcout(\quad_counter0.n13182 ),
            .ltout(),
            .carryin(\quad_counter0.n17207 ),
            .carryout(\quad_counter0.n17208 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_4_lut_LC_9_14_2 .C_ON=1'b1;
    defparam \quad_counter0.add_86_4_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_4_lut_LC_9_14_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_4_lut_LC_9_14_2  (
            .in0(N__26374),
            .in1(N__26373),
            .in2(N__26228),
            .in3(N__24949),
            .lcout(\quad_counter0.n13187 ),
            .ltout(),
            .carryin(\quad_counter0.n17208 ),
            .carryout(\quad_counter0.n17209 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_5_lut_LC_9_14_3 .C_ON=1'b1;
    defparam \quad_counter0.add_86_5_lut_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_5_lut_LC_9_14_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_5_lut_LC_9_14_3  (
            .in0(N__25126),
            .in1(N__25125),
            .in2(N__26232),
            .in3(N__24946),
            .lcout(\quad_counter0.n13194 ),
            .ltout(),
            .carryin(\quad_counter0.n17209 ),
            .carryout(\quad_counter0.n17210 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_6_lut_LC_9_14_4 .C_ON=1'b1;
    defparam \quad_counter0.add_86_6_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_6_lut_LC_9_14_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_6_lut_LC_9_14_4  (
            .in0(N__24942),
            .in1(N__24943),
            .in2(N__26229),
            .in3(N__24901),
            .lcout(\quad_counter0.n13197 ),
            .ltout(),
            .carryin(\quad_counter0.n17210 ),
            .carryout(\quad_counter0.n17211 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_7_lut_LC_9_14_5 .C_ON=1'b1;
    defparam \quad_counter0.add_86_7_lut_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_7_lut_LC_9_14_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_7_lut_LC_9_14_5  (
            .in0(N__25096),
            .in1(N__25095),
            .in2(N__26233),
            .in3(N__24898),
            .lcout(\quad_counter0.n13200 ),
            .ltout(),
            .carryin(\quad_counter0.n17211 ),
            .carryout(\quad_counter0.n17212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_8_lut_LC_9_14_6 .C_ON=1'b1;
    defparam \quad_counter0.add_86_8_lut_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_8_lut_LC_9_14_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_8_lut_LC_9_14_6  (
            .in0(N__25204),
            .in1(N__25203),
            .in2(N__26230),
            .in3(N__24895),
            .lcout(\quad_counter0.n13203 ),
            .ltout(),
            .carryin(\quad_counter0.n17212 ),
            .carryout(\quad_counter0.n17213 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_9_lut_LC_9_14_7 .C_ON=1'b1;
    defparam \quad_counter0.add_86_9_lut_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_9_lut_LC_9_14_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_9_lut_LC_9_14_7  (
            .in0(N__24891),
            .in1(N__24890),
            .in2(N__26234),
            .in3(N__24865),
            .lcout(\quad_counter0.n13214 ),
            .ltout(),
            .carryin(\quad_counter0.n17213 ),
            .carryout(\quad_counter0.n17214 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_10_lut_LC_9_15_0 .C_ON=1'b1;
    defparam \quad_counter0.add_86_10_lut_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_10_lut_LC_9_15_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_10_lut_LC_9_15_0  (
            .in0(N__25233),
            .in1(N__25232),
            .in2(N__26235),
            .in3(N__24862),
            .lcout(\quad_counter0.n13248 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\quad_counter0.n17215 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_11_lut_LC_9_15_1 .C_ON=1'b1;
    defparam \quad_counter0.add_86_11_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_11_lut_LC_9_15_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_11_lut_LC_9_15_1  (
            .in0(N__25153),
            .in1(N__25152),
            .in2(N__26239),
            .in3(N__24859),
            .lcout(\quad_counter0.n13251 ),
            .ltout(),
            .carryin(\quad_counter0.n17215 ),
            .carryout(\quad_counter0.n17216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_12_lut_LC_9_15_2 .C_ON=1'b1;
    defparam \quad_counter0.add_86_12_lut_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_12_lut_LC_9_15_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_12_lut_LC_9_15_2  (
            .in0(N__26031),
            .in1(N__26030),
            .in2(N__26236),
            .in3(N__25075),
            .lcout(\quad_counter0.n13254 ),
            .ltout(),
            .carryin(\quad_counter0.n17216 ),
            .carryout(\quad_counter0.n17217 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_13_lut_LC_9_15_3 .C_ON=1'b1;
    defparam \quad_counter0.add_86_13_lut_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_13_lut_LC_9_15_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_13_lut_LC_9_15_3  (
            .in0(N__25072),
            .in1(N__25071),
            .in2(N__26240),
            .in3(N__25039),
            .lcout(\quad_counter0.n13257 ),
            .ltout(),
            .carryin(\quad_counter0.n17217 ),
            .carryout(\quad_counter0.n17218 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_14_lut_LC_9_15_4 .C_ON=1'b1;
    defparam \quad_counter0.add_86_14_lut_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_14_lut_LC_9_15_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_14_lut_LC_9_15_4  (
            .in0(N__24985),
            .in1(N__24984),
            .in2(N__26237),
            .in3(N__25036),
            .lcout(\quad_counter0.n13260 ),
            .ltout(),
            .carryin(\quad_counter0.n17218 ),
            .carryout(\quad_counter0.n17219 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_15_lut_LC_9_15_5 .C_ON=1'b1;
    defparam \quad_counter0.add_86_15_lut_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_15_lut_LC_9_15_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_15_lut_LC_9_15_5  (
            .in0(N__25033),
            .in1(N__25032),
            .in2(N__26241),
            .in3(N__25000),
            .lcout(\quad_counter0.n13263 ),
            .ltout(),
            .carryin(\quad_counter0.n17219 ),
            .carryout(\quad_counter0.n17220 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_16_lut_LC_9_15_6 .C_ON=1'b1;
    defparam \quad_counter0.add_86_16_lut_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_16_lut_LC_9_15_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_16_lut_LC_9_15_6  (
            .in0(N__25258),
            .in1(N__25257),
            .in2(N__26238),
            .in3(N__24997),
            .lcout(\quad_counter0.n13266 ),
            .ltout(),
            .carryin(\quad_counter0.n17220 ),
            .carryout(\quad_counter0.n17221 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_86_17_lut_LC_9_15_7 .C_ON=1'b0;
    defparam \quad_counter0.add_86_17_lut_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_86_17_lut_LC_9_15_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.add_86_17_lut_LC_9_15_7  (
            .in0(N__26313),
            .in1(N__26314),
            .in2(N__26242),
            .in3(N__24994),
            .lcout(\quad_counter0.n13269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i12_LC_9_16_0 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i12_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i12_LC_9_16_0 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i12_LC_9_16_0  (
            .in0(N__26604),
            .in1(N__26486),
            .in2(_gnd_net_),
            .in3(N__24991),
            .lcout(\quad_counter0.b_delay_counter_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_LC_9_16_1 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_LC_9_16_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i12_4_lut_LC_9_16_1  (
            .in0(N__25256),
            .in1(N__24983),
            .in2(N__26366),
            .in3(N__25088),
            .lcout(\quad_counter0.n28_adj_2990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i0_LC_9_16_2 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i0_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i0_LC_9_16_2 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i0_LC_9_16_2  (
            .in0(N__26603),
            .in1(N__26485),
            .in2(_gnd_net_),
            .in3(N__24967),
            .lcout(\quad_counter0.b_delay_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i14_LC_9_16_3 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i14_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i14_LC_9_16_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i14_LC_9_16_3  (
            .in0(N__26488),
            .in1(N__26605),
            .in2(_gnd_net_),
            .in3(N__25264),
            .lcout(\quad_counter0.b_delay_counter_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i8_LC_9_16_4 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i8_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i8_LC_9_16_4 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i8_LC_9_16_4  (
            .in0(N__26607),
            .in1(N__26487),
            .in2(_gnd_net_),
            .in3(N__25240),
            .lcout(\quad_counter0.b_delay_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i6_LC_9_16_5 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i6_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i6_LC_9_16_5 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i6_LC_9_16_5  (
            .in0(N__26489),
            .in1(N__26606),
            .in2(_gnd_net_),
            .in3(N__25213),
            .lcout(\quad_counter0.b_delay_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_206_LC_9_16_6 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_206_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_206_LC_9_16_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter0.i9_4_lut_adj_206_LC_9_16_6  (
            .in0(N__25151),
            .in1(N__25118),
            .in2(N__25202),
            .in3(N__25172),
            .lcout(\quad_counter0.n25_adj_2993 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i9_LC_9_16_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i9_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i9_LC_9_16_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i9_LC_9_16_7  (
            .in0(N__26490),
            .in1(N__26608),
            .in2(_gnd_net_),
            .in3(N__25159),
            .lcout(\quad_counter0.b_delay_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70995),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i3_LC_9_17_1 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i3_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i3_LC_9_17_1 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i3_LC_9_17_1  (
            .in0(N__26541),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(N__25135),
            .lcout(\quad_counter0.b_delay_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70992),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i5_LC_9_17_5 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i5_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i5_LC_9_17_5 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i5_LC_9_17_5  (
            .in0(N__26542),
            .in1(N__26492),
            .in2(_gnd_net_),
            .in3(N__25105),
            .lcout(\quad_counter0.b_delay_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70992),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_9_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__29624),
            .in2(_gnd_net_),
            .in3(N__40542),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70996),
            .ce(),
            .sr(N__25318));
    defparam \c0.i1_2_lut_adj_435_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_435_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_435_LC_9_19_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_435_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__29816),
            .in2(_gnd_net_),
            .in3(N__41471),
            .lcout(\c0.n18639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_368_LC_9_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_368_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_368_LC_9_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_368_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__29618),
            .in2(_gnd_net_),
            .in3(N__41470),
            .lcout(\c0.n18649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i27_LC_9_20_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_9_20_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_9_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__40544),
            .in2(_gnd_net_),
            .in3(N__29817),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71008),
            .ce(),
            .sr(N__25306));
    defparam \c0.i1_2_lut_adj_247_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_247_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_247_LC_9_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_247_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__29423),
            .in2(_gnd_net_),
            .in3(N__41393),
            .lcout(\c0.n18663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i14_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_9_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_9_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__29424),
            .in2(_gnd_net_),
            .in3(N__40540),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71025),
            .ce(),
            .sr(N__25300));
    defparam \c0.i1_2_lut_adj_258_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_258_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_258_LC_9_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_258_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__27611),
            .in2(_gnd_net_),
            .in3(N__41469),
            .lcout(\c0.n18671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_9_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__40541),
            .in2(_gnd_net_),
            .in3(N__29771),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71046),
            .ce(),
            .sr(N__27952));
    defparam \quad_counter1.quadA_delayed_61_LC_10_4_3 .C_ON=1'b0;
    defparam \quad_counter1.quadA_delayed_61_LC_10_4_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadA_delayed_61_LC_10_4_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter1.quadA_delayed_61_LC_10_4_3  (
            .in0(N__28206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadA_delayed_adj_3584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71131),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_10_6_0 .C_ON=1'b0;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadA_I_0_73_2_lut_LC_10_6_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.quadA_I_0_73_2_lut_LC_10_6_0  (
            .in0(N__25598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25565),
            .lcout(a_delay_counter_15__N_2916),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_63_LC_10_6_2 .C_ON=1'b0;
    defparam \quad_counter0.A_63_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_63_LC_10_6_2 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \quad_counter0.A_63_LC_10_6_2  (
            .in0(N__25441),
            .in1(N__25567),
            .in2(N__25600),
            .in3(N__26880),
            .lcout(A_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71101),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_10_6_3.C_ON=1'b0;
    defparam i1_3_lut_LC_10_6_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_10_6_3.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_LC_10_6_3 (
            .in0(N__25566),
            .in1(N__25594),
            .in2(_gnd_net_),
            .in3(N__25440),
            .lcout(n12447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_delayed_61_LC_10_6_6 .C_ON=1'b0;
    defparam \quad_counter0.quadA_delayed_61_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadA_delayed_61_LC_10_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.quadA_delayed_61_LC_10_6_6  (
            .in0(N__25599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadA_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71101),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i7_4_lut_LC_10_7_0 .C_ON=1'b0;
    defparam \quad_counter0.i7_4_lut_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i7_4_lut_LC_10_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i7_4_lut_LC_10_7_0  (
            .in0(N__25554),
            .in1(N__25542),
            .in2(N__25531),
            .in3(N__25515),
            .lcout(),
            .ltout(\quad_counter0.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_LC_10_7_1 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_LC_10_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i9_4_lut_LC_10_7_1  (
            .in0(N__25503),
            .in1(N__25491),
            .in2(N__25480),
            .in3(N__25381),
            .lcout(),
            .ltout(\quad_counter0.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_4_lut_LC_10_7_2 .C_ON=1'b0;
    defparam \quad_counter0.i2_4_lut_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_4_lut_LC_10_7_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \quad_counter0.i2_4_lut_LC_10_7_2  (
            .in0(N__25324),
            .in1(N__25472),
            .in2(N__25456),
            .in3(N__25452),
            .lcout(n11349),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_adj_205_LC_10_7_5 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_adj_205_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_adj_205_LC_10_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i3_4_lut_adj_205_LC_10_7_5  (
            .in0(N__25431),
            .in1(N__25419),
            .in2(N__25408),
            .in3(N__25392),
            .lcout(\quad_counter0.n20954 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i1_LC_10_8_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i1_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i1_LC_10_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i1_LC_10_8_5  (
            .in0(N__35640),
            .in1(N__27326),
            .in2(_gnd_net_),
            .in3(N__25708),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71073),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_LC_10_8_6 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_LC_10_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_LC_10_8_6  (
            .in0(N__25374),
            .in1(N__25362),
            .in2(N__25351),
            .in3(N__25335),
            .lcout(\quad_counter0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i3_LC_10_8_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i3_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i3_LC_10_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i3_LC_10_8_7  (
            .in0(N__35641),
            .in1(N__25661),
            .in2(_gnd_net_),
            .in3(N__25642),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71073),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_1_LC_10_9_0 .C_ON=1'b1;
    defparam \quad_counter0.add_601_1_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_1_LC_10_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter0.add_601_1_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__25895),
            .in2(N__25955),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\quad_counter0.n17282 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_2_lut_LC_10_9_1 .C_ON=1'b1;
    defparam \quad_counter0.add_601_2_lut_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_2_lut_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_2_lut_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__25726),
            .in2(N__31140),
            .in3(N__25711),
            .lcout(n2279),
            .ltout(),
            .carryin(\quad_counter0.n17282 ),
            .carryout(\quad_counter0.n17283 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_3_lut_LC_10_9_2 .C_ON=1'b1;
    defparam \quad_counter0.add_601_3_lut_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_3_lut_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_3_lut_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__25896),
            .in2(N__27327),
            .in3(N__25702),
            .lcout(n2278),
            .ltout(),
            .carryin(\quad_counter0.n17283 ),
            .carryout(\quad_counter0.n17284 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_4_lut_LC_10_9_3 .C_ON=1'b1;
    defparam \quad_counter0.add_601_4_lut_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_4_lut_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_4_lut_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__25697),
            .in2(N__25954),
            .in3(N__25675),
            .lcout(n2277),
            .ltout(),
            .carryin(\quad_counter0.n17284 ),
            .carryout(\quad_counter0.n17285 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_5_lut_LC_10_9_4 .C_ON=1'b1;
    defparam \quad_counter0.add_601_5_lut_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_5_lut_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_5_lut_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__25900),
            .in2(N__25671),
            .in3(N__25636),
            .lcout(n2276),
            .ltout(),
            .carryin(\quad_counter0.n17285 ),
            .carryout(\quad_counter0.n17286 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_6_lut_LC_10_9_5 .C_ON=1'b1;
    defparam \quad_counter0.add_601_6_lut_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_6_lut_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_6_lut_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__25905),
            .in2(N__27211),
            .in3(N__25633),
            .lcout(n2275),
            .ltout(),
            .carryin(\quad_counter0.n17286 ),
            .carryout(\quad_counter0.n17287 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_7_lut_LC_10_9_6 .C_ON=1'b1;
    defparam \quad_counter0.add_601_7_lut_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_7_lut_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_7_lut_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__25901),
            .in2(N__26074),
            .in3(N__25630),
            .lcout(n2274),
            .ltout(),
            .carryin(\quad_counter0.n17287 ),
            .carryout(\quad_counter0.n17288 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_8_lut_LC_10_9_7 .C_ON=1'b1;
    defparam \quad_counter0.add_601_8_lut_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_8_lut_LC_10_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_8_lut_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__25906),
            .in2(N__27442),
            .in3(N__25627),
            .lcout(n2273),
            .ltout(),
            .carryin(\quad_counter0.n17288 ),
            .carryout(\quad_counter0.n17289 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_9_lut_LC_10_10_0 .C_ON=1'b1;
    defparam \quad_counter0.add_601_9_lut_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_9_lut_LC_10_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_9_lut_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__25907),
            .in2(N__27403),
            .in3(N__25753),
            .lcout(n2272),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\quad_counter0.n17290 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_10_lut_LC_10_10_1 .C_ON=1'b1;
    defparam \quad_counter0.add_601_10_lut_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_10_lut_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_10_lut_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__25911),
            .in2(N__30721),
            .in3(N__25750),
            .lcout(n2271),
            .ltout(),
            .carryin(\quad_counter0.n17290 ),
            .carryout(\quad_counter0.n17291 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_11_lut_LC_10_10_2 .C_ON=1'b1;
    defparam \quad_counter0.add_601_11_lut_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_11_lut_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_11_lut_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__25908),
            .in2(N__30790),
            .in3(N__25747),
            .lcout(n2270),
            .ltout(),
            .carryin(\quad_counter0.n17291 ),
            .carryout(\quad_counter0.n17292 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_12_lut_LC_10_10_3 .C_ON=1'b1;
    defparam \quad_counter0.add_601_12_lut_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_12_lut_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_12_lut_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__25912),
            .in2(N__27130),
            .in3(N__25744),
            .lcout(n2269),
            .ltout(),
            .carryin(\quad_counter0.n17292 ),
            .carryout(\quad_counter0.n17293 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_13_lut_LC_10_10_4 .C_ON=1'b1;
    defparam \quad_counter0.add_601_13_lut_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_13_lut_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_13_lut_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__25909),
            .in2(N__33258),
            .in3(N__25741),
            .lcout(n2268),
            .ltout(),
            .carryin(\quad_counter0.n17293 ),
            .carryout(\quad_counter0.n17294 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_14_lut_LC_10_10_5 .C_ON=1'b1;
    defparam \quad_counter0.add_601_14_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_14_lut_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_14_lut_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__25913),
            .in2(N__28842),
            .in3(N__25738),
            .lcout(n2267),
            .ltout(),
            .carryin(\quad_counter0.n17294 ),
            .carryout(\quad_counter0.n17295 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_15_lut_LC_10_10_6 .C_ON=1'b1;
    defparam \quad_counter0.add_601_15_lut_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_15_lut_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_15_lut_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__25910),
            .in2(N__28674),
            .in3(N__25735),
            .lcout(n2266),
            .ltout(),
            .carryin(\quad_counter0.n17295 ),
            .carryout(\quad_counter0.n17296 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_16_lut_LC_10_10_7 .C_ON=1'b1;
    defparam \quad_counter0.add_601_16_lut_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_16_lut_LC_10_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_16_lut_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__25914),
            .in2(N__27249),
            .in3(N__25732),
            .lcout(n2265),
            .ltout(),
            .carryin(\quad_counter0.n17296 ),
            .carryout(\quad_counter0.n17297 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_17_lut_LC_10_11_0 .C_ON=1'b1;
    defparam \quad_counter0.add_601_17_lut_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_17_lut_LC_10_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_17_lut_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__25956),
            .in2(N__27003),
            .in3(N__25729),
            .lcout(n2264),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\quad_counter0.n17298 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_18_lut_LC_10_11_1 .C_ON=1'b1;
    defparam \quad_counter0.add_601_18_lut_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_18_lut_LC_10_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_18_lut_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__25959),
            .in2(N__27273),
            .in3(N__25834),
            .lcout(n2263),
            .ltout(),
            .carryin(\quad_counter0.n17298 ),
            .carryout(\quad_counter0.n17299 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_19_lut_LC_10_11_2 .C_ON=1'b1;
    defparam \quad_counter0.add_601_19_lut_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_19_lut_LC_10_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_19_lut_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__28721),
            .in2(N__25977),
            .in3(N__25831),
            .lcout(n2262),
            .ltout(),
            .carryin(\quad_counter0.n17299 ),
            .carryout(\quad_counter0.n17300 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_20_lut_LC_10_11_3 .C_ON=1'b1;
    defparam \quad_counter0.add_601_20_lut_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_20_lut_LC_10_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_20_lut_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__25963),
            .in2(N__35760),
            .in3(N__25822),
            .lcout(n2261),
            .ltout(),
            .carryin(\quad_counter0.n17300 ),
            .carryout(\quad_counter0.n17301 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_21_lut_LC_10_11_4 .C_ON=1'b1;
    defparam \quad_counter0.add_601_21_lut_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_21_lut_LC_10_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_21_lut_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__25957),
            .in2(N__33003),
            .in3(N__25813),
            .lcout(n2260),
            .ltout(),
            .carryin(\quad_counter0.n17301 ),
            .carryout(\quad_counter0.n17302 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_22_lut_LC_10_11_5 .C_ON=1'b1;
    defparam \quad_counter0.add_601_22_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_22_lut_LC_10_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_22_lut_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__25964),
            .in2(N__27108),
            .in3(N__25804),
            .lcout(n2259),
            .ltout(),
            .carryin(\quad_counter0.n17302 ),
            .carryout(\quad_counter0.n17303 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_23_lut_LC_10_11_6 .C_ON=1'b1;
    defparam \quad_counter0.add_601_23_lut_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_23_lut_LC_10_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_23_lut_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__25958),
            .in2(N__33462),
            .in3(N__25795),
            .lcout(n2258),
            .ltout(),
            .carryin(\quad_counter0.n17303 ),
            .carryout(\quad_counter0.n17304 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_24_lut_LC_10_11_7 .C_ON=1'b1;
    defparam \quad_counter0.add_601_24_lut_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_24_lut_LC_10_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_24_lut_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__25965),
            .in2(N__25792),
            .in3(N__25765),
            .lcout(n2257),
            .ltout(),
            .carryin(\quad_counter0.n17304 ),
            .carryout(\quad_counter0.n17305 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_25_lut_LC_10_12_0 .C_ON=1'b1;
    defparam \quad_counter0.add_601_25_lut_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_25_lut_LC_10_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_25_lut_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__25966),
            .in2(N__33969),
            .in3(N__25756),
            .lcout(n2256),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\quad_counter0.n17306 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_26_lut_LC_10_12_1 .C_ON=1'b1;
    defparam \quad_counter0.add_601_26_lut_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_26_lut_LC_10_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_26_lut_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__25970),
            .in2(N__32889),
            .in3(N__26005),
            .lcout(n2255),
            .ltout(),
            .carryin(\quad_counter0.n17306 ),
            .carryout(\quad_counter0.n17307 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_27_lut_LC_10_12_2 .C_ON=1'b1;
    defparam \quad_counter0.add_601_27_lut_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_27_lut_LC_10_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_27_lut_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__25967),
            .in2(N__27153),
            .in3(N__25996),
            .lcout(n2254),
            .ltout(),
            .carryin(\quad_counter0.n17307 ),
            .carryout(\quad_counter0.n17308 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_28_lut_LC_10_12_3 .C_ON=1'b1;
    defparam \quad_counter0.add_601_28_lut_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_28_lut_LC_10_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_28_lut_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__25971),
            .in2(N__35895),
            .in3(N__25993),
            .lcout(n2253),
            .ltout(),
            .carryin(\quad_counter0.n17308 ),
            .carryout(\quad_counter0.n17309 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_29_lut_LC_10_12_4 .C_ON=1'b1;
    defparam \quad_counter0.add_601_29_lut_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_29_lut_LC_10_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_29_lut_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__25968),
            .in2(N__35547),
            .in3(N__25990),
            .lcout(n2252),
            .ltout(),
            .carryin(\quad_counter0.n17309 ),
            .carryout(\quad_counter0.n17310 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_30_lut_LC_10_12_5 .C_ON=1'b1;
    defparam \quad_counter0.add_601_30_lut_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_30_lut_LC_10_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_30_lut_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__25972),
            .in2(N__27297),
            .in3(N__25987),
            .lcout(n2251),
            .ltout(),
            .carryin(\quad_counter0.n17310 ),
            .carryout(\quad_counter0.n17311 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_31_lut_LC_10_12_6 .C_ON=1'b1;
    defparam \quad_counter0.add_601_31_lut_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_31_lut_LC_10_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_31_lut_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__25969),
            .in2(N__33354),
            .in3(N__25984),
            .lcout(n2250),
            .ltout(),
            .carryin(\quad_counter0.n17311 ),
            .carryout(\quad_counter0.n17312 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_32_lut_LC_10_12_7 .C_ON=1'b1;
    defparam \quad_counter0.add_601_32_lut_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_32_lut_LC_10_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_601_32_lut_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(N__25973),
            .in2(N__27051),
            .in3(N__25981),
            .lcout(n2249),
            .ltout(),
            .carryin(\quad_counter0.n17312 ),
            .carryout(\quad_counter0.n17313 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_601_33_lut_LC_10_13_0 .C_ON=1'b0;
    defparam \quad_counter0.add_601_33_lut_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_601_33_lut_LC_10_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.add_601_33_lut_LC_10_13_0  (
            .in0(N__43454),
            .in1(N__25978),
            .in2(_gnd_net_),
            .in3(N__25837),
            .lcout(n2248),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__0__5350_LC_10_13_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__0__5350_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__0__5350_LC_10_13_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_11__0__5350_LC_10_13_1  (
            .in0(N__30121),
            .in1(N__33606),
            .in2(_gnd_net_),
            .in3(N__46903),
            .lcout(data_out_frame_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i4_LC_10_13_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i4_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i4_LC_10_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i4_LC_10_13_2  (
            .in0(N__35709),
            .in1(N__27203),
            .in2(_gnd_net_),
            .in3(N__26119),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__3__5203_LC_10_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__3__5203_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__3__5203_LC_10_13_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.data_out_frame_29__3__5203_LC_10_13_3  (
            .in0(N__36033),
            .in1(N__46889),
            .in2(_gnd_net_),
            .in3(N__50362),
            .lcout(data_out_frame_29_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i7_LC_10_13_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i7_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i7_LC_10_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i7_LC_10_13_5  (
            .in0(N__27398),
            .in1(N__35711),
            .in2(_gnd_net_),
            .in3(N__26107),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i5_LC_10_13_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i5_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i5_LC_10_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \quad_counter0.count_i0_i5_LC_10_13_6  (
            .in0(N__35710),
            .in1(_gnd_net_),
            .in2(N__26073),
            .in3(N__26098),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i31_LC_10_13_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i31_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i31_LC_10_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i31_LC_10_13_7  (
            .in0(N__35719),
            .in1(N__43455),
            .in2(_gnd_net_),
            .in3(N__26089),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71016),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17718_4_lut_LC_10_14_1 .C_ON=1'b0;
    defparam \c0.i17718_4_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17718_4_lut_LC_10_14_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i17718_4_lut_LC_10_14_1  (
            .in0(N__26083),
            .in1(N__36953),
            .in2(N__33430),
            .in3(N__36700),
            .lcout(\c0.n21305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__5__5361_LC_10_14_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__5__5361_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__5__5361_LC_10_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_9__5__5361_LC_10_14_5  (
            .in0(N__26069),
            .in1(N__33102),
            .in2(_gnd_net_),
            .in3(N__46901),
            .lcout(data_out_frame_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71010),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21629_bdd_4_lut_LC_10_14_6 .C_ON=1'b0;
    defparam \c0.n21629_bdd_4_lut_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.n21629_bdd_4_lut_LC_10_14_6 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n21629_bdd_4_lut_LC_10_14_6  (
            .in0(N__36699),
            .in1(N__26046),
            .in2(N__27226),
            .in3(N__26125),
            .lcout(\c0.n21632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__6__5360_LC_10_14_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__6__5360_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__6__5360_LC_10_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_9__6__5360_LC_10_14_7  (
            .in0(N__26047),
            .in1(N__27435),
            .in2(_gnd_net_),
            .in3(N__46902),
            .lcout(data_out_frame_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71010),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i10_LC_10_15_1 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i10_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i10_LC_10_15_1 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i10_LC_10_15_1  (
            .in0(N__26473),
            .in1(N__26610),
            .in2(_gnd_net_),
            .in3(N__26038),
            .lcout(\quad_counter0.b_delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71003),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i15_LC_10_15_3 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i15_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i15_LC_10_15_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i15_LC_10_15_3  (
            .in0(N__26474),
            .in1(N__26611),
            .in2(_gnd_net_),
            .in3(N__26320),
            .lcout(\quad_counter0.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71003),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__6__5352_LC_10_15_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__6__5352_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__6__5352_LC_10_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__6__5352_LC_10_15_4  (
            .in0(N__30646),
            .in1(N__26134),
            .in2(_gnd_net_),
            .in3(N__46723),
            .lcout(data_out_frame_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71003),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_LC_10_15_5 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_LC_10_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_LC_10_15_5  (
            .in0(N__26290),
            .in1(N__26281),
            .in2(N__26272),
            .in3(N__26263),
            .lcout(n11347),
            .ltout(n11347_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i18016_4_lut_3_lut_LC_10_15_6 .C_ON=1'b0;
    defparam \quad_counter0.i18016_4_lut_3_lut_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i18016_4_lut_3_lut_LC_10_15_6 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \quad_counter0.i18016_4_lut_3_lut_LC_10_15_6  (
            .in0(N__26612),
            .in1(_gnd_net_),
            .in2(N__26245),
            .in3(N__26472),
            .lcout(\quad_counter0.n21603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18044_LC_10_15_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18044_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18044_LC_10_15_7 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18044_LC_10_15_7  (
            .in0(N__26133),
            .in1(N__40857),
            .in2(N__28651),
            .in3(N__36701),
            .lcout(\c0.n21629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_10_16_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_10_16_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_10_16_0  (
            .in0(N__29282),
            .in1(N__29145),
            .in2(_gnd_net_),
            .in3(N__27556),
            .lcout(\c0.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70998),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__4__5354_LC_10_16_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__4__5354_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__4__5354_LC_10_16_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__4__5354_LC_10_16_1  (
            .in0(N__36082),
            .in1(N__27472),
            .in2(_gnd_net_),
            .in3(N__46939),
            .lcout(data_out_frame_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70998),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__7__5367_LC_10_16_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__7__5367_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__7__5367_LC_10_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__7__5367_LC_10_16_2  (
            .in0(N__46938),
            .in1(N__27004),
            .in2(_gnd_net_),
            .in3(N__27168),
            .lcout(data_out_frame_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70998),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_10_16_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_10_16_3 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_10_16_3  (
            .in0(N__29328),
            .in1(N__34065),
            .in2(N__29163),
            .in3(N__27523),
            .lcout(\c0.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70998),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i2_LC_10_16_6 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i2_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i2_LC_10_16_6 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \quad_counter0.b_delay_counter__i2_LC_10_16_6  (
            .in0(N__26609),
            .in1(N__26471),
            .in2(_gnd_net_),
            .in3(N__26383),
            .lcout(\quad_counter0.b_delay_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70998),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i17744_3_lut_LC_10_17_0 .C_ON=1'b0;
    defparam \c0.tx.i17744_3_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i17744_3_lut_LC_10_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.tx.i17744_3_lut_LC_10_17_0  (
            .in0(N__28939),
            .in1(N__34161),
            .in2(_gnd_net_),
            .in3(N__34064),
            .lcout(),
            .ltout(\c0.n21331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13772_4_lut_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.i13772_4_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i13772_4_lut_LC_10_17_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.i13772_4_lut_LC_10_17_1  (
            .in0(N__29280),
            .in1(N__27412),
            .in2(N__26347),
            .in3(N__29005),
            .lcout(),
            .ltout(\c0.n17354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_10_17_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_10_17_2  (
            .in0(N__29032),
            .in1(N__26341),
            .in2(N__26344),
            .in3(N__29281),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70994),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17934_2_lut_LC_10_17_4 .C_ON=1'b0;
    defparam \c0.i17934_2_lut_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17934_2_lut_LC_10_17_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i17934_2_lut_LC_10_17_4  (
            .in0(N__29159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27543),
            .lcout(\c0.n21521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_10_17_5 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx.i2_4_lut_LC_10_17_5  (
            .in0(N__26712),
            .in1(N__26667),
            .in2(N__26731),
            .in3(N__26697),
            .lcout(),
            .ltout(\c0.tx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i12488_4_lut_LC_10_17_6 .C_ON=1'b0;
    defparam \c0.tx.i12488_4_lut_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i12488_4_lut_LC_10_17_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx.i12488_4_lut_LC_10_17_6  (
            .in0(N__26682),
            .in1(N__26652),
            .in2(N__26335),
            .in3(N__26637),
            .lcout(\c0.n15938 ),
            .ltout(\c0.n15938_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_4_lut_LC_10_17_7 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_4_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_4_lut_LC_10_17_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \c0.tx.i1_4_lut_4_lut_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__34062),
            .in2(N__26332),
            .in3(N__29158),
            .lcout(\c0.tx.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_10_18_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i0_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_10_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__26329),
            .in2(_gnd_net_),
            .in3(N__26323),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\c0.tx.n17274 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i1_LC_10_18_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i1_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__26730),
            .in2(_gnd_net_),
            .in3(N__26716),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx.n17274 ),
            .carryout(\c0.tx.n17275 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i2_LC_10_18_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i2_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__26713),
            .in2(_gnd_net_),
            .in3(N__26701),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx.n17275 ),
            .carryout(\c0.tx.n17276 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i3_LC_10_18_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i3_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_10_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__26698),
            .in2(_gnd_net_),
            .in3(N__26686),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx.n17276 ),
            .carryout(\c0.tx.n17277 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i4_LC_10_18_4 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i4_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_10_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__26683),
            .in2(_gnd_net_),
            .in3(N__26671),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx.n17277 ),
            .carryout(\c0.tx.n17278 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i5_LC_10_18_5 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i5_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_10_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__26668),
            .in2(_gnd_net_),
            .in3(N__26656),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx.n17278 ),
            .carryout(\c0.tx.n17279 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i6_LC_10_18_6 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i6_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__26653),
            .in2(_gnd_net_),
            .in3(N__26641),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx.n17279 ),
            .carryout(\c0.tx.n17280 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i7_LC_10_18_7 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i7_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_10_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__26638),
            .in2(_gnd_net_),
            .in3(N__26626),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx.n17280 ),
            .carryout(\c0.tx.n17281 ),
            .clk(N__70999),
            .ce(N__29199),
            .sr(N__27651));
    defparam \c0.tx.r_Clock_Count__i8_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__27681),
            .in2(_gnd_net_),
            .in3(N__26623),
            .lcout(\c0.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71004),
            .ce(N__29203),
            .sr(N__27655));
    defparam \c0.FRAME_MATCHER_state_i21_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_10_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_10_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__31506),
            .in2(_gnd_net_),
            .in3(N__40480),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71017),
            .ce(),
            .sr(N__31480));
    defparam \c0.FRAME_MATCHER_state_i6_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_10_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_10_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__29548),
            .in2(_gnd_net_),
            .in3(N__40524),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71027),
            .ce(),
            .sr(N__27568));
    defparam \c0.FRAME_MATCHER_state_i10_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_10_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_10_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__27612),
            .in2(_gnd_net_),
            .in3(N__40525),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71036),
            .ce(),
            .sr(N__26755));
    defparam \c0.FRAME_MATCHER_state_i13_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_10_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_10_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__27770),
            .in2(_gnd_net_),
            .in3(N__40527),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71048),
            .ce(),
            .sr(N__27751));
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_10_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__29591),
            .in2(_gnd_net_),
            .in3(N__40529),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71060),
            .ce(),
            .sr(N__26746));
    defparam \c0.i1_2_lut_adj_485_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_485_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_485_LC_10_26_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_485_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(N__29590),
            .in2(_gnd_net_),
            .in3(N__41476),
            .lcout(\c0.n18617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadB_I_0_79_2_lut_LC_11_4_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadB_I_0_79_2_lut_LC_11_4_0  (
            .in0(N__26815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26780),
            .lcout(b_delay_counter_15__N_2933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_delayed_62_LC_11_4_1 .C_ON=1'b0;
    defparam \quad_counter1.quadB_delayed_62_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadB_delayed_62_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.quadB_delayed_62_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26816),
            .lcout(quadB_delayed_adj_3585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71148),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_LC_11_5_2 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_LC_11_5_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter1.i9_4_lut_LC_11_5_2  (
            .in0(N__28026),
            .in1(N__27867),
            .in2(N__28075),
            .in3(N__27926),
            .lcout(),
            .ltout(\quad_counter1.n25_adj_3577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_LC_11_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_LC_11_5_3  (
            .in0(N__26824),
            .in1(N__26767),
            .in2(N__26734),
            .in3(N__26761),
            .lcout(n11343),
            .ltout(n11343_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_11_5_4.C_ON=1'b0;
    defparam i1_4_lut_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_11_5_4.LUT_INIT=16'b1111111110010000;
    LogicCell40 i1_4_lut_LC_11_5_4 (
            .in0(N__26781),
            .in1(N__26817),
            .in2(N__26830),
            .in3(N__28231),
            .lcout(n12417),
            .ltout(n12417_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i0_LC_11_5_5 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i0_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i0_LC_11_5_5 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \quad_counter1.b_delay_counter__i0_LC_11_5_5  (
            .in0(N__27927),
            .in1(N__28245),
            .in2(N__26827),
            .in3(N__27913),
            .lcout(b_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71132),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_LC_11_5_6 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_LC_11_5_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i12_4_lut_LC_11_5_6  (
            .in0(N__28089),
            .in1(N__28056),
            .in2(N__27886),
            .in3(N__28302),
            .lcout(\quad_counter1.n28_adj_3574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_65_LC_11_5_7 .C_ON=1'b0;
    defparam \quad_counter1.B_65_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_65_LC_11_5_7 .LUT_INIT=16'b1100111011001000;
    LogicCell40 \quad_counter1.B_65_LC_11_5_7  (
            .in0(N__26818),
            .in1(N__29903),
            .in2(N__26791),
            .in3(N__26782),
            .lcout(B_filtered_adj_3582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71132),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_LC_11_6_0 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_LC_11_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_LC_11_6_0  (
            .in0(N__28284),
            .in1(N__28317),
            .in2(N__27904),
            .in3(N__28041),
            .lcout(\quad_counter1.n26_adj_3575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_LC_11_6_7 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_LC_11_6_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_LC_11_6_7  (
            .in0(N__27996),
            .in1(N__28011),
            .in2(N__27982),
            .in3(N__27852),
            .lcout(\quad_counter1.n27_adj_3576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_63_LC_11_7_6 .C_ON=1'b0;
    defparam \quad_counter1.A_63_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_63_LC_11_7_6 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \quad_counter1.A_63_LC_11_7_6  (
            .in0(N__26938),
            .in1(N__28213),
            .in2(N__28174),
            .in3(N__29857),
            .lcout(A_filtered_adj_3581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71102),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_951_LC_11_7_7.C_ON=1'b0;
    defparam i1_3_lut_adj_951_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_951_LC_11_7_7.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_adj_951_LC_11_7_7 (
            .in0(N__28212),
            .in1(N__28170),
            .in2(_gnd_net_),
            .in3(N__26937),
            .lcout(n12477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_LC_11_8_5 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_LC_11_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i3_4_lut_LC_11_8_5  (
            .in0(N__28428),
            .in1(N__28530),
            .in2(N__28597),
            .in3(N__26890),
            .lcout(),
            .ltout(\quad_counter1.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_946_LC_11_8_6 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_946_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_946_LC_11_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_946_LC_11_8_6  (
            .in0(N__28443),
            .in1(N__28398),
            .in2(N__26944),
            .in3(N__26848),
            .lcout(),
            .ltout(\quad_counter1.n24_adj_3578_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_947_LC_11_8_7 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_947_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_947_LC_11_8_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_adj_947_LC_11_8_7  (
            .in0(N__28116),
            .in1(N__28563),
            .in2(N__26941),
            .in3(N__28147),
            .lcout(n11351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i30_LC_11_9_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i30_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i30_LC_11_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i30_LC_11_9_0  (
            .in0(N__36247),
            .in1(N__30638),
            .in2(_gnd_net_),
            .in3(N__30616),
            .lcout(encoder1_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71075),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_LC_11_9_1 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_LC_11_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter0.i3_4_lut_LC_11_9_1  (
            .in0(N__26854),
            .in1(N__26883),
            .in2(N__26929),
            .in3(N__26908),
            .lcout(count_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_LC_11_9_2 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_LC_11_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i2_2_lut_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__28548),
            .in2(_gnd_net_),
            .in3(N__28383),
            .lcout(\quad_counter1.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_delayed_67_LC_11_9_3 .C_ON=1'b0;
    defparam \quad_counter0.A_delayed_67_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_delayed_67_LC_11_9_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \quad_counter0.A_delayed_67_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__26884),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71075),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_945_LC_11_9_7 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_945_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_945_LC_11_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i9_4_lut_adj_945_LC_11_9_7  (
            .in0(N__28578),
            .in1(N__28413),
            .in2(N__28369),
            .in3(N__28332),
            .lcout(\quad_counter1.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i10_LC_11_10_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i10_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i10_LC_11_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i10_LC_11_10_0  (
            .in0(N__35632),
            .in1(N__27128),
            .in2(_gnd_net_),
            .in3(N__26842),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i11_LC_11_10_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i11_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i11_LC_11_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i11_LC_11_10_1  (
            .in0(N__33257),
            .in1(N__35636),
            .in2(_gnd_net_),
            .in3(N__26836),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i12_LC_11_10_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i12_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i12_LC_11_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i12_LC_11_10_2  (
            .in0(N__35633),
            .in1(N__28838),
            .in2(_gnd_net_),
            .in3(N__27028),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i13_LC_11_10_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i13_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i13_LC_11_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i13_LC_11_10_3  (
            .in0(N__28673),
            .in1(N__35637),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i14_LC_11_10_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i14_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i14_LC_11_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i14_LC_11_10_4  (
            .in0(N__35634),
            .in1(N__27245),
            .in2(_gnd_net_),
            .in3(N__27016),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i15_LC_11_10_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i15_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i15_LC_11_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i15_LC_11_10_5  (
            .in0(N__26996),
            .in1(N__35638),
            .in2(_gnd_net_),
            .in3(N__27010),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i16_LC_11_10_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i16_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i16_LC_11_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i16_LC_11_10_6  (
            .in0(N__35635),
            .in1(N__27269),
            .in2(_gnd_net_),
            .in3(N__26974),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i17_LC_11_10_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i17_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i17_LC_11_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i17_LC_11_10_7  (
            .in0(N__28725),
            .in1(N__35639),
            .in2(_gnd_net_),
            .in3(N__26968),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71061),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i18_LC_11_11_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i18_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i18_LC_11_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i18_LC_11_11_1  (
            .in0(N__33290),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(N__30427),
            .lcout(encoder1_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__3__5387_LC_11_11_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__3__5387_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__3__5387_LC_11_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_6__3__5387_LC_11_11_3  (
            .in0(N__35548),
            .in1(N__35499),
            .in2(_gnd_net_),
            .in3(N__46934),
            .lcout(data_out_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__4__5386_LC_11_11_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__4__5386_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__4__5386_LC_11_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_6__4__5386_LC_11_11_4  (
            .in0(N__46931),
            .in1(N__27298),
            .in2(_gnd_net_),
            .in3(N__26958),
            .lcout(data_out_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__1__5389_LC_11_11_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__1__5389_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__1__5389_LC_11_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_6__1__5389_LC_11_11_5  (
            .in0(N__27345),
            .in1(N__27154),
            .in2(_gnd_net_),
            .in3(N__46933),
            .lcout(data_out_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__2__5372_LC_11_11_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__2__5372_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__2__5372_LC_11_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__2__5372_LC_11_11_6  (
            .in0(N__46932),
            .in1(N__27129),
            .in2(_gnd_net_),
            .in3(N__28459),
            .lcout(data_out_frame_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__4__5378_LC_11_11_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__4__5378_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__4__5378_LC_11_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__4__5378_LC_11_11_7  (
            .in0(N__27109),
            .in1(N__27081),
            .in2(_gnd_net_),
            .in3(N__46935),
            .lcout(data_out_frame_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71049),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i26_LC_11_12_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i26_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i26_LC_11_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i26_LC_11_12_0  (
            .in0(N__35728),
            .in1(N__35891),
            .in2(_gnd_net_),
            .in3(N__27067),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i4_LC_11_12_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i4_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i4_LC_11_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i4_LC_11_12_1  (
            .in0(N__30908),
            .in1(N__36258),
            .in2(_gnd_net_),
            .in3(N__30055),
            .lcout(encoder1_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i19_LC_11_12_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i19_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i19_LC_11_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i19_LC_11_12_2  (
            .in0(N__36256),
            .in1(N__30407),
            .in2(_gnd_net_),
            .in3(N__30388),
            .lcout(encoder1_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i30_LC_11_12_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i30_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i30_LC_11_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i30_LC_11_12_4  (
            .in0(N__35729),
            .in1(N__27047),
            .in2(_gnd_net_),
            .in3(N__27061),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17712_4_lut_LC_11_12_5 .C_ON=1'b0;
    defparam \c0.i17712_4_lut_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17712_4_lut_LC_11_12_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \c0.i17712_4_lut_LC_11_12_5  (
            .in0(N__33307),
            .in1(N__32749),
            .in2(N__36986),
            .in3(N__40919),
            .lcout(\c0.n21299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i7_LC_11_12_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i7_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i7_LC_11_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i7_LC_11_12_6  (
            .in0(N__36257),
            .in1(N__29978),
            .in2(_gnd_net_),
            .in3(N__29959),
            .lcout(encoder1_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i8_LC_11_12_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i8_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i8_LC_11_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i8_LC_11_12_7  (
            .in0(N__36356),
            .in1(N__36259),
            .in2(_gnd_net_),
            .in3(N__29944),
            .lcout(encoder1_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71037),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_11_13_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_11_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_11_13_0  (
            .in0(N__28704),
            .in1(N__27346),
            .in2(_gnd_net_),
            .in3(N__40905),
            .lcout(\c0.n5_adj_3102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__1__5365_LC_11_13_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__1__5365_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__1__5365_LC_11_13_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_9__1__5365_LC_11_13_1  (
            .in0(N__27331),
            .in1(N__31242),
            .in2(_gnd_net_),
            .in3(N__46736),
            .lcout(data_out_frame_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71028),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i28_LC_11_13_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i28_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i28_LC_11_13_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i28_LC_11_13_2  (
            .in0(N__27293),
            .in1(N__35688),
            .in2(_gnd_net_),
            .in3(N__27304),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71028),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__0__5382_LC_11_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__0__5382_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__0__5382_LC_11_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__0__5382_LC_11_13_3  (
            .in0(N__27274),
            .in1(N__33321),
            .in2(_gnd_net_),
            .in3(N__46735),
            .lcout(\c0.data_out_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71028),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__6__5368_LC_11_13_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__6__5368_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__6__5368_LC_11_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__6__5368_LC_11_13_4  (
            .in0(N__46733),
            .in1(N__27250),
            .in2(_gnd_net_),
            .in3(N__27225),
            .lcout(data_out_frame_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71028),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__4__5362_LC_11_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__4__5362_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__4__5362_LC_11_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_9__4__5362_LC_11_13_6  (
            .in0(N__46734),
            .in1(N__27207),
            .in2(_gnd_net_),
            .in3(N__30828),
            .lcout(data_out_frame_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71028),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17982_4_lut_LC_11_14_0 .C_ON=1'b0;
    defparam \c0.i17982_4_lut_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17982_4_lut_LC_11_14_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.i17982_4_lut_LC_11_14_0  (
            .in0(N__36765),
            .in1(N__36952),
            .in2(N__27367),
            .in3(N__27184),
            .lcout(\c0.n21570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17714_4_lut_LC_11_14_2 .C_ON=1'b0;
    defparam \c0.i17714_4_lut_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17714_4_lut_LC_11_14_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.i17714_4_lut_LC_11_14_2  (
            .in0(N__29071),
            .in1(N__28693),
            .in2(N__37465),
            .in3(N__27178),
            .lcout(\c0.n21301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21623_bdd_4_lut_LC_11_14_3 .C_ON=1'b0;
    defparam \c0.n21623_bdd_4_lut_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.n21623_bdd_4_lut_LC_11_14_3 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n21623_bdd_4_lut_LC_11_14_3  (
            .in0(N__27375),
            .in1(N__33217),
            .in2(N__36766),
            .in3(N__27169),
            .lcout(),
            .ltout(\c0.n21626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17984_4_lut_LC_11_14_4 .C_ON=1'b0;
    defparam \c0.i17984_4_lut_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17984_4_lut_LC_11_14_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i17984_4_lut_LC_11_14_4  (
            .in0(N__36764),
            .in1(N__27358),
            .in2(N__27406),
            .in3(N__36951),
            .lcout(\c0.n21572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__7__5359_LC_11_14_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__7__5359_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__7__5359_LC_11_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_9__7__5359_LC_11_14_5  (
            .in0(N__27376),
            .in1(N__27402),
            .in2(_gnd_net_),
            .in3(N__46930),
            .lcout(data_out_frame_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71018),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__3__5347_LC_11_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__3__5347_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__3__5347_LC_11_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_11__3__5347_LC_11_14_6  (
            .in0(N__46929),
            .in1(N__30411),
            .in2(_gnd_net_),
            .in3(N__28869),
            .lcout(data_out_frame_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71018),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_11_15_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_11_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_11_15_0  (
            .in0(N__40855),
            .in1(N__28815),
            .in2(_gnd_net_),
            .in3(N__28741),
            .lcout(\c0.n11_adj_3472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_15_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_15_1  (
            .in0(N__28960),
            .in1(N__28881),
            .in2(_gnd_net_),
            .in3(N__40853),
            .lcout(\c0.n11_adj_3479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_11_15_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_11_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_11_15_3  (
            .in0(N__30889),
            .in1(N__37027),
            .in2(_gnd_net_),
            .in3(N__40854),
            .lcout(),
            .ltout(\c0.n11_adj_3444_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17702_4_lut_LC_11_15_4 .C_ON=1'b0;
    defparam \c0.i17702_4_lut_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17702_4_lut_LC_11_15_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.i17702_4_lut_LC_11_15_4  (
            .in0(N__36930),
            .in1(N__36702),
            .in2(N__27352),
            .in3(N__27460),
            .lcout(),
            .ltout(\c0.n21289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17989_4_lut_LC_11_15_5 .C_ON=1'b0;
    defparam \c0.i17989_4_lut_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17989_4_lut_LC_11_15_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.i17989_4_lut_LC_11_15_5  (
            .in0(N__36703),
            .in1(N__30802),
            .in2(N__27349),
            .in3(N__36931),
            .lcout(\c0.n21577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_220_LC_11_15_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_220_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_220_LC_11_15_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_220_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__29144),
            .in2(_gnd_net_),
            .in3(N__30955),
            .lcout(n6866),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_11_16_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_651_LC_11_16_1 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_651_LC_11_16_1  (
            .in0(N__27687),
            .in1(N__34063),
            .in2(_gnd_net_),
            .in3(N__27514),
            .lcout(\c0.n55 ),
            .ltout(\c0.n55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_11_16_2 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_11_16_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \c0.tx.i1_2_lut_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27490),
            .in3(N__29143),
            .lcout(),
            .ltout(\c0.n14301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_11_16_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_11_16_3 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_11_16_3  (
            .in0(N__29284),
            .in1(N__27484),
            .in2(N__27487),
            .in3(N__34085),
            .lcout(r_SM_Main_1_adj_3592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71005),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12492_2_lut_3_lut_LC_11_16_4 .C_ON=1'b0;
    defparam \c0.i12492_2_lut_3_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12492_2_lut_3_lut_LC_11_16_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i12492_2_lut_3_lut_LC_11_16_4  (
            .in0(N__27515),
            .in1(N__29142),
            .in2(_gnd_net_),
            .in3(N__27688),
            .lcout(\c0.n15942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_11_16_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_11_16_5 .LUT_INIT=16'b0101010011110000;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_11_16_5  (
            .in0(N__29283),
            .in1(N__27478),
            .in2(N__31295),
            .in3(N__29233),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71005),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17701_3_lut_LC_11_16_6 .C_ON=1'b0;
    defparam \c0.i17701_3_lut_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17701_3_lut_LC_11_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i17701_3_lut_LC_11_16_6  (
            .in0(N__28768),
            .in1(N__27471),
            .in2(_gnd_net_),
            .in3(N__40856),
            .lcout(\c0.n21288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i6_LC_11_16_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i6_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i6_LC_11_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i6_LC_11_16_7  (
            .in0(N__35687),
            .in1(N__27431),
            .in2(_gnd_net_),
            .in3(N__27454),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71005),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17930_3_lut_LC_11_17_0 .C_ON=1'b0;
    defparam \c0.i17930_3_lut_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17930_3_lut_LC_11_17_0 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \c0.i17930_3_lut_LC_11_17_0  (
            .in0(N__34060),
            .in1(N__29162),
            .in2(_gnd_net_),
            .in3(N__29056),
            .lcout(\c0.n21517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_LC_11_17_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.tx.i2_3_lut_LC_11_17_1  (
            .in0(N__29269),
            .in1(N__34059),
            .in2(_gnd_net_),
            .in3(N__27516),
            .lcout(\c0.tx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17919_2_lut_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.i17919_2_lut_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17919_2_lut_LC_11_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i17919_2_lut_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__34226),
            .in2(_gnd_net_),
            .in3(N__29057),
            .lcout(),
            .ltout(\c0.n21506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_11_17_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_11_17_3 .LUT_INIT=16'b0010100011001100;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_11_17_3  (
            .in0(N__29272),
            .in1(N__27542),
            .in2(N__27559),
            .in3(N__28988),
            .lcout(\c0.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70997),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17898_4_lut_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.i17898_4_lut_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17898_4_lut_LC_11_17_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i17898_4_lut_LC_11_17_4  (
            .in0(N__34228),
            .in1(N__27555),
            .in2(N__27544),
            .in3(N__29055),
            .lcout(),
            .ltout(\c0.n21414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_4_lut_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.i25_4_lut_4_lut_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_4_lut_LC_11_17_5 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.i25_4_lut_4_lut_LC_11_17_5  (
            .in0(N__29270),
            .in1(N__30943),
            .in2(N__27526),
            .in3(N__34061),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_11_17_6 .LUT_INIT=16'b0110110000001100;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_11_17_6  (
            .in0(N__34229),
            .in1(N__29058),
            .in2(N__28993),
            .in3(N__29271),
            .lcout(\c0.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__70997),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21611_bdd_4_lut_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.n21611_bdd_4_lut_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.n21611_bdd_4_lut_LC_11_17_7 .LUT_INIT=16'b1100111011000010;
    LogicCell40 \c0.n21611_bdd_4_lut_LC_11_17_7  (
            .in0(N__31186),
            .in1(N__33991),
            .in2(N__34233),
            .in3(N__28945),
            .lcout(\c0.n21614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_5164_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.tx_transmit_5164_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_5164_LC_11_18_0 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \c0.tx_transmit_5164_LC_11_18_0  (
            .in0(N__39492),
            .in1(N__39071),
            .in2(N__38985),
            .in3(N__31519),
            .lcout(\c0.r_SM_Main_2_N_2547_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71006),
            .ce(),
            .sr(N__31447));
    defparam \c0.i12472_2_lut_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.i12472_2_lut_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12472_2_lut_LC_11_18_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i12472_2_lut_LC_11_18_2  (
            .in0(N__27517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27678),
            .lcout(\c0.n15920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_4_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_4_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_4_lut_LC_11_18_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i2_2_lut_4_lut_LC_11_18_4  (
            .in0(N__29161),
            .in1(N__34096),
            .in2(N__30952),
            .in3(N__29303),
            .lcout(n9377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_adj_219_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_adj_219_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_adj_219_LC_11_18_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.tx.i2_3_lut_adj_219_LC_11_18_5  (
            .in0(N__27679),
            .in1(N__29160),
            .in2(_gnd_net_),
            .in3(N__27496),
            .lcout(),
            .ltout(\c0.tx.n21179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i18012_4_lut_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.tx.i18012_4_lut_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i18012_4_lut_LC_11_18_6 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \c0.tx.i18012_4_lut_LC_11_18_6  (
            .in0(N__27697),
            .in1(N__34097),
            .in2(N__27691),
            .in3(N__27680),
            .lcout(\c0.tx.n12759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i26_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_11_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_11_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__27798),
            .in2(_gnd_net_),
            .in3(N__40533),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71011),
            .ce(),
            .sr(N__27784));
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_11_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__40543),
            .in2(_gnd_net_),
            .in3(N__27737),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71019),
            .ce(),
            .sr(N__27838));
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_11_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__29356),
            .in2(_gnd_net_),
            .in3(N__40443),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71029),
            .ce(),
            .sr(N__29083));
    defparam \c0.i4_4_lut_adj_688_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_688_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_688_LC_11_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_688_LC_11_22_0  (
            .in0(N__27771),
            .in1(N__27634),
            .in2(N__27613),
            .in3(N__27590),
            .lcout(\c0.n10_adj_3488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i11_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_11_22_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_11_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__27592),
            .in2(_gnd_net_),
            .in3(N__40522),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71038),
            .ce(),
            .sr(N__27580));
    defparam \c0.i1_2_lut_adj_267_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_267_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_267_LC_11_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_267_LC_11_22_3  (
            .in0(N__27591),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41456),
            .lcout(\c0.n18669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_268_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_268_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_268_LC_11_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_268_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__27718),
            .in2(_gnd_net_),
            .in3(N__41457),
            .lcout(\c0.n18651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_269_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_269_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_269_LC_11_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_269_LC_11_22_6  (
            .in0(N__41458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29553),
            .lcout(\c0.n18679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_363_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_363_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_363_LC_11_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_363_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__27739),
            .in2(_gnd_net_),
            .in3(N__41459),
            .lcout(\c0.n18637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_686_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_686_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_686_LC_11_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_686_LC_11_23_0  (
            .in0(N__27804),
            .in1(N__31502),
            .in2(N__29500),
            .in3(N__27824),
            .lcout(\c0.n10_adj_3438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_11_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_11_23_1  (
            .in0(N__27826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40523),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71050),
            .ce(),
            .sr(N__27814));
    defparam \c0.i1_2_lut_adj_346_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_346_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_346_LC_11_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_346_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__27825),
            .in2(_gnd_net_),
            .in3(N__41462),
            .lcout(\c0.n18635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_370_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_370_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_370_LC_11_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_370_LC_11_23_4  (
            .in0(N__27805),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41463),
            .lcout(\c0.n18623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_260_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_260_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_260_LC_11_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_260_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__27772),
            .in2(_gnd_net_),
            .in3(N__41460),
            .lcout(\c0.n18665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_263_LC_11_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_263_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_263_LC_11_23_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_263_LC_11_23_7  (
            .in0(N__41461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29797),
            .lcout(\c0.n18641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_677_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_677_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_677_LC_11_24_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_677_LC_11_24_0  (
            .in0(N__34932),
            .in1(N__27738),
            .in2(N__31666),
            .in3(N__27710),
            .lcout(\c0.n16_adj_3484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i20_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_11_24_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_11_24_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_11_24_1  (
            .in0(N__40526),
            .in1(_gnd_net_),
            .in2(N__27717),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71062),
            .ce(),
            .sr(N__27964));
    defparam \c0.i1_2_lut_adj_366_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_366_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_366_LC_11_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_366_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__29775),
            .in2(_gnd_net_),
            .in3(N__41464),
            .lcout(\c0.n18625 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_851_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_851_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_851_LC_11_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_851_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__29735),
            .in2(_gnd_net_),
            .in3(N__41465),
            .lcout(\c0.n18677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i19_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_11_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_11_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_11_25_0  (
            .in0(N__40528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29796),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71074),
            .ce(),
            .sr(N__27940));
    defparam \c0.FRAME_MATCHER_state_i3_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_11_26_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_11_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__29452),
            .in2(_gnd_net_),
            .in3(N__40553),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71087),
            .ce(),
            .sr(N__29437));
    defparam \quad_counter1.add_86_2_lut_LC_12_5_0 .C_ON=1'b1;
    defparam \quad_counter1.add_86_2_lut_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_86_2_lut_LC_12_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_86_2_lut_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__27928),
            .in2(_gnd_net_),
            .in3(N__27907),
            .lcout(n187),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\quad_counter1.n17237 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i1_LC_12_5_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i1_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i1_LC_12_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i1_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__27903),
            .in2(_gnd_net_),
            .in3(N__27889),
            .lcout(\quad_counter1.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n17237 ),
            .carryout(\quad_counter1.n17238 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i2_LC_12_5_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i2_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i2_LC_12_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i2_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__27885),
            .in2(_gnd_net_),
            .in3(N__27871),
            .lcout(\quad_counter1.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n17238 ),
            .carryout(\quad_counter1.n17239 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i3_LC_12_5_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i3_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i3_LC_12_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i3_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__27868),
            .in2(_gnd_net_),
            .in3(N__27856),
            .lcout(\quad_counter1.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n17239 ),
            .carryout(\quad_counter1.n17240 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i4_LC_12_5_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i4_LC_12_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i4_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__27853),
            .in2(_gnd_net_),
            .in3(N__27841),
            .lcout(\quad_counter1.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n17240 ),
            .carryout(\quad_counter1.n17241 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i5_LC_12_5_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i5_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i5_LC_12_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i5_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__28090),
            .in2(_gnd_net_),
            .in3(N__28078),
            .lcout(\quad_counter1.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n17241 ),
            .carryout(\quad_counter1.n17242 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i6_LC_12_5_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i6_LC_12_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i6_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__28074),
            .in2(_gnd_net_),
            .in3(N__28060),
            .lcout(\quad_counter1.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n17242 ),
            .carryout(\quad_counter1.n17243 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i7_LC_12_5_7 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i7_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i7_LC_12_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i7_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__28057),
            .in2(_gnd_net_),
            .in3(N__28045),
            .lcout(\quad_counter1.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n17243 ),
            .carryout(\quad_counter1.n17244 ),
            .clk(N__71149),
            .ce(N__28273),
            .sr(N__28244));
    defparam \quad_counter1.b_delay_counter__i8_LC_12_6_0 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i8_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i8_LC_12_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i8_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__28042),
            .in2(_gnd_net_),
            .in3(N__28030),
            .lcout(\quad_counter1.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\quad_counter1.n17245 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i9_LC_12_6_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i9_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i9_LC_12_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i9_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__28027),
            .in2(_gnd_net_),
            .in3(N__28015),
            .lcout(\quad_counter1.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n17245 ),
            .carryout(\quad_counter1.n17246 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i10_LC_12_6_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i10_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i10_LC_12_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i10_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__28012),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(\quad_counter1.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n17246 ),
            .carryout(\quad_counter1.n17247 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i11_LC_12_6_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i11_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i11_LC_12_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i11_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__27997),
            .in2(_gnd_net_),
            .in3(N__27985),
            .lcout(\quad_counter1.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n17247 ),
            .carryout(\quad_counter1.n17248 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i12_LC_12_6_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i12_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i12_LC_12_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i12_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__27981),
            .in2(_gnd_net_),
            .in3(N__27967),
            .lcout(\quad_counter1.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n17248 ),
            .carryout(\quad_counter1.n17249 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i13_LC_12_6_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i13_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i13_LC_12_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i13_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__28318),
            .in2(_gnd_net_),
            .in3(N__28306),
            .lcout(\quad_counter1.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n17249 ),
            .carryout(\quad_counter1.n17250 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i14_LC_12_6_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i14_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i14_LC_12_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i14_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__28303),
            .in2(_gnd_net_),
            .in3(N__28291),
            .lcout(\quad_counter1.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n17250 ),
            .carryout(\quad_counter1.n17251 ),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.b_delay_counter__i15_LC_12_6_7 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i15_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i15_LC_12_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i15_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__28285),
            .in2(_gnd_net_),
            .in3(N__28288),
            .lcout(\quad_counter1.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71134),
            .ce(N__28266),
            .sr(N__28246));
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_12_7_0 .C_ON=1'b0;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadA_I_0_73_2_lut_LC_12_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter1.quadA_I_0_73_2_lut_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__28205),
            .in2(_gnd_net_),
            .in3(N__28169),
            .lcout(a_delay_counter_15__N_2916_adj_3589),
            .ltout(a_delay_counter_15__N_2916_adj_3589_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i0_LC_12_7_1 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i0_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i0_LC_12_7_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \quad_counter1.a_delay_counter__i0_LC_12_7_1  (
            .in0(N__28126),
            .in1(N__28140),
            .in2(N__28150),
            .in3(N__28508),
            .lcout(a_delay_counter_0_adj_3583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71118),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i7_3_lut_LC_12_7_3 .C_ON=1'b0;
    defparam \quad_counter1.i7_3_lut_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i7_3_lut_LC_12_7_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \quad_counter1.i7_3_lut_LC_12_7_3  (
            .in0(N__28351),
            .in1(N__28139),
            .in2(_gnd_net_),
            .in3(N__28101),
            .lcout(\quad_counter1.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_85_2_lut_LC_12_8_0 .C_ON=1'b1;
    defparam \quad_counter1.add_85_2_lut_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_85_2_lut_LC_12_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_85_2_lut_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__28141),
            .in2(_gnd_net_),
            .in3(N__28120),
            .lcout(n39_adj_3587),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\quad_counter1.n17252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i1_LC_12_8_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i1_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i1_LC_12_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__28117),
            .in2(_gnd_net_),
            .in3(N__28105),
            .lcout(\quad_counter1.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n17252 ),
            .carryout(\quad_counter1.n17253 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i2_LC_12_8_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i2_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i2_LC_12_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i2_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__28102),
            .in2(_gnd_net_),
            .in3(N__28447),
            .lcout(\quad_counter1.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n17253 ),
            .carryout(\quad_counter1.n17254 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i3_LC_12_8_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i3_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i3_LC_12_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i3_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__28444),
            .in2(_gnd_net_),
            .in3(N__28432),
            .lcout(\quad_counter1.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n17254 ),
            .carryout(\quad_counter1.n17255 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i4_LC_12_8_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i4_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i4_LC_12_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i4_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__28429),
            .in2(_gnd_net_),
            .in3(N__28417),
            .lcout(\quad_counter1.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n17255 ),
            .carryout(\quad_counter1.n17256 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i5_LC_12_8_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i5_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i5_LC_12_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i5_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__28414),
            .in2(_gnd_net_),
            .in3(N__28402),
            .lcout(\quad_counter1.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n17256 ),
            .carryout(\quad_counter1.n17257 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i6_LC_12_8_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i6_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i6_LC_12_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i6_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__28399),
            .in2(_gnd_net_),
            .in3(N__28387),
            .lcout(\quad_counter1.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n17257 ),
            .carryout(\quad_counter1.n17258 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i7_LC_12_8_7 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i7_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i7_LC_12_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i7_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__28384),
            .in2(_gnd_net_),
            .in3(N__28372),
            .lcout(\quad_counter1.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n17258 ),
            .carryout(\quad_counter1.n17259 ),
            .clk(N__71104),
            .ce(N__28515),
            .sr(N__28491));
    defparam \quad_counter1.a_delay_counter__i8_LC_12_9_0 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i8_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i8_LC_12_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i8_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__28368),
            .in2(_gnd_net_),
            .in3(N__28354),
            .lcout(\quad_counter1.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\quad_counter1.n17260 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i9_LC_12_9_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i9_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i9_LC_12_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i9_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__28350),
            .in2(_gnd_net_),
            .in3(N__28336),
            .lcout(\quad_counter1.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n17260 ),
            .carryout(\quad_counter1.n17261 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i10_LC_12_9_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i10_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i10_LC_12_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i10_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__28333),
            .in2(_gnd_net_),
            .in3(N__28321),
            .lcout(\quad_counter1.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n17261 ),
            .carryout(\quad_counter1.n17262 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i11_LC_12_9_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i11_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i11_LC_12_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i11_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__28596),
            .in2(_gnd_net_),
            .in3(N__28582),
            .lcout(\quad_counter1.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n17262 ),
            .carryout(\quad_counter1.n17263 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i12_LC_12_9_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i12_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i12_LC_12_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i12_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__28579),
            .in2(_gnd_net_),
            .in3(N__28567),
            .lcout(\quad_counter1.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n17263 ),
            .carryout(\quad_counter1.n17264 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i13_LC_12_9_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i13_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i13_LC_12_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i13_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__28564),
            .in2(_gnd_net_),
            .in3(N__28552),
            .lcout(\quad_counter1.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n17264 ),
            .carryout(\quad_counter1.n17265 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i14_LC_12_9_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i14_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i14_LC_12_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i14_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__28549),
            .in2(_gnd_net_),
            .in3(N__28537),
            .lcout(\quad_counter1.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n17265 ),
            .carryout(\quad_counter1.n17266 ),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.a_delay_counter__i15_LC_12_9_7 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i15_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i15_LC_12_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i15_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__28531),
            .in2(_gnd_net_),
            .in3(N__28534),
            .lcout(\quad_counter1.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71088),
            .ce(N__28519),
            .sr(N__28492));
    defparam \quad_counter1.count_i0_i9_LC_12_10_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i9_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i9_LC_12_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i9_LC_12_10_0  (
            .in0(N__36177),
            .in1(N__31163),
            .in2(_gnd_net_),
            .in3(N__29929),
            .lcout(encoder1_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i10_LC_12_10_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i10_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i10_LC_12_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i10_LC_12_10_1  (
            .in0(N__30287),
            .in1(N__36178),
            .in2(_gnd_net_),
            .in3(N__30268),
            .lcout(encoder1_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i11_LC_12_10_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i11_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i11_LC_12_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i11_LC_12_10_2  (
            .in0(N__36174),
            .in1(N__30251),
            .in2(_gnd_net_),
            .in3(N__30232),
            .lcout(encoder1_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21647_bdd_4_lut_LC_12_10_3 .C_ON=1'b0;
    defparam \c0.n21647_bdd_4_lut_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.n21647_bdd_4_lut_LC_12_10_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n21647_bdd_4_lut_LC_12_10_3  (
            .in0(N__28474),
            .in1(N__36756),
            .in2(N__32824),
            .in3(N__28458),
            .lcout(\c0.n21650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i13_LC_12_10_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i13_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i13_LC_12_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i13_LC_12_10_4  (
            .in0(N__36175),
            .in1(N__30218),
            .in2(_gnd_net_),
            .in3(N__30196),
            .lcout(encoder1_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i14_LC_12_10_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i14_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i14_LC_12_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i14_LC_12_10_5  (
            .in0(N__30185),
            .in1(N__36179),
            .in2(_gnd_net_),
            .in3(N__30163),
            .lcout(encoder1_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i15_LC_12_10_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i15_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i15_LC_12_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i15_LC_12_10_6  (
            .in0(N__36176),
            .in1(N__30149),
            .in2(_gnd_net_),
            .in3(N__30130),
            .lcout(encoder1_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i16_LC_12_10_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i16_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i16_LC_12_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i16_LC_12_10_7  (
            .in0(N__30116),
            .in1(N__36180),
            .in2(_gnd_net_),
            .in3(N__30094),
            .lcout(encoder1_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71076),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17976_4_lut_LC_12_11_2 .C_ON=1'b0;
    defparam \c0.i17976_4_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17976_4_lut_LC_12_11_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.i17976_4_lut_LC_12_11_2  (
            .in0(N__36954),
            .in1(N__28618),
            .in2(N__36760),
            .in3(N__31006),
            .lcout(),
            .ltout(\c0.n21564_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_4_lut_adj_607_LC_12_11_3 .C_ON=1'b0;
    defparam \c0.i24_3_lut_4_lut_adj_607_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_4_lut_adj_607_LC_12_11_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \c0.i24_3_lut_4_lut_adj_607_LC_12_11_3  (
            .in0(N__37336),
            .in1(N__37450),
            .in2(N__28612),
            .in3(N__35779),
            .lcout(n10_adj_3593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i20_LC_12_11_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i20_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i20_LC_12_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i20_LC_12_11_4  (
            .in0(N__30368),
            .in1(N__36246),
            .in2(_gnd_net_),
            .in3(N__30349),
            .lcout(encoder1_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71063),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i9_LC_12_11_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i9_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i9_LC_12_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i9_LC_12_11_5  (
            .in0(N__30782),
            .in1(N__35730),
            .in2(_gnd_net_),
            .in3(N__28609),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71063),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i22_LC_12_11_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i22_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i22_LC_12_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i22_LC_12_11_7  (
            .in0(N__36245),
            .in1(N__30335),
            .in2(_gnd_net_),
            .in3(N__30316),
            .lcout(encoder1_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71063),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i17_LC_12_12_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i17_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i17_LC_12_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i17_LC_12_12_0  (
            .in0(N__31052),
            .in1(N__36224),
            .in2(_gnd_net_),
            .in3(N__30085),
            .lcout(encoder1_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i29_LC_12_12_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i29_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i29_LC_12_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i29_LC_12_12_1  (
            .in0(N__33350),
            .in1(N__35724),
            .in2(_gnd_net_),
            .in3(N__28687),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i24_LC_12_12_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i24_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i24_LC_12_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \quad_counter1.count_i0_i24_LC_12_12_2  (
            .in0(N__36221),
            .in1(_gnd_net_),
            .in2(N__30762),
            .in3(N__30304),
            .lcout(encoder1_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__5__5337_LC_12_12_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__5__5337_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__5__5337_LC_12_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_12__5__5337_LC_12_12_3  (
            .in0(N__30220),
            .in1(N__30439),
            .in2(_gnd_net_),
            .in3(N__46732),
            .lcout(data_out_frame_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i26_LC_12_12_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i26_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i26_LC_12_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i26_LC_12_12_4  (
            .in0(N__36222),
            .in1(N__32799),
            .in2(_gnd_net_),
            .in3(N__30694),
            .lcout(encoder1_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i27_LC_12_12_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i27_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i27_LC_12_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i27_LC_12_12_5  (
            .in0(N__30661),
            .in1(N__36223),
            .in2(_gnd_net_),
            .in3(N__30680),
            .lcout(encoder1_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__5__5369_LC_12_12_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__5__5369_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__5__5369_LC_12_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__5__5369_LC_12_12_6  (
            .in0(N__46730),
            .in1(N__28678),
            .in2(_gnd_net_),
            .in3(N__33126),
            .lcout(data_out_frame_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__6__5344_LC_12_12_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__6__5344_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__6__5344_LC_12_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_11__6__5344_LC_12_12_7  (
            .in0(N__30336),
            .in1(N__28644),
            .in2(_gnd_net_),
            .in3(N__46731),
            .lcout(data_out_frame_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71051),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i8_LC_12_13_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i8_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i8_LC_12_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i8_LC_12_13_0  (
            .in0(N__28630),
            .in1(N__35723),
            .in2(_gnd_net_),
            .in3(N__30714),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i2_LC_12_13_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i2_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i2_LC_12_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i2_LC_12_13_1  (
            .in0(N__36260),
            .in1(N__31079),
            .in2(_gnd_net_),
            .in3(N__30073),
            .lcout(encoder1_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__4__5346_LC_12_13_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__4__5346_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__4__5346_LC_12_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_11__4__5346_LC_12_13_2  (
            .in0(N__30373),
            .in1(N__28767),
            .in2(_gnd_net_),
            .in3(N__46726),
            .lcout(data_out_frame_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_12_13_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_12_13_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_12_13_3  (
            .in0(N__36475),
            .in1(N__36939),
            .in2(N__28753),
            .in3(N__36698),
            .lcout(\c0.n21653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__6__5336_LC_12_13_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__6__5336_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__6__5336_LC_12_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_12__6__5336_LC_12_13_4  (
            .in0(N__30187),
            .in1(N__28740),
            .in2(_gnd_net_),
            .in3(N__46727),
            .lcout(data_out_frame_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i6_LC_12_13_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i6_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i6_LC_12_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i6_LC_12_13_5  (
            .in0(N__36261),
            .in1(N__30029),
            .in2(_gnd_net_),
            .in3(N__30007),
            .lcout(encoder1_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__1__5381_LC_12_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__1__5381_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__1__5381_LC_12_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__1__5381_LC_12_13_6  (
            .in0(N__28726),
            .in1(N__28705),
            .in2(_gnd_net_),
            .in3(N__46728),
            .lcout(data_out_frame_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71039),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_475_LC_12_13_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_475_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_475_LC_12_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i2_2_lut_adj_475_LC_12_13_7  (
            .in0(N__40975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36940),
            .lcout(\c0.n6_adj_3324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__2__5340_LC_12_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__2__5340_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__2__5340_LC_12_14_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame_12__2__5340_LC_12_14_0  (
            .in0(N__30292),
            .in1(N__46923),
            .in2(_gnd_net_),
            .in3(N__31018),
            .lcout(data_out_frame_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71030),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__3__5331_LC_12_14_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__3__5331_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__3__5331_LC_12_14_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame_13__3__5331_LC_12_14_1  (
            .in0(N__46920),
            .in1(_gnd_net_),
            .in2(N__28894),
            .in3(N__33036),
            .lcout(data_out_frame_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71030),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__3__5355_LC_12_14_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__3__5355_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__3__5355_LC_12_14_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame_10__3__5355_LC_12_14_2  (
            .in0(N__30685),
            .in1(N__46922),
            .in2(_gnd_net_),
            .in3(N__28855),
            .lcout(data_out_frame_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71030),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_12_14_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_12_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_12_14_4  (
            .in0(N__40881),
            .in1(N__28890),
            .in2(_gnd_net_),
            .in3(N__28909),
            .lcout(\c0.n11_adj_3404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__7__5335_LC_12_14_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__7__5335_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__7__5335_LC_12_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_12__7__5335_LC_12_14_5  (
            .in0(N__46919),
            .in1(N__30154),
            .in2(_gnd_net_),
            .in3(N__28882),
            .lcout(data_out_frame_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71030),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18054_LC_12_14_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18054_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18054_LC_12_14_6 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18054_LC_12_14_6  (
            .in0(N__40880),
            .in1(N__36746),
            .in2(N__28870),
            .in3(N__28854),
            .lcout(\c0.n21641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__4__5370_LC_12_14_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__4__5370_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__4__5370_LC_12_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__4__5370_LC_12_14_7  (
            .in0(N__46921),
            .in1(N__28846),
            .in2(_gnd_net_),
            .in3(N__30814),
            .lcout(data_out_frame_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71030),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__6__5328_LC_12_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__6__5328_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__6__5328_LC_12_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_13__6__5328_LC_12_15_1  (
            .in0(N__30033),
            .in1(N__28816),
            .in2(_gnd_net_),
            .in3(N__46737),
            .lcout(data_out_frame_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71020),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_3_lut_4_lut_adj_609_LC_12_15_2 .C_ON=1'b0;
    defparam \c0.i21_3_lut_4_lut_adj_609_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_3_lut_4_lut_adj_609_LC_12_15_2 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.i21_3_lut_4_lut_adj_609_LC_12_15_2  (
            .in0(N__28804),
            .in1(N__33556),
            .in2(N__37451),
            .in3(N__37341),
            .lcout(\c0.n7_adj_3333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21653_bdd_4_lut_4_lut_LC_12_15_3 .C_ON=1'b0;
    defparam \c0.n21653_bdd_4_lut_4_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.n21653_bdd_4_lut_4_lut_LC_12_15_3 .LUT_INIT=16'b1100110010011000;
    LogicCell40 \c0.n21653_bdd_4_lut_4_lut_LC_12_15_3  (
            .in0(N__40824),
            .in1(N__28798),
            .in2(N__30736),
            .in3(N__36908),
            .lcout(n21656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17720_4_lut_LC_12_15_4 .C_ON=1'b0;
    defparam \c0.i17720_4_lut_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17720_4_lut_LC_12_15_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.i17720_4_lut_LC_12_15_4  (
            .in0(N__37423),
            .in1(N__37523),
            .in2(N__35839),
            .in3(N__28789),
            .lcout(),
            .ltout(\c0.n21307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_4_lut_adj_619_LC_12_15_5 .C_ON=1'b0;
    defparam \c0.i23_3_lut_4_lut_adj_619_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_4_lut_adj_619_LC_12_15_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.i23_3_lut_4_lut_adj_619_LC_12_15_5  (
            .in0(N__37342),
            .in1(N__28777),
            .in2(N__28771),
            .in3(N__37428),
            .lcout(n9_adj_3588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17990_4_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \c0.i17990_4_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17990_4_lut_LC_12_15_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.i17990_4_lut_LC_12_15_6  (
            .in0(N__37422),
            .in1(N__37522),
            .in2(N__33073),
            .in3(N__28975),
            .lcout(),
            .ltout(n21578_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i23_4_lut_adj_953_LC_12_15_7.C_ON=1'b0;
    defparam i23_4_lut_adj_953_LC_12_15_7.SEQ_MODE=4'b0000;
    defparam i23_4_lut_adj_953_LC_12_15_7.LUT_INIT=16'b1111000111100000;
    LogicCell40 i23_4_lut_adj_953_LC_12_15_7 (
            .in0(N__37340),
            .in1(N__37424),
            .in2(N__28969),
            .in3(N__28966),
            .lcout(n9_adj_3591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__7__5327_LC_12_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__7__5327_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__7__5327_LC_12_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_13__7__5327_LC_12_16_0  (
            .in0(N__46622),
            .in1(N__29991),
            .in2(_gnd_net_),
            .in3(N__28959),
            .lcout(data_out_frame_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71012),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17927_2_lut_LC_12_16_1 .C_ON=1'b0;
    defparam \c0.i17927_2_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17927_2_lut_LC_12_16_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i17927_2_lut_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__31199),
            .in2(_gnd_net_),
            .in3(N__34084),
            .lcout(\c0.n21467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i17743_3_lut_LC_12_16_2 .C_ON=1'b0;
    defparam \c0.tx.i17743_3_lut_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i17743_3_lut_LC_12_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i17743_3_lut_LC_12_16_2  (
            .in0(N__34227),
            .in1(N__33931),
            .in2(_gnd_net_),
            .in3(N__28920),
            .lcout(\c0.tx.n21330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_12_16_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_12_16_4 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_12_16_4  (
            .in0(N__33785),
            .in1(N__28921),
            .in2(N__33886),
            .in3(N__28927),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71012),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_643_LC_12_16_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_643_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_643_LC_12_16_5 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i2_3_lut_adj_643_LC_12_16_5  (
            .in0(N__36876),
            .in1(N__37316),
            .in2(_gnd_net_),
            .in3(N__36621),
            .lcout(\c0.n9753 ),
            .ltout(\c0.n9753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_647_LC_12_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_647_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_647_LC_12_16_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_647_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28912),
            .in3(N__40823),
            .lcout(\c0.n9755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__3__5339_LC_12_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__3__5339_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__3__5339_LC_12_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_12__3__5339_LC_12_16_7  (
            .in0(N__30259),
            .in1(N__28908),
            .in2(_gnd_net_),
            .in3(N__46623),
            .lcout(data_out_frame_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71012),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17972_3_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.i17972_3_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17972_3_lut_LC_12_17_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.i17972_3_lut_LC_12_17_0  (
            .in0(N__37301),
            .in1(N__40739),
            .in2(_gnd_net_),
            .in3(N__36588),
            .lcout(\c0.n21456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.i20_3_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_LC_12_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i20_3_lut_LC_12_17_1  (
            .in0(N__29059),
            .in1(N__29020),
            .in2(_gnd_net_),
            .in3(N__29038),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i17742_3_lut_LC_12_17_2 .C_ON=1'b0;
    defparam \c0.tx.i17742_3_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i17742_3_lut_LC_12_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i17742_3_lut_LC_12_17_2  (
            .in0(N__34220),
            .in1(N__30853),
            .in2(_gnd_net_),
            .in3(N__29214),
            .lcout(\c0.n21329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_12_17_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_12_17_5 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_12_17_5  (
            .in0(N__29304),
            .in1(N__28992),
            .in2(_gnd_net_),
            .in3(N__34222),
            .lcout(\c0.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71002),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_2__I_0_i2_3_lut_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_2__I_0_i2_3_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_2__I_0_i2_3_lut_LC_12_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Bit_Index_2__I_0_i2_3_lut_LC_12_17_6  (
            .in0(N__34221),
            .in1(N__31362),
            .in2(_gnd_net_),
            .in3(N__31323),
            .lcout(),
            .ltout(\c0.n2_adj_3556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_3_lut_adj_904_LC_12_17_7 .C_ON=1'b0;
    defparam \c0.i21_3_lut_adj_904_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i21_3_lut_adj_904_LC_12_17_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.i21_3_lut_adj_904_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__34098),
            .in2(N__29023),
            .in3(N__34160),
            .lcout(\c0.n7_adj_3557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_935_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_935_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_935_LC_12_18_0 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \c0.i11_4_lut_adj_935_LC_12_18_0  (
            .in0(N__34168),
            .in1(N__29186),
            .in2(N__29170),
            .in3(N__29014),
            .lcout(),
            .ltout(\c0.n19001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_3_lut_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.i31_3_lut_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i31_3_lut_LC_12_18_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.i31_3_lut_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__29298),
            .in2(N__29008),
            .in3(N__29089),
            .lcout(\c0.n30_adj_3559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_690_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_690_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_690_LC_12_18_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i2_2_lut_adj_690_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__39590),
            .in2(_gnd_net_),
            .in3(N__38968),
            .lcout(\c0.n6_adj_3338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_4_lut_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_4_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_4_lut_LC_12_18_3 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \c0.tx.i2_4_lut_4_lut_LC_12_18_3  (
            .in0(N__34095),
            .in1(N__29302),
            .in2(N__29329),
            .in3(N__29169),
            .lcout(\c0.n12498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_18_4 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \c0.tx.i1_3_lut_4_lut_LC_12_18_4  (
            .in0(N__29168),
            .in1(N__29324),
            .in2(N__29305),
            .in3(N__34094),
            .lcout(n4_adj_3580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_12_18_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_12_18_5 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_12_18_5  (
            .in0(N__33765),
            .in1(N__29215),
            .in2(N__33877),
            .in3(N__29224),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71013),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_1_lut_LC_12_18_6 .C_ON=1'b0;
    defparam \c0.tx.i1_1_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_1_lut_LC_12_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.i1_1_lut_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34092),
            .lcout(\c0.n12512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.i12_3_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_LC_12_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \c0.i12_3_lut_LC_12_18_7  (
            .in0(N__34093),
            .in1(N__29164),
            .in2(_gnd_net_),
            .in3(N__34169),
            .lcout(\c0.n19023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_691_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_691_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_691_LC_12_19_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_691_LC_12_19_1  (
            .in0(N__37149),
            .in1(N__29527),
            .in2(_gnd_net_),
            .in3(N__37128),
            .lcout(\c0.n19052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_12_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.i2_2_lut_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__56126),
            .in2(_gnd_net_),
            .in3(N__39232),
            .lcout(\c0.rx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_390_Select_2_i2_4_lut_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.select_390_Select_2_i2_4_lut_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_390_Select_2_i2_4_lut_LC_12_19_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.select_390_Select_2_i2_4_lut_LC_12_19_5  (
            .in0(N__38972),
            .in1(N__42505),
            .in2(N__39076),
            .in3(N__35419),
            .lcout(n8112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12190_4_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.i12190_4_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i12190_4_lut_LC_12_19_6 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \c0.i12190_4_lut_LC_12_19_6  (
            .in0(N__29650),
            .in1(N__40284),
            .in2(N__38167),
            .in3(N__38194),
            .lcout(\c0.n4812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_229_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_229_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_229_LC_12_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_229_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__29355),
            .in2(_gnd_net_),
            .in3(N__41404),
            .lcout(\c0.n18609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17645_2_lut_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.i17645_2_lut_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17645_2_lut_LC_12_21_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i17645_2_lut_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__39486),
            .in2(_gnd_net_),
            .in3(N__29523),
            .lcout(\c0.n21231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_915_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_915_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_915_LC_12_21_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_915_LC_12_21_2  (
            .in0(N__31575),
            .in1(N__38245),
            .in2(N__31429),
            .in3(N__38325),
            .lcout(\c0.n21053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_425_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_425_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_425_LC_12_21_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_425_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__38361),
            .in2(_gnd_net_),
            .in3(N__35208),
            .lcout(\c0.FRAME_MATCHER_state_31_N_1864_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_22_i6_2_lut_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.select_357_Select_22_i6_2_lut_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_22_i6_2_lut_LC_12_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_22_i6_2_lut_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__60695),
            .in2(_gnd_net_),
            .in3(N__34390),
            .lcout(\c0.n6_adj_3178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_689_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_689_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_689_LC_12_22_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i5_3_lut_adj_689_LC_12_22_0  (
            .in0(N__29425),
            .in1(N__29404),
            .in2(_gnd_net_),
            .in3(N__29377),
            .lcout(\c0.n15850 ),
            .ltout(\c0.n15850_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_12_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_4_lut_LC_12_22_1  (
            .in0(N__29469),
            .in1(N__29560),
            .in2(N__29371),
            .in3(N__29335),
            .lcout(\c0.n11427 ),
            .ltout(\c0.n11427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_279_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_279_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_279_LC_12_22_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_279_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29368),
            .in3(N__39568),
            .lcout(n11289),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_682_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_682_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_682_LC_12_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_682_LC_12_22_3  (
            .in0(N__40324),
            .in1(N__29365),
            .in2(N__29749),
            .in3(N__29354),
            .lcout(\c0.n19045 ),
            .ltout(\c0.n19045_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_586_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_586_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_586_LC_12_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_586_LC_12_22_4  (
            .in0(N__41505),
            .in1(N__29736),
            .in2(N__29338),
            .in3(N__29549),
            .lcout(\c0.n4_adj_3046 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_577_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_577_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_577_LC_12_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_577_LC_12_22_5  (
            .in0(N__29569),
            .in1(N__29626),
            .in2(N__29635),
            .in3(N__29599),
            .lcout(\c0.n70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_687_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_687_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_687_LC_12_22_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i5_3_lut_adj_687_LC_12_22_6  (
            .in0(N__29625),
            .in1(N__29598),
            .in2(_gnd_net_),
            .in3(N__29568),
            .lcout(\c0.n19050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_594_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_594_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_594_LC_12_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_594_LC_12_22_7  (
            .in0(N__29737),
            .in1(N__29470),
            .in2(N__29554),
            .in3(N__41506),
            .lcout(\c0.n63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_12_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_12_23_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_12_23_2  (
            .in0(N__29509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71064),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_511_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_511_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_511_LC_12_23_3 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \c0.i1_4_lut_adj_511_LC_12_23_3  (
            .in0(N__42518),
            .in1(N__37960),
            .in2(N__29695),
            .in3(N__31543),
            .lcout(\c0.n18601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_251_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_251_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_251_LC_12_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_251_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__29495),
            .in2(_gnd_net_),
            .in3(N__41435),
            .lcout(\c0.n18659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i16_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_12_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_12_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__29496),
            .in2(_gnd_net_),
            .in3(N__40545),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71077),
            .ce(),
            .sr(N__29476));
    defparam \c0.i3_4_lut_adj_674_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_674_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_674_LC_12_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_674_LC_12_25_0  (
            .in0(N__31627),
            .in1(N__35472),
            .in2(N__31690),
            .in3(N__29450),
            .lcout(\c0.n19146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_858_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_858_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_858_LC_12_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_858_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__29451),
            .in2(_gnd_net_),
            .in3(N__41467),
            .lcout(\c0.n18633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_680_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_680_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_680_LC_12_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_680_LC_12_25_3  (
            .in0(N__29824),
            .in1(N__29792),
            .in2(N__29694),
            .in3(N__29776),
            .lcout(\c0.n17_adj_3486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_923_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_923_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_923_LC_12_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_923_LC_12_25_5  (
            .in0(N__41468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31688),
            .lcout(\c0.n18681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_12_26_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_12_26_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_12_26_6  (
            .in0(_gnd_net_),
            .in1(N__29729),
            .in2(_gnd_net_),
            .in3(N__40548),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71103),
            .ce(),
            .sr(N__29707));
    defparam \c0.FRAME_MATCHER_state_i30_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_12_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_12_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_12_27_0  (
            .in0(_gnd_net_),
            .in1(N__40549),
            .in2(_gnd_net_),
            .in3(N__29687),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71117),
            .ce(),
            .sr(N__29665));
    defparam \c0.FRAME_MATCHER_state_i4_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_12_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_12_28_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_12_28_0  (
            .in0(N__40550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31626),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71133),
            .ce(),
            .sr(N__31606));
    defparam \c0.FRAME_MATCHER_i_i3_LC_13_6_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i3_LC_13_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_13_6_0 .LUT_INIT=16'b1111111111010101;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_13_6_0  (
            .in0(N__38670),
            .in1(N__60710),
            .in2(N__40084),
            .in3(N__31723),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71150),
            .ce(),
            .sr(N__46937));
    defparam \c0.select_357_Select_2_i6_2_lut_LC_13_6_1 .C_ON=1'b0;
    defparam \c0.select_357_Select_2_i6_2_lut_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_2_i6_2_lut_LC_13_6_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.select_357_Select_2_i6_2_lut_LC_13_6_1  (
            .in0(N__60709),
            .in1(_gnd_net_),
            .in2(N__59944),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n6_adj_3143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_13_6_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i2_LC_13_6_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_13_6_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_13_6_2  (
            .in0(N__38984),
            .in1(N__31594),
            .in2(N__29653),
            .in3(N__35437),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71150),
            .ce(),
            .sr(N__46937));
    defparam \c0.i1_2_lut_3_lut_adj_675_LC_13_6_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_675_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_675_LC_13_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_675_LC_13_6_3  (
            .in0(N__59921),
            .in1(N__60048),
            .in2(_gnd_net_),
            .in3(N__40071),
            .lcout(\c0.n4_adj_3227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_63_i9_2_lut_3_lut_LC_13_6_6 .C_ON=1'b0;
    defparam \c0.equal_63_i9_2_lut_3_lut_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_63_i9_2_lut_3_lut_LC_13_6_6 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \c0.equal_63_i9_2_lut_3_lut_LC_13_6_6  (
            .in0(N__60049),
            .in1(_gnd_net_),
            .in2(N__60263),
            .in3(N__59923),
            .lcout(\c0.n9_adj_3351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_64_i9_2_lut_3_lut_LC_13_6_7 .C_ON=1'b0;
    defparam \c0.equal_64_i9_2_lut_3_lut_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.equal_64_i9_2_lut_3_lut_LC_13_6_7 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.equal_64_i9_2_lut_3_lut_LC_13_6_7  (
            .in0(N__59922),
            .in1(N__60242),
            .in2(_gnd_net_),
            .in3(N__60047),
            .lcout(\c0.n9_adj_3251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_adj_948_LC_13_7_4 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_adj_948_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_adj_948_LC_13_7_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter1.i3_4_lut_adj_948_LC_13_7_4  (
            .in0(N__29913),
            .in1(N__29884),
            .in2(N__29869),
            .in3(N__29920),
            .lcout(count_enable_adj_3586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_delayed_67_LC_13_7_7 .C_ON=1'b0;
    defparam \quad_counter1.A_delayed_67_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_delayed_67_LC_13_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.A_delayed_67_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29866),
            .lcout(\quad_counter1.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71136),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_13_8_1 .C_ON=1'b0;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_13_8_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter1.A_filtered_I_0_2_lut_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__29883),
            .in2(_gnd_net_),
            .in3(N__29868),
            .lcout(\quad_counter1.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_delayed_68_LC_13_8_2 .C_ON=1'b0;
    defparam \quad_counter1.B_delayed_68_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_delayed_68_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.B_delayed_68_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29914),
            .lcout(\quad_counter1.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71120),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1063_1_lut_2_lut_LC_13_8_7 .C_ON=1'b0;
    defparam \quad_counter1.i1063_1_lut_2_lut_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1063_1_lut_2_lut_LC_13_8_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter1.i1063_1_lut_2_lut_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__29882),
            .in2(_gnd_net_),
            .in3(N__29867),
            .lcout(\quad_counter1.n2301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_1_LC_13_9_0 .C_ON=1'b1;
    defparam \quad_counter1.add_635_1_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_1_LC_13_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter1.add_635_1_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__30498),
            .in2(N__30564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\quad_counter1.n17314 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_2_lut_LC_13_9_1 .C_ON=1'b1;
    defparam \quad_counter1.add_635_2_lut_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_2_lut_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_2_lut_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__29833),
            .in2(N__37212),
            .in3(N__29827),
            .lcout(n2345),
            .ltout(),
            .carryin(\quad_counter1.n17314 ),
            .carryout(\quad_counter1.n17315 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_3_lut_LC_13_9_2 .C_ON=1'b1;
    defparam \quad_counter1.add_635_3_lut_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_3_lut_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_3_lut_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__30499),
            .in2(N__33702),
            .in3(N__30076),
            .lcout(n2344),
            .ltout(),
            .carryin(\quad_counter1.n17315 ),
            .carryout(\quad_counter1.n17316 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_4_lut_LC_13_9_3 .C_ON=1'b1;
    defparam \quad_counter1.add_635_4_lut_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_4_lut_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_4_lut_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__30505),
            .in2(N__31090),
            .in3(N__30061),
            .lcout(n2343),
            .ltout(),
            .carryin(\quad_counter1.n17316 ),
            .carryout(\quad_counter1.n17317 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_5_lut_LC_13_9_4 .C_ON=1'b1;
    defparam \quad_counter1.add_635_5_lut_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_5_lut_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_5_lut_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__30500),
            .in2(N__33037),
            .in3(N__30058),
            .lcout(n2342),
            .ltout(),
            .carryin(\quad_counter1.n17317 ),
            .carryout(\quad_counter1.n17318 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_6_lut_LC_13_9_5 .C_ON=1'b1;
    defparam \quad_counter1.add_635_6_lut_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_6_lut_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_6_lut_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__30506),
            .in2(N__30919),
            .in3(N__30043),
            .lcout(n2341),
            .ltout(),
            .carryin(\quad_counter1.n17318 ),
            .carryout(\quad_counter1.n17319 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_7_lut_LC_13_9_6 .C_ON=1'b1;
    defparam \quad_counter1.add_635_7_lut_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_7_lut_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_7_lut_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__30501),
            .in2(N__32853),
            .in3(N__30040),
            .lcout(n2340),
            .ltout(),
            .carryin(\quad_counter1.n17319 ),
            .carryout(\quad_counter1.n17320 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_8_lut_LC_13_9_7 .C_ON=1'b1;
    defparam \quad_counter1.add_635_8_lut_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_8_lut_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_8_lut_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__30507),
            .in2(N__30037),
            .in3(N__29995),
            .lcout(n2339),
            .ltout(),
            .carryin(\quad_counter1.n17320 ),
            .carryout(\quad_counter1.n17321 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_9_lut_LC_13_10_0 .C_ON=1'b1;
    defparam \quad_counter1.add_635_9_lut_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_9_lut_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_9_lut_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__30565),
            .in2(N__29992),
            .in3(N__29947),
            .lcout(n2338),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\quad_counter1.n17322 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_10_lut_LC_13_10_1 .C_ON=1'b1;
    defparam \quad_counter1.add_635_10_lut_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_10_lut_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_10_lut_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__30569),
            .in2(N__36369),
            .in3(N__29932),
            .lcout(n2337),
            .ltout(),
            .carryin(\quad_counter1.n17322 ),
            .carryout(\quad_counter1.n17323 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_11_lut_LC_13_10_2 .C_ON=1'b1;
    defparam \quad_counter1.add_635_11_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_11_lut_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_11_lut_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__30566),
            .in2(N__31167),
            .in3(N__29923),
            .lcout(n2336),
            .ltout(),
            .carryin(\quad_counter1.n17323 ),
            .carryout(\quad_counter1.n17324 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_12_lut_LC_13_10_3 .C_ON=1'b1;
    defparam \quad_counter1.add_635_12_lut_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_12_lut_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_12_lut_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__30570),
            .in2(N__30291),
            .in3(N__30262),
            .lcout(n2335),
            .ltout(),
            .carryin(\quad_counter1.n17324 ),
            .carryout(\quad_counter1.n17325 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_13_lut_LC_13_10_4 .C_ON=1'b1;
    defparam \quad_counter1.add_635_13_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_13_lut_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_13_lut_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__30567),
            .in2(N__30255),
            .in3(N__30226),
            .lcout(n2334),
            .ltout(),
            .carryin(\quad_counter1.n17325 ),
            .carryout(\quad_counter1.n17326 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_14_lut_LC_13_10_5 .C_ON=1'b1;
    defparam \quad_counter1.add_635_14_lut_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_14_lut_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_14_lut_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__30571),
            .in2(N__37060),
            .in3(N__30223),
            .lcout(n2333),
            .ltout(),
            .carryin(\quad_counter1.n17326 ),
            .carryout(\quad_counter1.n17327 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_15_lut_LC_13_10_6 .C_ON=1'b1;
    defparam \quad_counter1.add_635_15_lut_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_15_lut_LC_13_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_15_lut_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__30568),
            .in2(N__30219),
            .in3(N__30190),
            .lcout(n2332),
            .ltout(),
            .carryin(\quad_counter1.n17327 ),
            .carryout(\quad_counter1.n17328 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_16_lut_LC_13_10_7 .C_ON=1'b1;
    defparam \quad_counter1.add_635_16_lut_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_16_lut_LC_13_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_16_lut_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__30572),
            .in2(N__30186),
            .in3(N__30157),
            .lcout(n2331),
            .ltout(),
            .carryin(\quad_counter1.n17328 ),
            .carryout(\quad_counter1.n17329 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_17_lut_LC_13_11_0 .C_ON=1'b1;
    defparam \quad_counter1.add_635_17_lut_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_17_lut_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_17_lut_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__30573),
            .in2(N__30153),
            .in3(N__30124),
            .lcout(n2330),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\quad_counter1.n17330 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_18_lut_LC_13_11_1 .C_ON=1'b1;
    defparam \quad_counter1.add_635_18_lut_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_18_lut_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_18_lut_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__30577),
            .in2(N__30117),
            .in3(N__30088),
            .lcout(n2329),
            .ltout(),
            .carryin(\quad_counter1.n17330 ),
            .carryout(\quad_counter1.n17331 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_19_lut_LC_13_11_2 .C_ON=1'b1;
    defparam \quad_counter1.add_635_19_lut_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_19_lut_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_19_lut_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__30574),
            .in2(N__31056),
            .in3(N__30079),
            .lcout(n2328),
            .ltout(),
            .carryin(\quad_counter1.n17331 ),
            .carryout(\quad_counter1.n17332 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_20_lut_LC_13_11_3 .C_ON=1'b1;
    defparam \quad_counter1.add_635_20_lut_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_20_lut_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_20_lut_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__30578),
            .in2(N__33294),
            .in3(N__30418),
            .lcout(n2327),
            .ltout(),
            .carryin(\quad_counter1.n17332 ),
            .carryout(\quad_counter1.n17333 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_21_lut_LC_13_11_4 .C_ON=1'b1;
    defparam \quad_counter1.add_635_21_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_21_lut_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_21_lut_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__30575),
            .in2(N__30415),
            .in3(N__30376),
            .lcout(n2326),
            .ltout(),
            .carryin(\quad_counter1.n17333 ),
            .carryout(\quad_counter1.n17334 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_22_lut_LC_13_11_5 .C_ON=1'b1;
    defparam \quad_counter1.add_635_22_lut_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_22_lut_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_22_lut_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__30579),
            .in2(N__30372),
            .in3(N__30343),
            .lcout(n2325),
            .ltout(),
            .carryin(\quad_counter1.n17334 ),
            .carryout(\quad_counter1.n17335 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_23_lut_LC_13_11_6 .C_ON=1'b1;
    defparam \quad_counter1.add_635_23_lut_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_23_lut_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_23_lut_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__30576),
            .in2(N__32965),
            .in3(N__30340),
            .lcout(n2324),
            .ltout(),
            .carryin(\quad_counter1.n17335 ),
            .carryout(\quad_counter1.n17336 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_24_lut_LC_13_11_7 .C_ON=1'b1;
    defparam \quad_counter1.add_635_24_lut_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_24_lut_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_24_lut_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__30580),
            .in2(N__30337),
            .in3(N__30310),
            .lcout(n2323),
            .ltout(),
            .carryin(\quad_counter1.n17336 ),
            .carryout(\quad_counter1.n17337 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_25_lut_LC_13_12_0 .C_ON=1'b1;
    defparam \quad_counter1.add_635_25_lut_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_25_lut_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_25_lut_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__30581),
            .in2(N__36322),
            .in3(N__30307),
            .lcout(n2322),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\quad_counter1.n17338 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_26_lut_LC_13_12_1 .C_ON=1'b1;
    defparam \quad_counter1.add_635_26_lut_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_26_lut_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_26_lut_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__30752),
            .in2(N__30598),
            .in3(N__30298),
            .lcout(n2321),
            .ltout(),
            .carryin(\quad_counter1.n17338 ),
            .carryout(\quad_counter1.n17339 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_27_lut_LC_13_12_2 .C_ON=1'b1;
    defparam \quad_counter1.add_635_27_lut_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_27_lut_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_27_lut_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__30585),
            .in2(N__31111),
            .in3(N__30295),
            .lcout(n2320),
            .ltout(),
            .carryin(\quad_counter1.n17339 ),
            .carryout(\quad_counter1.n17340 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_28_lut_LC_13_12_3 .C_ON=1'b1;
    defparam \quad_counter1.add_635_28_lut_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_28_lut_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_28_lut_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__32798),
            .in2(N__30599),
            .in3(N__30688),
            .lcout(n2319),
            .ltout(),
            .carryin(\quad_counter1.n17340 ),
            .carryout(\quad_counter1.n17341 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_29_lut_LC_13_12_4 .C_ON=1'b1;
    defparam \quad_counter1.add_635_29_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_29_lut_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_29_lut_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__30589),
            .in2(N__30684),
            .in3(N__30655),
            .lcout(n2318),
            .ltout(),
            .carryin(\quad_counter1.n17341 ),
            .carryout(\quad_counter1.n17342 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_30_lut_LC_13_12_5 .C_ON=1'b1;
    defparam \quad_counter1.add_635_30_lut_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_30_lut_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_30_lut_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__36078),
            .in2(N__30600),
            .in3(N__30652),
            .lcout(n2317),
            .ltout(),
            .carryin(\quad_counter1.n17342 ),
            .carryout(\quad_counter1.n17343 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_31_lut_LC_13_12_6 .C_ON=1'b1;
    defparam \quad_counter1.add_635_31_lut_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_31_lut_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_31_lut_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__30593),
            .in2(N__33391),
            .in3(N__30649),
            .lcout(n2316),
            .ltout(),
            .carryin(\quad_counter1.n17343 ),
            .carryout(\quad_counter1.n17344 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_32_lut_LC_13_12_7 .C_ON=1'b1;
    defparam \quad_counter1.add_635_32_lut_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_32_lut_LC_13_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_635_32_lut_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__30642),
            .in2(N__30601),
            .in3(N__30604),
            .lcout(n2315),
            .ltout(),
            .carryin(\quad_counter1.n17344 ),
            .carryout(\quad_counter1.n17345 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_635_33_lut_LC_13_13_0 .C_ON=1'b0;
    defparam \quad_counter1.add_635_33_lut_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_635_33_lut_LC_13_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter1.add_635_33_lut_LC_13_13_0  (
            .in0(N__30869),
            .in1(N__30597),
            .in2(_gnd_net_),
            .in3(N__30457),
            .lcout(n2314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i31_LC_13_13_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i31_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i31_LC_13_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i31_LC_13_13_1  (
            .in0(N__36229),
            .in1(N__30454),
            .in2(_gnd_net_),
            .in3(N__30870),
            .lcout(encoder1_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71052),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i0_LC_13_13_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i0_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i0_LC_13_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i0_LC_13_13_2  (
            .in0(N__30448),
            .in1(N__36230),
            .in2(_gnd_net_),
            .in3(N__37211),
            .lcout(encoder1_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71052),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_13_13_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_13_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_13_13_3  (
            .in0(N__30970),
            .in1(N__30438),
            .in2(_gnd_net_),
            .in3(N__40884),
            .lcout(\c0.n11_adj_3462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__4__5330_LC_13_13_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__4__5330_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__4__5330_LC_13_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_13__4__5330_LC_13_13_5  (
            .in0(N__46724),
            .in1(N__30918),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(data_out_frame_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71052),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__7__5351_LC_13_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__7__5351_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__7__5351_LC_13_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__7__5351_LC_13_13_6  (
            .in0(N__30871),
            .in1(N__33231),
            .in2(_gnd_net_),
            .in3(N__46725),
            .lcout(data_out_frame_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71052),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i25_LC_13_13_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i25_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i25_LC_13_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i25_LC_13_13_7  (
            .in0(N__36228),
            .in1(N__31109),
            .in2(_gnd_net_),
            .in3(N__30859),
            .lcout(encoder1_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71052),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_13_14_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_14_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_13_14_0  (
            .in0(N__33799),
            .in1(N__33873),
            .in2(N__30852),
            .in3(N__37243),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17700_3_lut_LC_13_14_1 .C_ON=1'b0;
    defparam \c0.i17700_3_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17700_3_lut_LC_13_14_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i17700_3_lut_LC_13_14_1  (
            .in0(N__30832),
            .in1(N__30813),
            .in2(_gnd_net_),
            .in3(N__40885),
            .lcout(\c0.n21287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__1__5373_LC_13_14_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__1__5373_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__1__5373_LC_13_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_8__1__5373_LC_13_14_2  (
            .in0(N__46646),
            .in1(N__30786),
            .in2(_gnd_net_),
            .in3(N__31218),
            .lcout(data_out_frame_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__0__5358_LC_13_14_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__0__5358_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__0__5358_LC_13_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__0__5358_LC_13_14_3  (
            .in0(N__30763),
            .in1(N__33628),
            .in2(_gnd_net_),
            .in3(N__46648),
            .lcout(data_out_frame_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__4__5434_LC_13_14_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__4__5434_LC_13_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__4__5434_LC_13_14_4 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \c0.data_out_frame_0__4__5434_LC_13_14_4  (
            .in0(N__39493),
            .in1(N__30735),
            .in2(N__38996),
            .in3(N__37091),
            .lcout(\c0.data_out_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__0__5374_LC_13_14_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__0__5374_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__0__5374_LC_13_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_8__0__5374_LC_13_14_5  (
            .in0(N__30713),
            .in1(N__33591),
            .in2(_gnd_net_),
            .in3(N__46650),
            .lcout(data_out_frame_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__0__5366_LC_13_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__0__5366_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__0__5366_LC_13_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_9__0__5366_LC_13_14_6  (
            .in0(N__46647),
            .in1(N__31144),
            .in2(_gnd_net_),
            .in3(N__33573),
            .lcout(data_out_frame_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__1__5357_LC_13_14_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__1__5357_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__1__5357_LC_13_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__1__5357_LC_13_14_7  (
            .in0(N__31110),
            .in1(N__30994),
            .in2(_gnd_net_),
            .in3(N__46649),
            .lcout(data_out_frame_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71040),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__2__5332_LC_13_15_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__2__5332_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__2__5332_LC_13_15_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame_13__2__5332_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__46651),
            .in2(N__31033),
            .in3(N__31086),
            .lcout(data_out_frame_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71031),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__1__5349_LC_13_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__1__5349_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__1__5349_LC_13_15_1 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.data_out_frame_11__1__5349_LC_13_15_1  (
            .in0(N__30981),
            .in1(N__31060),
            .in2(N__46765),
            .in3(_gnd_net_),
            .lcout(data_out_frame_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71031),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_15_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_15_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_15_2  (
            .in0(N__40883),
            .in1(_gnd_net_),
            .in2(N__31032),
            .in3(N__31017),
            .lcout(\c0.n11_adj_3108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18029_LC_13_15_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18029_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18029_LC_13_15_3 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18029_LC_13_15_3  (
            .in0(N__30993),
            .in1(N__40882),
            .in2(N__30982),
            .in3(N__36633),
            .lcout(\c0.n21605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i276_3_lut_4_lut_LC_13_15_4 .C_ON=1'b0;
    defparam \c0.i276_3_lut_4_lut_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i276_3_lut_4_lut_LC_13_15_4 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \c0.i276_3_lut_4_lut_LC_13_15_4  (
            .in0(N__30953),
            .in1(N__33507),
            .in2(N__31302),
            .in3(N__31272),
            .lcout(\c0.n700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__5__5329_LC_13_15_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__5__5329_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__5__5329_LC_13_15_5 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame_13__5__5329_LC_13_15_5  (
            .in0(N__32857),
            .in1(N__30969),
            .in2(N__46766),
            .in3(_gnd_net_),
            .lcout(data_out_frame_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71031),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18009_3_lut_4_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \c0.i18009_3_lut_4_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i18009_3_lut_4_lut_LC_13_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.i18009_3_lut_4_lut_LC_13_15_6  (
            .in0(N__30954),
            .in1(N__33508),
            .in2(N__31303),
            .in3(N__31273),
            .lcout(\c0.tx_transmit_N_2443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_264_LC_13_16_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_264_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_264_LC_13_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i3_4_lut_adj_264_LC_13_16_0  (
            .in0(N__37412),
            .in1(N__36864),
            .in2(N__37335),
            .in3(N__34264),
            .lcout(\c0.n15842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17978_4_lut_LC_13_16_1 .C_ON=1'b0;
    defparam \c0.i17978_4_lut_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17978_4_lut_LC_13_16_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.i17978_4_lut_LC_13_16_1  (
            .in0(N__36624),
            .in1(N__31264),
            .in2(N__36926),
            .in3(N__33163),
            .lcout(\c0.n21566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_13_16_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_13_16_3 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_13_16_3  (
            .in0(N__33800),
            .in1(N__31201),
            .in2(N__33885),
            .in3(N__31252),
            .lcout(\c0.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71021),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21605_bdd_4_lut_LC_13_16_4 .C_ON=1'b0;
    defparam \c0.n21605_bdd_4_lut_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.n21605_bdd_4_lut_LC_13_16_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n21605_bdd_4_lut_LC_13_16_4  (
            .in0(N__31246),
            .in1(N__31228),
            .in2(N__31222),
            .in3(N__36622),
            .lcout(),
            .ltout(\c0.n21608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17974_4_lut_LC_13_16_5 .C_ON=1'b0;
    defparam \c0.i17974_4_lut_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17974_4_lut_LC_13_16_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.i17974_4_lut_LC_13_16_5  (
            .in0(N__36623),
            .in1(N__36885),
            .in2(N__31204),
            .in3(N__31342),
            .lcout(\c0.n21562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_16_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_16_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17959_2_lut_2_lut_LC_13_16_7 .C_ON=1'b0;
    defparam \c0.i17959_2_lut_2_lut_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17959_2_lut_2_lut_LC_13_16_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i17959_2_lut_2_lut_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__31200),
            .in2(_gnd_net_),
            .in3(N__34083),
            .lcout(\c0.n21466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__1__5341_LC_13_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__1__5341_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__1__5341_LC_13_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_12__1__5341_LC_13_17_0  (
            .in0(N__31174),
            .in1(N__31351),
            .in2(_gnd_net_),
            .in3(N__46645),
            .lcout(data_out_frame_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71009),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__5__5393_LC_13_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__5__5393_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__5__5393_LC_13_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_5__5__5393_LC_13_17_1  (
            .in0(N__46644),
            .in1(N__36448),
            .in2(_gnd_net_),
            .in3(N__33735),
            .lcout(data_out_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71009),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_4_lut_adj_610_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.i24_3_lut_4_lut_adj_610_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_4_lut_adj_610_LC_13_17_2 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.i24_3_lut_4_lut_adj_610_LC_13_17_2  (
            .in0(N__37312),
            .in1(N__31375),
            .in2(N__37443),
            .in3(N__35953),
            .lcout(),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_13_17_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_13_17_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_13_17_3  (
            .in0(N__33861),
            .in1(N__31366),
            .in2(N__31369),
            .in3(N__33798),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71009),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_13_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_13_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_13_17_6  (
            .in0(N__33670),
            .in1(N__31350),
            .in2(_gnd_net_),
            .in3(N__40738),
            .lcout(\c0.n11_adj_3104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_13_17_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_17_7 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_13_17_7  (
            .in0(N__31324),
            .in1(N__33797),
            .in2(N__33878),
            .in3(N__31336),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71009),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1399__i0_LC_13_18_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i0_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i0_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i0_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__31536),
            .in2(N__40825),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\c0.n17346 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i1_LC_13_18_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i1_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i1_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__36589),
            .in2(_gnd_net_),
            .in3(N__31312),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n17346 ),
            .carryout(\c0.n17347 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i2_LC_13_18_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i2_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i2_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i2_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__36925),
            .in2(_gnd_net_),
            .in3(N__31309),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(\c0.n17347 ),
            .carryout(\c0.n17348 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i3_LC_13_18_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i3_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i3_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i3_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__37311),
            .in2(_gnd_net_),
            .in3(N__31306),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(\c0.n17348 ),
            .carryout(\c0.n17349 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i4_LC_13_18_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i4_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i4_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i4_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__37408),
            .in2(_gnd_net_),
            .in3(N__31459),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(\c0.n17349 ),
            .carryout(\c0.n17350 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i5_LC_13_18_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i5_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i5_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i5_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__33848),
            .in2(_gnd_net_),
            .in3(N__31456),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(\c0.n17350 ),
            .carryout(\c0.n17351 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i6_LC_13_18_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1399__i6_LC_13_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i6_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i6_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__33540),
            .in2(_gnd_net_),
            .in3(N__31453),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(\c0.n17351 ),
            .carryout(\c0.n17352 ),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.byte_transmit_counter_1399__i7_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1399__i7_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1399__i7_LC_13_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1399__i7_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__33522),
            .in2(_gnd_net_),
            .in3(N__31450),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71022),
            .ce(N__31408),
            .sr(N__31393));
    defparam \c0.i18005_4_lut_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.i18005_4_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i18005_4_lut_LC_13_19_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \c0.i18005_4_lut_LC_13_19_1  (
            .in0(N__42512),
            .in1(N__31440),
            .in2(N__31428),
            .in3(N__31468),
            .lcout(\c0.n12326 ),
            .ltout(\c0.n12326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18001_2_lut_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.i18001_2_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i18001_2_lut_LC_13_19_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \c0.i18001_2_lut_LC_13_19_2  (
            .in0(N__39595),
            .in1(_gnd_net_),
            .in2(N__31396),
            .in3(_gnd_net_),
            .lcout(\c0.n12758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_741_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_741_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_741_LC_13_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_741_LC_13_19_3  (
            .in0(N__40092),
            .in1(N__40267),
            .in2(N__59965),
            .in3(N__38193),
            .lcout(),
            .ltout(\c0.n4_adj_3263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12196_4_lut_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.i12196_4_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12196_4_lut_LC_13_19_4 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \c0.i12196_4_lut_LC_13_19_4  (
            .in0(N__38153),
            .in1(N__60272),
            .in2(N__31381),
            .in3(N__60115),
            .lcout(\c0.n936 ),
            .ltout(\c0.n936_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_671_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_671_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_671_LC_13_19_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_671_LC_13_19_5  (
            .in0(N__42516),
            .in1(_gnd_net_),
            .in2(N__31378),
            .in3(N__42330),
            .lcout(\c0.n10_adj_3081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17902_4_lut_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.i17902_4_lut_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17902_4_lut_LC_13_19_7 .LUT_INIT=16'b1000000010110000;
    LogicCell40 \c0.i17902_4_lut_LC_13_19_7  (
            .in0(N__31537),
            .in1(N__39596),
            .in2(N__42520),
            .in3(N__38848),
            .lcout(\c0.n21420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_18_i6_2_lut_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.select_357_Select_18_i6_2_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_18_i6_2_lut_LC_13_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_357_Select_18_i6_2_lut_LC_13_20_0  (
            .in0(N__60692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38046),
            .lcout(\c0.n6_adj_3186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_313_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_313_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_313_LC_13_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_313_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__31507),
            .in2(_gnd_net_),
            .in3(N__41403),
            .lcout(\c0.n18627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_13_i6_2_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.select_357_Select_13_i6_2_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_13_i6_2_lut_LC_13_20_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_357_Select_13_i6_2_lut_LC_13_20_2  (
            .in0(N__60691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34848),
            .lcout(\c0.n6_adj_3162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_949_LC_13_20_4.C_ON=1'b0;
    defparam i2_4_lut_adj_949_LC_13_20_4.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_949_LC_13_20_4.LUT_INIT=16'b0000000010100010;
    LogicCell40 i2_4_lut_adj_949_LC_13_20_4 (
            .in0(N__42506),
            .in1(N__39075),
            .in2(N__38977),
            .in3(N__35418),
            .lcout(n20764),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_20_i6_2_lut_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.select_357_Select_20_i6_2_lut_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_20_i6_2_lut_LC_13_20_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_20_i6_2_lut_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__60694),
            .in2(_gnd_net_),
            .in3(N__34483),
            .lcout(\c0.n6_adj_3182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_19_i6_2_lut_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.select_357_Select_19_i6_2_lut_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_19_i6_2_lut_LC_13_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_19_i6_2_lut_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__34594),
            .in2(_gnd_net_),
            .in3(N__60693),
            .lcout(\c0.n6_adj_3184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_21_i6_2_lut_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.select_357_Select_21_i6_2_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_21_i6_2_lut_LC_13_21_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_357_Select_21_i6_2_lut_LC_13_21_0  (
            .in0(N__60690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35079),
            .lcout(\c0.n6_adj_3180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16066_2_lut_4_lut_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.i16066_2_lut_4_lut_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16066_2_lut_4_lut_LC_13_21_2 .LUT_INIT=16'b1111011111110010;
    LogicCell40 \c0.i16066_2_lut_4_lut_LC_13_21_2  (
            .in0(N__38925),
            .in1(N__38841),
            .in2(N__39597),
            .in3(N__39064),
            .lcout(\c0.n19650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_13_21_4 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \c0.i1_4_lut_LC_13_21_4  (
            .in0(N__38380),
            .in1(N__35095),
            .in2(N__34729),
            .in3(N__38326),
            .lcout(\c0.n5_adj_2999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_17_i6_2_lut_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.select_357_Select_17_i6_2_lut_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_17_i6_2_lut_LC_13_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_17_i6_2_lut_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__60689),
            .in2(_gnd_net_),
            .in3(N__35055),
            .lcout(\c0.n6_adj_3188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16054_2_lut_3_lut_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.i16054_2_lut_3_lut_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16054_2_lut_3_lut_LC_13_22_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i16054_2_lut_3_lut_LC_13_22_0  (
            .in0(N__42508),
            .in1(N__31571),
            .in2(_gnd_net_),
            .in3(N__42323),
            .lcout(\c0.n19638 ),
            .ltout(\c0.n19638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17686_3_lut_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i17686_3_lut_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17686_3_lut_LC_13_22_1 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \c0.i17686_3_lut_LC_13_22_1  (
            .in0(N__38362),
            .in1(_gnd_net_),
            .in2(N__31588),
            .in3(N__34757),
            .lcout(\c0.n21273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_583_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_583_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_583_LC_13_22_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_583_LC_13_22_2  (
            .in0(N__38247),
            .in1(N__38927),
            .in2(N__42519),
            .in3(N__39594),
            .lcout(\c0.n11432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_877_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_877_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_877_LC_13_22_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_877_LC_13_22_3  (
            .in0(N__42479),
            .in1(N__38926),
            .in2(N__39598),
            .in3(N__38246),
            .lcout(\c0.n63_adj_3146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_390_Select_2_i6_3_lut_4_lut_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.select_390_Select_2_i6_3_lut_4_lut_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_390_Select_2_i6_3_lut_4_lut_LC_13_22_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.select_390_Select_2_i6_3_lut_4_lut_LC_13_22_5  (
            .in0(N__42324),
            .in1(N__34727),
            .in2(N__42507),
            .in3(N__35209),
            .lcout(),
            .ltout(\c0.n6_adj_3521_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_13_22_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_13_22_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_13_22_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_13_22_6  (
            .in0(N__34758),
            .in1(N__31585),
            .in2(N__31579),
            .in3(N__31696),
            .lcout(FRAME_MATCHER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71065),
            .ce(),
            .sr(N__46738));
    defparam \c0.i1_3_lut_4_lut_adj_913_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_913_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_913_LC_13_23_2 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_913_LC_13_23_2  (
            .in0(N__42329),
            .in1(N__38284),
            .in2(N__31576),
            .in3(N__38321),
            .lcout(\c0.n11_adj_3370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_254_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_254_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_254_LC_13_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_254_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__31662),
            .in2(_gnd_net_),
            .in3(N__41434),
            .lcout(\c0.n18657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_797_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_797_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_797_LC_13_23_5 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_797_LC_13_23_5  (
            .in0(N__35155),
            .in1(N__34951),
            .in2(N__35134),
            .in3(N__35207),
            .lcout(),
            .ltout(\c0.n6_adj_3515_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_753_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_753_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_753_LC_13_23_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \c0.i1_4_lut_adj_753_LC_13_23_6  (
            .in0(N__38476),
            .in1(N__31708),
            .in2(N__31699),
            .in3(N__38524),
            .lcout(\c0.n5_adj_3516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_13_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__40490),
            .in2(_gnd_net_),
            .in3(N__34931),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71089),
            .ce(),
            .sr(N__35218));
    defparam \c0.FRAME_MATCHER_state_i5_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_13_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_13_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__31689),
            .in2(_gnd_net_),
            .in3(N__40515),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71105),
            .ce(),
            .sr(N__31672));
    defparam \c0.FRAME_MATCHER_state_i17_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_13_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_13_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__40546),
            .in2(_gnd_net_),
            .in3(N__31658),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71119),
            .ce(),
            .sr(N__31636));
    defparam \c0.FRAME_MATCHER_state_i8_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_13_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_13_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__35471),
            .in2(_gnd_net_),
            .in3(N__40547),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71135),
            .ce(),
            .sr(N__35449));
    defparam \c0.i1_2_lut_adj_860_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_860_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_860_LC_13_28_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_860_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(N__31625),
            .in2(_gnd_net_),
            .in3(N__41466),
            .lcout(\c0.n18629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_2_lut_LC_14_5_0 .C_ON=1'b1;
    defparam \c0.add_80_2_lut_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_2_lut_LC_14_5_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_80_2_lut_LC_14_5_0  (
            .in0(N__42170),
            .in1(N__60208),
            .in2(N__41829),
            .in3(_gnd_net_),
            .lcout(n16),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\c0.n17176 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i1_LC_14_5_1 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i1_LC_14_5_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_14_5_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_14_5_1  (
            .in0(N__42196),
            .in1(N__60041),
            .in2(_gnd_net_),
            .in3(N__31597),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(\c0.n17176 ),
            .carryout(\c0.n17177 ),
            .clk(N__71177),
            .ce(),
            .sr(N__60511));
    defparam \c0.add_80_4_lut_LC_14_5_2 .C_ON=1'b1;
    defparam \c0.add_80_4_lut_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_4_lut_LC_14_5_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_80_4_lut_LC_14_5_2  (
            .in0(N__42171),
            .in1(N__59927),
            .in2(_gnd_net_),
            .in3(N__31726),
            .lcout(\c0.n2_adj_3144 ),
            .ltout(),
            .carryin(\c0.n17177 ),
            .carryout(\c0.n17178 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_5_lut_LC_14_5_3 .C_ON=1'b1;
    defparam \c0.add_80_5_lut_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_5_lut_LC_14_5_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_80_5_lut_LC_14_5_3  (
            .in0(N__42195),
            .in1(N__40062),
            .in2(_gnd_net_),
            .in3(N__31717),
            .lcout(\c0.n2_adj_3145 ),
            .ltout(),
            .carryin(\c0.n17178 ),
            .carryout(\c0.n17179 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_6_lut_LC_14_5_4 .C_ON=1'b1;
    defparam \c0.add_80_6_lut_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_6_lut_LC_14_5_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_80_6_lut_LC_14_5_4  (
            .in0(N__42169),
            .in1(N__40266),
            .in2(_gnd_net_),
            .in3(N__31714),
            .lcout(\c0.n2_adj_3147 ),
            .ltout(),
            .carryin(\c0.n17179 ),
            .carryout(\c0.n17180 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_6_THRU_CRY_0_LC_14_5_5 .C_ON=1'b1;
    defparam \c0.add_80_6_THRU_CRY_0_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_6_THRU_CRY_0_LC_14_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_6_THRU_CRY_0_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__32614),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17180 ),
            .carryout(\c0.n17180_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_6_THRU_CRY_1_LC_14_5_6 .C_ON=1'b1;
    defparam \c0.add_80_6_THRU_CRY_1_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_6_THRU_CRY_1_LC_14_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_6_THRU_CRY_1_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32704),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17180_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17180_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_6_THRU_CRY_2_LC_14_5_7 .C_ON=1'b1;
    defparam \c0.add_80_6_THRU_CRY_2_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_6_THRU_CRY_2_LC_14_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_6_THRU_CRY_2_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__32618),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17180_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17180_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_14_6_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i5_LC_14_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_14_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_14_6_0  (
            .in0(N__42197),
            .in1(N__49618),
            .in2(_gnd_net_),
            .in3(N__31711),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\c0.n17181 ),
            .clk(N__71165),
            .ce(),
            .sr(N__49597));
    defparam \c0.add_80_7_THRU_CRY_0_LC_14_6_1 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_0_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_0_LC_14_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_0_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__32601),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181 ),
            .carryout(\c0.n17181_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_1_LC_14_6_2 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_1_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_1_LC_14_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_1_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_2_LC_14_6_3 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_2_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_2_LC_14_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_2_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__32605),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_3_LC_14_6_4 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_3_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_3_LC_14_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_3_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32702),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_4_LC_14_6_5 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_4_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_4_LC_14_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_4_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__32609),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_5_LC_14_6_6 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_5_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_5_LC_14_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_5_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32703),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_7_THRU_CRY_6_LC_14_6_7 .C_ON=1'b1;
    defparam \c0.add_80_7_THRU_CRY_6_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_7_THRU_CRY_6_LC_14_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_7_THRU_CRY_6_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__32613),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17181_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17181_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_14_7_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i6_LC_14_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_14_7_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_14_7_0  (
            .in0(N__42200),
            .in1(N__40164),
            .in2(_gnd_net_),
            .in3(N__31729),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\c0.n17182 ),
            .clk(N__71152),
            .ce(),
            .sr(N__35803));
    defparam \c0.add_80_8_THRU_CRY_0_LC_14_7_1 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_0_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_0_LC_14_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_0_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__32588),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182 ),
            .carryout(\c0.n17182_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_1_LC_14_7_2 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_1_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_1_LC_14_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_1_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32698),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_2_LC_14_7_3 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_2_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_2_LC_14_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_2_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__32592),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_3_LC_14_7_4 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_3_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_3_LC_14_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_3_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32699),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_4_LC_14_7_5 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_4_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_4_LC_14_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_4_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__32596),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_5_LC_14_7_6 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_5_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_5_LC_14_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_5_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32700),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_8_THRU_CRY_6_LC_14_7_7 .C_ON=1'b1;
    defparam \c0.add_80_8_THRU_CRY_6_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_8_THRU_CRY_6_LC_14_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_8_THRU_CRY_6_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__32600),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17182_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17182_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_14_8_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i7_LC_14_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_14_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_14_8_0  (
            .in0(N__42199),
            .in1(N__34424),
            .in2(_gnd_net_),
            .in3(N__31732),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\c0.n17183 ),
            .clk(N__71138),
            .ce(),
            .sr(N__33481));
    defparam \c0.add_80_9_THRU_CRY_0_LC_14_8_1 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_0_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_0_LC_14_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_0_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__32566),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183 ),
            .carryout(\c0.n17183_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_1_LC_14_8_2 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_1_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_1_LC_14_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_1_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32695),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_2_LC_14_8_3 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_2_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_2_LC_14_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_2_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__32570),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_3_LC_14_8_4 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_3_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_3_LC_14_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_3_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32696),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_4_LC_14_8_5 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_4_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_4_LC_14_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_4_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__32574),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_5_LC_14_8_6 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_5_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_5_LC_14_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_5_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32697),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_9_THRU_CRY_6_LC_14_8_7 .C_ON=1'b1;
    defparam \c0.add_80_9_THRU_CRY_6_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_9_THRU_CRY_6_LC_14_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_9_THRU_CRY_6_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__32578),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17183_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17183_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i8_LC_14_9_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i8_LC_14_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_14_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_14_9_0  (
            .in0(N__42198),
            .in1(N__34610),
            .in2(_gnd_net_),
            .in3(N__31735),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\c0.n17184 ),
            .clk(N__71122),
            .ce(),
            .sr(N__32773));
    defparam \c0.add_80_10_THRU_CRY_0_LC_14_9_1 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_0_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_0_LC_14_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_0_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__32408),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184 ),
            .carryout(\c0.n17184_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_1_LC_14_9_2 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_1_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_1_LC_14_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_1_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_2_LC_14_9_3 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_2_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_2_LC_14_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_2_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__32412),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_3_LC_14_9_4 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_3_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_3_LC_14_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_3_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_4_LC_14_9_5 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_4_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_4_LC_14_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_4_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__32416),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_5_LC_14_9_6 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_5_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_5_LC_14_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_5_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_10_THRU_CRY_6_LC_14_9_7 .C_ON=1'b1;
    defparam \c0.add_80_10_THRU_CRY_6_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_10_THRU_CRY_6_LC_14_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_10_THRU_CRY_6_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__32420),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17184_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17184_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_14_10_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i9_LC_14_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_14_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_14_10_0  (
            .in0(N__42224),
            .in1(N__34802),
            .in2(_gnd_net_),
            .in3(N__31738),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\c0.n17185 ),
            .clk(N__71106),
            .ce(),
            .sr(N__31885));
    defparam \c0.add_80_11_THRU_CRY_0_LC_14_10_1 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_0_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_0_LC_14_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_0_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__32395),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185 ),
            .carryout(\c0.n17185_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_1_LC_14_10_2 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_1_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_1_LC_14_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_1_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_2_LC_14_10_3 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_2_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_2_LC_14_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_2_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__32399),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_3_LC_14_10_4 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_3_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_3_LC_14_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_3_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32583),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_4_LC_14_10_5 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_4_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_4_LC_14_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_4_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__32403),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_5_LC_14_10_6 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_5_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_5_LC_14_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_5_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_11_THRU_CRY_6_LC_14_10_7 .C_ON=1'b1;
    defparam \c0.add_80_11_THRU_CRY_6_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_11_THRU_CRY_6_LC_14_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_11_THRU_CRY_6_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__32407),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17185_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17185_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_14_11_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i10_LC_14_11_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_14_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_14_11_0  (
            .in0(N__42227),
            .in1(N__34892),
            .in2(_gnd_net_),
            .in3(N__31744),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\c0.n17186 ),
            .clk(N__71090),
            .ce(),
            .sr(N__33400));
    defparam \c0.add_80_12_THRU_CRY_0_LC_14_11_1 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_0_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_0_LC_14_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_0_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__32382),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186 ),
            .carryout(\c0.n17186_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_1_LC_14_11_2 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_1_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_1_LC_14_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_1_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_2_LC_14_11_3 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_2_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_2_LC_14_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_2_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__32386),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_3_LC_14_11_4 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_3_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_3_LC_14_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_3_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_4_LC_14_11_5 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_4_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_4_LC_14_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_4_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__32390),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_5_LC_14_11_6 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_5_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_5_LC_14_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_5_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32581),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_12_THRU_CRY_6_LC_14_11_7 .C_ON=1'b1;
    defparam \c0.add_80_12_THRU_CRY_6_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_12_THRU_CRY_6_LC_14_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_12_THRU_CRY_6_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__32394),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17186_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17186_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_14_12_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i11_LC_14_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_14_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_14_12_0  (
            .in0(N__42226),
            .in1(N__34323),
            .in2(_gnd_net_),
            .in3(N__31741),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\c0.n17187 ),
            .clk(N__71078),
            .ce(),
            .sr(N__34405));
    defparam \c0.add_80_13_THRU_CRY_0_LC_14_12_1 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_0_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_0_LC_14_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_0_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__32348),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187 ),
            .carryout(\c0.n17187_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_1_LC_14_12_2 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_1_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_1_LC_14_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_1_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32563),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_2_LC_14_12_3 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_2_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_2_LC_14_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_2_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__32352),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_3_LC_14_12_4 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_3_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_3_LC_14_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_3_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_4_LC_14_12_5 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_4_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_4_LC_14_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_4_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__32356),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_5_LC_14_12_6 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_5_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_5_LC_14_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_5_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32565),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_13_THRU_CRY_6_LC_14_12_7 .C_ON=1'b1;
    defparam \c0.add_80_13_THRU_CRY_6_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_13_THRU_CRY_6_LC_14_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_13_THRU_CRY_6_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__32360),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17187_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17187_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_14_13_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i12_LC_14_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_14_13_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_14_13_0  (
            .in0(N__42225),
            .in1(N__34497),
            .in2(_gnd_net_),
            .in3(N__31747),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\c0.n17188 ),
            .clk(N__71066),
            .ce(),
            .sr(N__34573));
    defparam \c0.add_80_14_THRU_CRY_0_LC_14_13_1 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_0_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_0_LC_14_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_0_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__32193),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188 ),
            .carryout(\c0.n17188_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_1_LC_14_13_2 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_1_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_1_LC_14_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_1_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32379),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_2_LC_14_13_3 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_2_LC_14_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_2_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__32197),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_3_LC_14_13_4 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_3_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_3_LC_14_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_3_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32380),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_4_LC_14_13_5 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_4_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_4_LC_14_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_4_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__32201),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_5_LC_14_13_6 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_5_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_5_LC_14_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_5_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32381),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_14_THRU_CRY_6_LC_14_13_7 .C_ON=1'b1;
    defparam \c0.add_80_14_THRU_CRY_6_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_14_THRU_CRY_6_LC_14_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_14_THRU_CRY_6_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__32205),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17188_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17188_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i13_LC_14_14_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i13_LC_14_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_14_14_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_14_14_0  (
            .in0(N__42249),
            .in1(N__34835),
            .in2(_gnd_net_),
            .in3(N__31762),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\c0.n17189 ),
            .clk(N__71053),
            .ce(),
            .sr(N__31759));
    defparam \c0.add_80_15_THRU_CRY_0_LC_14_14_1 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_0_LC_14_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_0_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__32180),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189 ),
            .carryout(\c0.n17189_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_1_LC_14_14_2 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_1_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_1_LC_14_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_1_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32376),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_2_LC_14_14_3 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_2_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_2_LC_14_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_2_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__32184),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_3_LC_14_14_4 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_3_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_3_LC_14_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_3_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32377),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_4_LC_14_14_5 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_4_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_4_LC_14_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_4_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__32188),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_5_LC_14_14_6 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_5_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_5_LC_14_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_5_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_15_THRU_CRY_6_LC_14_14_7 .C_ON=1'b1;
    defparam \c0.add_80_15_THRU_CRY_6_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_15_THRU_CRY_6_LC_14_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_15_THRU_CRY_6_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__32192),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17189_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17189_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i14_LC_14_15_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i14_LC_14_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_14_15_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_14_15_0  (
            .in0(N__42252),
            .in1(N__34455),
            .in2(_gnd_net_),
            .in3(N__31765),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\c0.n17190 ),
            .clk(N__71041),
            .ce(),
            .sr(N__34522));
    defparam \c0.add_80_16_THRU_CRY_0_LC_14_15_1 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_0_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_0_LC_14_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_0_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__32000),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190 ),
            .carryout(\c0.n17190_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_1_LC_14_15_2 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_1_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_1_LC_14_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_1_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32071),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_2_LC_14_15_3 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_2_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_2_LC_14_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_2_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__32004),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_3_LC_14_15_4 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_3_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_3_LC_14_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_3_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32072),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_4_LC_14_15_5 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_4_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_4_LC_14_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_4_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__32008),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_5_LC_14_15_6 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_5_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_5_LC_14_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_5_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__32073),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_16_THRU_CRY_6_LC_14_15_7 .C_ON=1'b1;
    defparam \c0.add_80_16_THRU_CRY_6_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_16_THRU_CRY_6_LC_14_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_16_THRU_CRY_6_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__32012),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17190_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17190_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_14_16_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i15_LC_14_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_14_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_14_16_0  (
            .in0(N__42251),
            .in1(N__34868),
            .in2(_gnd_net_),
            .in3(N__31768),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\c0.n17191 ),
            .clk(N__71032),
            .ce(),
            .sr(N__33712));
    defparam \c0.add_80_17_THRU_CRY_0_LC_14_16_1 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_0_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_0_LC_14_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_0_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__31993),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191 ),
            .carryout(\c0.n17191_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_1_LC_14_16_2 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_1_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_1_LC_14_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_1_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__31997),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_2_LC_14_16_3 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_2_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_2_LC_14_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_2_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__31994),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_3_LC_14_16_4 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_3_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_3_LC_14_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_3_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__31998),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_4_LC_14_16_5 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_4_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_4_LC_14_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_4_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__31995),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_5_LC_14_16_6 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_5_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_5_LC_14_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_5_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__31999),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_17_THRU_CRY_6_LC_14_16_7 .C_ON=1'b1;
    defparam \c0.add_80_17_THRU_CRY_6_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_17_THRU_CRY_6_LC_14_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_17_THRU_CRY_6_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__31996),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17191_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17191_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_14_17_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i16_LC_14_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_14_17_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_14_17_0  (
            .in0(N__42250),
            .in1(N__34355),
            .in2(_gnd_net_),
            .in3(N__31771),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\c0.n17192 ),
            .clk(N__71015),
            .ce(),
            .sr(N__33655));
    defparam \c0.add_80_18_THRU_CRY_0_LC_14_17_1 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_0_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_0_LC_14_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_0_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__32013),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192 ),
            .carryout(\c0.n17192_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_1_LC_14_17_2 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_1_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_1_LC_14_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_1_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__32017),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_2_LC_14_17_3 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_2_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_2_LC_14_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_2_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__32014),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_3_LC_14_17_4 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_3_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_3_LC_14_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_3_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__32018),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_4_LC_14_17_5 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_4_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_4_LC_14_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_4_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__32015),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_5_LC_14_17_6 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_5_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_5_LC_14_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_5_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__32019),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_18_THRU_CRY_6_LC_14_17_7 .C_ON=1'b1;
    defparam \c0.add_80_18_THRU_CRY_6_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_18_THRU_CRY_6_LC_14_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_18_THRU_CRY_6_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__32016),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17192_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17192_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i17_LC_14_18_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i17_LC_14_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_14_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_14_18_0  (
            .in0(N__42265),
            .in1(N__35042),
            .in2(_gnd_net_),
            .in3(N__31786),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\c0.n17193 ),
            .clk(N__71033),
            .ce(),
            .sr(N__31783));
    defparam \c0.add_80_19_THRU_CRY_0_LC_14_18_1 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_0_LC_14_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__32148),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193 ),
            .carryout(\c0.n17193_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_1_LC_14_18_2 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_1_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_1_LC_14_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_1_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__32152),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_2_LC_14_18_3 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_2_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_2_LC_14_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_2_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__32149),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_3_LC_14_18_4 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_3_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_3_LC_14_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_3_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__32153),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_4_LC_14_18_5 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_4_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_4_LC_14_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_4_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__32150),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_5_LC_14_18_6 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_5_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_5_LC_14_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_5_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__32154),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_19_THRU_CRY_6_LC_14_18_7 .C_ON=1'b1;
    defparam \c0.add_80_19_THRU_CRY_6_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_19_THRU_CRY_6_LC_14_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_19_THRU_CRY_6_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__32151),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17193_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17193_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_14_19_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i18_LC_14_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_14_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_14_19_0  (
            .in0(N__42266),
            .in1(N__38045),
            .in2(_gnd_net_),
            .in3(N__31798),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\c0.n17194 ),
            .clk(N__71042),
            .ce(),
            .sr(N__31795));
    defparam \c0.add_80_20_THRU_CRY_0_LC_14_19_1 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_0_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_0_LC_14_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_0_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__32155),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194 ),
            .carryout(\c0.n17194_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_1_LC_14_19_2 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_1_LC_14_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_1_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__32159),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_2_LC_14_19_3 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_2_LC_14_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_2_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__32156),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_3_LC_14_19_4 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_3_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_3_LC_14_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_3_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__32160),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_4_LC_14_19_5 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_4_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_4_LC_14_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_4_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__32157),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_5_LC_14_19_6 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_5_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_5_LC_14_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_5_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__32161),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_20_THRU_CRY_6_LC_14_19_7 .C_ON=1'b1;
    defparam \c0.add_80_20_THRU_CRY_6_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_20_THRU_CRY_6_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_20_THRU_CRY_6_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__32158),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17194_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17194_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i19_LC_14_20_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i19_LC_14_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_14_20_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_14_20_0  (
            .in0(N__42268),
            .in1(N__34589),
            .in2(_gnd_net_),
            .in3(N__31816),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\c0.n17195 ),
            .clk(N__71054),
            .ce(),
            .sr(N__31813));
    defparam \c0.add_80_21_THRU_CRY_0_LC_14_20_1 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_0_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_0_LC_14_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_0_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__32258),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195 ),
            .carryout(\c0.n17195_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_1_LC_14_20_2 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_1_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_1_LC_14_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_1_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__32262),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_2_LC_14_20_3 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_2_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_2_LC_14_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_2_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__32259),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_3_LC_14_20_4 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_3_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_3_LC_14_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_3_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__32263),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_4_LC_14_20_5 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_4_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_4_LC_14_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_4_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__32260),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_5_LC_14_20_6 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_5_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_5_LC_14_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_5_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__32264),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_21_THRU_CRY_6_LC_14_20_7 .C_ON=1'b1;
    defparam \c0.add_80_21_THRU_CRY_6_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_21_THRU_CRY_6_LC_14_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_21_THRU_CRY_6_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__32261),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17195_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17195_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i20_LC_14_21_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i20_LC_14_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_14_21_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_14_21_0  (
            .in0(N__42267),
            .in1(N__34482),
            .in2(_gnd_net_),
            .in3(N__31801),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\c0.n17196 ),
            .clk(N__71067),
            .ce(),
            .sr(N__31834));
    defparam \c0.add_80_22_THRU_CRY_0_LC_14_21_1 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_0_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_0_LC_14_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_0_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__32458),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196 ),
            .carryout(\c0.n17196_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_1_LC_14_21_2 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_1_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_1_LC_14_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_1_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__32462),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_2_LC_14_21_3 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_2_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_2_LC_14_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_2_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__32459),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_3_LC_14_21_4 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_3_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_3_LC_14_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_3_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__32463),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_4_LC_14_21_5 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_4_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_4_LC_14_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_4_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__32460),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_5_LC_14_21_6 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_5_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_5_LC_14_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_5_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__32464),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_22_THRU_CRY_6_LC_14_21_7 .C_ON=1'b1;
    defparam \c0.add_80_22_THRU_CRY_6_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_22_THRU_CRY_6_LC_14_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_22_THRU_CRY_6_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__32461),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17196_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17196_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i21_LC_14_22_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i21_LC_14_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_14_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_14_22_0  (
            .in0(N__42140),
            .in1(N__35078),
            .in2(_gnd_net_),
            .in3(N__31828),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\c0.n17197 ),
            .clk(N__71079),
            .ce(),
            .sr(N__31825));
    defparam \c0.add_80_23_THRU_CRY_0_LC_14_22_1 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_0_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_0_LC_14_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_0_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__32465),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197 ),
            .carryout(\c0.n17197_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_1_LC_14_22_2 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_1_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_1_LC_14_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_1_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__32469),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_2_LC_14_22_3 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_2_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_2_LC_14_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_2_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__32466),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_3_LC_14_22_4 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_3_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_3_LC_14_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_3_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__32470),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_4_LC_14_22_5 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_4_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_4_LC_14_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_4_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__32467),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_5_LC_14_22_6 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_5_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_5_LC_14_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_5_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__32471),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_23_THRU_CRY_6_LC_14_22_7 .C_ON=1'b1;
    defparam \c0.add_80_23_THRU_CRY_6_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_23_THRU_CRY_6_LC_14_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_23_THRU_CRY_6_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__32468),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17197_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17197_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i22_LC_14_23_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i22_LC_14_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_14_23_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_14_23_0  (
            .in0(N__42145),
            .in1(N__34382),
            .in2(_gnd_net_),
            .in3(N__31849),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\c0.n17198 ),
            .clk(N__71091),
            .ce(),
            .sr(N__31846));
    defparam \c0.add_80_24_THRU_CRY_0_LC_14_23_1 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_0_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_0_LC_14_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_0_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__32472),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198 ),
            .carryout(\c0.n17198_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_1_LC_14_23_2 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_1_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_1_LC_14_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_1_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__32476),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_2_LC_14_23_3 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_2_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_2_LC_14_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_2_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__32473),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_3_LC_14_23_4 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_3_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_3_LC_14_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_3_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__32477),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_4_LC_14_23_5 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_4_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_4_LC_14_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_4_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__32474),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_5_LC_14_23_6 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_5_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_5_LC_14_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_5_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__32478),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_24_THRU_CRY_6_LC_14_23_7 .C_ON=1'b1;
    defparam \c0.add_80_24_THRU_CRY_6_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_24_THRU_CRY_6_LC_14_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_24_THRU_CRY_6_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__32475),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17198_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17198_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i23_LC_14_24_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i23_LC_14_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_14_24_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_14_24_0  (
            .in0(N__42141),
            .in1(N__38018),
            .in2(_gnd_net_),
            .in3(N__31852),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\c0.n17199 ),
            .clk(N__71107),
            .ce(),
            .sr(N__35164));
    defparam \c0.add_80_25_THRU_CRY_0_LC_14_24_1 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_0_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_0_LC_14_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_0_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__32479),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199 ),
            .carryout(\c0.n17199_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_1_LC_14_24_2 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_1_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_1_LC_14_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_1_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__32483),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_2_LC_14_24_3 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_2_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_2_LC_14_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_2_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__32480),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_3_LC_14_24_4 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_3_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_3_LC_14_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_3_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__32484),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_4_LC_14_24_5 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_4_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_4_LC_14_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_4_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__32481),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_5_LC_14_24_6 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_5_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_5_LC_14_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_5_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__32485),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_25_THRU_CRY_6_LC_14_24_7 .C_ON=1'b1;
    defparam \c0.add_80_25_THRU_CRY_6_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_25_THRU_CRY_6_LC_14_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_25_THRU_CRY_6_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__32482),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17199_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17199_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i24_LC_14_25_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i24_LC_14_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_14_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_14_25_0  (
            .in0(N__42127),
            .in1(N__35013),
            .in2(_gnd_net_),
            .in3(N__31855),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\c0.n17200 ),
            .clk(N__71121),
            .ce(),
            .sr(N__34996));
    defparam \c0.add_80_26_THRU_CRY_0_LC_14_25_1 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_0_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_0_LC_14_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_0_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__32619),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200 ),
            .carryout(\c0.n17200_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_1_LC_14_25_2 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_1_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_1_LC_14_25_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_1_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__32623),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_2_LC_14_25_3 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_2_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_2_LC_14_25_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_2_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__32620),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_3_LC_14_25_4 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_3_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_3_LC_14_25_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_3_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__32624),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_4_LC_14_25_5 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_4_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_4_LC_14_25_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_4_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__32621),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_5_LC_14_25_6 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_5_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_5_LC_14_25_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_5_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__32625),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_26_THRU_CRY_6_LC_14_25_7 .C_ON=1'b1;
    defparam \c0.add_80_26_THRU_CRY_6_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_26_THRU_CRY_6_LC_14_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_26_THRU_CRY_6_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__32622),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17200_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17200_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_14_26_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i25_LC_14_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_14_26_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_14_26_0  (
            .in0(N__42142),
            .in1(N__34551),
            .in2(_gnd_net_),
            .in3(N__31858),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\c0.n17201 ),
            .clk(N__71137),
            .ce(),
            .sr(N__34537));
    defparam \c0.add_80_27_THRU_CRY_0_LC_14_26_1 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_0_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_0_LC_14_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_0_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__32626),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201 ),
            .carryout(\c0.n17201_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_1_LC_14_26_2 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_1_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_1_LC_14_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_1_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__32630),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_2_LC_14_26_3 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_2_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_2_LC_14_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_2_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__32627),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_3_LC_14_26_4 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_3_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_3_LC_14_26_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_3_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__32631),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_4_LC_14_26_5 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_4_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_4_LC_14_26_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_4_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__32628),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_5_LC_14_26_6 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_5_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_5_LC_14_26_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_5_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__32632),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_27_THRU_CRY_6_LC_14_26_7 .C_ON=1'b1;
    defparam \c0.add_80_27_THRU_CRY_6_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_27_THRU_CRY_6_LC_14_26_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_27_THRU_CRY_6_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(N__32629),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17201_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17201_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i26_LC_14_27_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i26_LC_14_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_14_27_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_14_27_0  (
            .in0(N__42143),
            .in1(N__35375),
            .in2(_gnd_net_),
            .in3(N__31861),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\c0.n17202 ),
            .clk(N__71151),
            .ce(),
            .sr(N__35353));
    defparam \c0.add_80_28_THRU_CRY_0_LC_14_27_1 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_0_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_0_LC_14_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_0_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__32633),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202 ),
            .carryout(\c0.n17202_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_1_LC_14_27_2 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_1_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_1_LC_14_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_1_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(N__32637),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_2_LC_14_27_3 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_2_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_2_LC_14_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_2_LC_14_27_3  (
            .in0(_gnd_net_),
            .in1(N__32634),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_3_LC_14_27_4 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_3_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_3_LC_14_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_3_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__32638),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_4_LC_14_27_5 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_4_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_4_LC_14_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_4_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(N__32635),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_5_LC_14_27_6 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_5_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_5_LC_14_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_5_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(N__32639),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_28_THRU_CRY_6_LC_14_27_7 .C_ON=1'b1;
    defparam \c0.add_80_28_THRU_CRY_6_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_28_THRU_CRY_6_LC_14_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_28_THRU_CRY_6_LC_14_27_7  (
            .in0(_gnd_net_),
            .in1(N__32636),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17202_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17202_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i27_LC_14_28_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i27_LC_14_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_14_28_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_14_28_0  (
            .in0(N__42125),
            .in1(N__35327),
            .in2(_gnd_net_),
            .in3(N__31864),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(\c0.n17203 ),
            .clk(N__71164),
            .ce(),
            .sr(N__35308));
    defparam \c0.add_80_29_THRU_CRY_0_LC_14_28_1 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_0_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_0_LC_14_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_0_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(N__32640),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203 ),
            .carryout(\c0.n17203_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_1_LC_14_28_2 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_1_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_1_LC_14_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_1_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__32644),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_2_LC_14_28_3 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_2_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_2_LC_14_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_2_LC_14_28_3  (
            .in0(_gnd_net_),
            .in1(N__32641),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_3_LC_14_28_4 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_3_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_3_LC_14_28_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_3_LC_14_28_4  (
            .in0(_gnd_net_),
            .in1(N__32645),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_4_LC_14_28_5 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_4_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_4_LC_14_28_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_4_LC_14_28_5  (
            .in0(_gnd_net_),
            .in1(N__32642),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_5_LC_14_28_6 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_5_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_5_LC_14_28_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_5_LC_14_28_6  (
            .in0(_gnd_net_),
            .in1(N__32646),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_29_THRU_CRY_6_LC_14_28_7 .C_ON=1'b1;
    defparam \c0.add_80_29_THRU_CRY_6_LC_14_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_29_THRU_CRY_6_LC_14_28_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_29_THRU_CRY_6_LC_14_28_7  (
            .in0(_gnd_net_),
            .in1(N__32643),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17203_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17203_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i28_LC_14_29_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i28_LC_14_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_14_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_14_29_0  (
            .in0(N__42126),
            .in1(N__35291),
            .in2(_gnd_net_),
            .in3(N__31870),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(bfn_14_29_0_),
            .carryout(\c0.n17204 ),
            .clk(N__71176),
            .ce(),
            .sr(N__35272));
    defparam \c0.add_80_30_THRU_CRY_0_LC_14_29_1 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_0_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_0_LC_14_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_0_LC_14_29_1  (
            .in0(_gnd_net_),
            .in1(N__32705),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204 ),
            .carryout(\c0.n17204_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_1_LC_14_29_2 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_1_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_1_LC_14_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_1_LC_14_29_2  (
            .in0(_gnd_net_),
            .in1(N__32709),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_2_LC_14_29_3 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_2_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_2_LC_14_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_2_LC_14_29_3  (
            .in0(_gnd_net_),
            .in1(N__32706),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_3_LC_14_29_4 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_3_LC_14_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_3_LC_14_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_3_LC_14_29_4  (
            .in0(_gnd_net_),
            .in1(N__32710),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_4_LC_14_29_5 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_4_LC_14_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_4_LC_14_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_4_LC_14_29_5  (
            .in0(_gnd_net_),
            .in1(N__32707),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_5_LC_14_29_6 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_5_LC_14_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_5_LC_14_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_5_LC_14_29_6  (
            .in0(_gnd_net_),
            .in1(N__32711),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_30_THRU_CRY_6_LC_14_29_7 .C_ON=1'b1;
    defparam \c0.add_80_30_THRU_CRY_6_LC_14_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_30_THRU_CRY_6_LC_14_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_30_THRU_CRY_6_LC_14_29_7  (
            .in0(_gnd_net_),
            .in1(N__32708),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17204_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17204_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i29_LC_14_30_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i29_LC_14_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_14_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_14_30_0  (
            .in0(N__42131),
            .in1(N__37985),
            .in2(_gnd_net_),
            .in3(N__31867),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(bfn_14_30_0_),
            .carryout(\c0.n17205 ),
            .clk(N__71188),
            .ce(),
            .sr(N__35344));
    defparam \c0.add_80_31_THRU_CRY_0_LC_14_30_1 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_0_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_0_LC_14_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_0_LC_14_30_1  (
            .in0(_gnd_net_),
            .in1(N__32712),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205 ),
            .carryout(\c0.n17205_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_1_LC_14_30_2 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_1_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_1_LC_14_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_1_LC_14_30_2  (
            .in0(_gnd_net_),
            .in1(N__32716),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_2_LC_14_30_3 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_2_LC_14_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_2_LC_14_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_2_LC_14_30_3  (
            .in0(_gnd_net_),
            .in1(N__32713),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_3_LC_14_30_4 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_3_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_3_LC_14_30_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_3_LC_14_30_4  (
            .in0(_gnd_net_),
            .in1(N__32717),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_4_LC_14_30_5 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_4_LC_14_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_4_LC_14_30_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_4_LC_14_30_5  (
            .in0(_gnd_net_),
            .in1(N__32714),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_5_LC_14_30_6 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_5_LC_14_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_5_LC_14_30_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_5_LC_14_30_6  (
            .in0(_gnd_net_),
            .in1(N__32718),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_31_THRU_CRY_6_LC_14_30_7 .C_ON=1'b1;
    defparam \c0.add_80_31_THRU_CRY_6_LC_14_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_31_THRU_CRY_6_LC_14_30_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_31_THRU_CRY_6_LC_14_30_7  (
            .in0(_gnd_net_),
            .in1(N__32715),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17205_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17205_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i30_LC_14_31_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i30_LC_14_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_14_31_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_14_31_0  (
            .in0(N__42121),
            .in1(N__35246),
            .in2(_gnd_net_),
            .in3(N__31873),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(bfn_14_31_0_),
            .carryout(\c0.n17206 ),
            .clk(N__71199),
            .ce(),
            .sr(N__35227));
    defparam \c0.add_80_32_THRU_CRY_0_LC_14_31_1 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_0_LC_14_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_0_LC_14_31_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_0_LC_14_31_1  (
            .in0(_gnd_net_),
            .in1(N__32719),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206 ),
            .carryout(\c0.n17206_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_1_LC_14_31_2 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_1_LC_14_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_1_LC_14_31_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_1_LC_14_31_2  (
            .in0(_gnd_net_),
            .in1(N__32723),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_2_LC_14_31_3 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_2_LC_14_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_2_LC_14_31_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_2_LC_14_31_3  (
            .in0(_gnd_net_),
            .in1(N__32720),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_3_LC_14_31_4 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_3_LC_14_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_3_LC_14_31_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_3_LC_14_31_4  (
            .in0(_gnd_net_),
            .in1(N__32724),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_4_LC_14_31_5 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_4_LC_14_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_4_LC_14_31_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_4_LC_14_31_5  (
            .in0(_gnd_net_),
            .in1(N__32721),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_5_LC_14_31_6 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_5_LC_14_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_5_LC_14_31_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_5_LC_14_31_6  (
            .in0(_gnd_net_),
            .in1(N__32725),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_80_32_THRU_CRY_6_LC_14_31_7 .C_ON=1'b1;
    defparam \c0.add_80_32_THRU_CRY_6_LC_14_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_80_32_THRU_CRY_6_LC_14_31_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_80_32_THRU_CRY_6_LC_14_31_7  (
            .in0(_gnd_net_),
            .in1(N__32722),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n17206_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n17206_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i31_LC_14_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_14_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_14_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_14_32_0  (
            .in0(N__42144),
            .in1(N__38135),
            .in2(_gnd_net_),
            .in3(N__31915),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71212),
            .ce(),
            .sr(N__35263));
    defparam \c0.FRAME_MATCHER_i_i0_LC_15_8_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i0_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_i_i0_LC_15_8_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_15_8_0  (
            .in0(N__60652),
            .in1(N__31912),
            .in2(N__60235),
            .in3(N__31897),
            .lcout(FRAME_MATCHER_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71154),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_9_i6_2_lut_LC_15_8_1 .C_ON=1'b0;
    defparam \c0.select_357_Select_9_i6_2_lut_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_9_i6_2_lut_LC_15_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_9_i6_2_lut_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__34809),
            .in2(_gnd_net_),
            .in3(N__60651),
            .lcout(\c0.n6_adj_3155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__5__5345_LC_15_8_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__5__5345_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__5__5345_LC_15_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_11__5__5345_LC_15_8_3  (
            .in0(N__32964),
            .in1(N__33141),
            .in2(_gnd_net_),
            .in3(N__46692),
            .lcout(data_out_frame_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71154),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__0__5390_LC_15_8_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__0__5390_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__0__5390_LC_15_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_6__0__5390_LC_15_8_4  (
            .in0(N__46691),
            .in1(N__32896),
            .in2(_gnd_net_),
            .in3(N__32763),
            .lcout(data_out_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71154),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i5_LC_15_9_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i5_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i5_LC_15_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i5_LC_15_9_1  (
            .in0(N__36254),
            .in1(N__32843),
            .in2(_gnd_net_),
            .in3(N__32866),
            .lcout(encoder1_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71139),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_9_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_9_2 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_9_2  (
            .in0(N__32781),
            .in1(N__40924),
            .in2(N__33646),
            .in3(N__36758),
            .lcout(\c0.n21647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__2__5356_LC_15_9_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__2__5356_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__2__5356_LC_15_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_10__2__5356_LC_15_9_3  (
            .in0(N__32806),
            .in1(N__32782),
            .in2(_gnd_net_),
            .in3(N__46914),
            .lcout(data_out_frame_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71139),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_8_i6_2_lut_LC_15_9_6 .C_ON=1'b0;
    defparam \c0.select_357_Select_8_i6_2_lut_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_8_i6_2_lut_LC_15_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_8_i6_2_lut_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__60650),
            .in2(_gnd_net_),
            .in3(N__34614),
            .lcout(\c0.n6_adj_3154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__5__5209_LC_15_9_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__5__5209_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__5__5209_LC_15_9_7 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \c0.data_out_frame_28__5__5209_LC_15_9_7  (
            .in0(N__37488),
            .in1(N__62180),
            .in2(N__54479),
            .in3(N__46915),
            .lcout(data_out_frame_28_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71139),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13745_4_lut_LC_15_10_0 .C_ON=1'b0;
    defparam \c0.i13745_4_lut_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13745_4_lut_LC_15_10_0 .LUT_INIT=16'b1010000000001100;
    LogicCell40 \c0.i13745_4_lut_LC_15_10_0  (
            .in0(N__32764),
            .in1(N__40925),
            .in2(N__36987),
            .in3(N__36755),
            .lcout(\c0.n6_adj_3321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i1_LC_15_10_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i1_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i1_LC_15_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i1_LC_15_10_2  (
            .in0(N__33689),
            .in1(N__36226),
            .in2(_gnd_net_),
            .in3(N__32737),
            .lcout(encoder1_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71123),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__4__5210_LC_15_10_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__4__5210_LC_15_10_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__4__5210_LC_15_10_3 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \c0.data_out_frame_28__4__5210_LC_15_10_3  (
            .in0(N__46860),
            .in1(N__62182),
            .in2(N__61132),
            .in3(N__33063),
            .lcout(data_out_frame_28_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71123),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_210_LC_15_10_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_210_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_210_LC_15_10_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_210_LC_15_10_6  (
            .in0(N__37231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39352),
            .lcout(n11461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i3_LC_15_10_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i3_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i3_LC_15_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i3_LC_15_10_7  (
            .in0(N__36225),
            .in1(N__33023),
            .in2(_gnd_net_),
            .in3(N__33049),
            .lcout(encoder1_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71123),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__3__5379_LC_15_11_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__3__5379_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__3__5379_LC_15_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__3__5379_LC_15_11_0  (
            .in0(N__33004),
            .in1(N__35515),
            .in2(_gnd_net_),
            .in3(N__46799),
            .lcout(data_out_frame_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71108),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_15_11_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_15_11_1 .LUT_INIT=16'b1111010101000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_15_11_1  (
            .in0(N__36966),
            .in1(N__33439),
            .in2(N__33088),
            .in3(N__40904),
            .lcout(),
            .ltout(\c0.n6_adj_3379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17727_4_lut_LC_15_11_2 .C_ON=1'b0;
    defparam \c0.i17727_4_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17727_4_lut_LC_15_11_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i17727_4_lut_LC_15_11_2  (
            .in0(N__36731),
            .in1(N__35485),
            .in2(N__32980),
            .in3(N__36967),
            .lcout(\c0.n21314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i21_LC_15_11_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i21_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i21_LC_15_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i21_LC_15_11_3  (
            .in0(N__36249),
            .in1(N__32977),
            .in2(_gnd_net_),
            .in3(N__32957),
            .lcout(encoder1_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71108),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i45_2_lut_LC_15_11_5 .C_ON=1'b0;
    defparam \c0.i45_2_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i45_2_lut_LC_15_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i45_2_lut_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__52996),
            .in2(_gnd_net_),
            .in3(N__38786),
            .lcout(\c0.n160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17733_4_lut_LC_15_11_6 .C_ON=1'b0;
    defparam \c0.i17733_4_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17733_4_lut_LC_15_11_6 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.i17733_4_lut_LC_15_11_6  (
            .in0(N__32938),
            .in1(N__32923),
            .in2(N__36757),
            .in3(N__36968),
            .lcout(\c0.n21320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i23_LC_15_11_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i23_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i23_LC_15_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i23_LC_15_11_7  (
            .in0(N__36250),
            .in1(N__36311),
            .in2(_gnd_net_),
            .in3(N__32911),
            .lcout(encoder1_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71108),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_15_12_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_15_12_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_15_12_0  (
            .in0(N__37810),
            .in1(N__37870),
            .in2(N__53036),
            .in3(N__34273),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71092),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__3__5371_LC_15_12_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__3__5371_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__3__5371_LC_15_12_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame_8__3__5371_LC_15_12_1  (
            .in0(N__46796),
            .in1(_gnd_net_),
            .in2(N__33178),
            .in3(N__33265),
            .lcout(data_out_frame_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71092),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18039_LC_15_12_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18039_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18039_LC_15_12_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18039_LC_15_12_2  (
            .in0(N__36723),
            .in1(N__33235),
            .in2(N__36292),
            .in3(N__40908),
            .lcout(\c0.n21623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21641_bdd_4_lut_LC_15_12_3 .C_ON=1'b0;
    defparam \c0.n21641_bdd_4_lut_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.n21641_bdd_4_lut_LC_15_12_3 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n21641_bdd_4_lut_LC_15_12_3  (
            .in0(N__33205),
            .in1(N__33190),
            .in2(N__33177),
            .in3(N__36726),
            .lcout(\c0.n21644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5165_LC_15_12_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5165_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5165_LC_15_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.FRAME_MATCHER_rx_data_ready_prev_5165_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53011),
            .lcout(\c0.FRAME_MATCHER_rx_data_ready_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71092),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18049_LC_15_12_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18049_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18049_LC_15_12_5 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18049_LC_15_12_5  (
            .in0(N__40907),
            .in1(N__33366),
            .in2(N__33148),
            .in3(N__36724),
            .lcout(),
            .ltout(\c0.n21635_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21635_bdd_4_lut_LC_15_12_6 .C_ON=1'b0;
    defparam \c0.n21635_bdd_4_lut_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.n21635_bdd_4_lut_LC_15_12_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n21635_bdd_4_lut_LC_15_12_6  (
            .in0(N__36725),
            .in1(N__33127),
            .in2(N__33112),
            .in3(N__33109),
            .lcout(\c0.n21638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__3__5395_LC_15_12_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__3__5395_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__3__5395_LC_15_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_5__3__5395_LC_15_12_7  (
            .in0(N__46795),
            .in1(N__38740),
            .in2(_gnd_net_),
            .in3(N__33087),
            .lcout(data_out_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71092),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__3__5211_LC_15_13_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__3__5211_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__3__5211_LC_15_13_1 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \c0.data_out_frame_28__3__5211_LC_15_13_1  (
            .in0(N__61131),
            .in1(N__36019),
            .in2(N__56860),
            .in3(N__46798),
            .lcout(\c0.data_out_frame_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71080),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17910_2_lut_LC_15_13_2 .C_ON=1'b0;
    defparam \c0.i17910_2_lut_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17910_2_lut_LC_15_13_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i17910_2_lut_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__35814),
            .in2(_gnd_net_),
            .in3(N__36736),
            .lcout(\c0.n21470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i179_LC_15_13_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i179_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i179_LC_15_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i179_LC_15_13_3  (
            .in0(N__68612),
            .in1(N__67526),
            .in2(_gnd_net_),
            .in3(N__58871),
            .lcout(data_in_frame_22_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71080),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17955_3_lut_LC_15_13_4 .C_ON=1'b0;
    defparam \c0.i17955_3_lut_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17955_3_lut_LC_15_13_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i17955_3_lut_LC_15_13_4  (
            .in0(N__36048),
            .in1(N__36976),
            .in2(_gnd_net_),
            .in3(N__40900),
            .lcout(\c0.n21542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i29_LC_15_13_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i29_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i29_LC_15_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i29_LC_15_13_5  (
            .in0(N__36227),
            .in1(N__33383),
            .in2(_gnd_net_),
            .in3(N__33412),
            .lcout(encoder1_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71080),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_10_i6_2_lut_LC_15_13_6 .C_ON=1'b0;
    defparam \c0.select_357_Select_10_i6_2_lut_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_10_i6_2_lut_LC_15_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_10_i6_2_lut_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__34896),
            .in2(_gnd_net_),
            .in3(N__60688),
            .lcout(\c0.n6_adj_3156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__5__5353_LC_15_13_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__5__5353_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__5__5353_LC_15_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_10__5__5353_LC_15_13_7  (
            .in0(N__33367),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__46797),
            .lcout(data_out_frame_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71080),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__5__5385_LC_15_14_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__5__5385_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__5__5385_LC_15_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_6__5__5385_LC_15_14_1  (
            .in0(N__46779),
            .in1(N__33355),
            .in2(_gnd_net_),
            .in3(N__33906),
            .lcout(data_out_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71068),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13744_3_lut_LC_15_14_2 .C_ON=1'b0;
    defparam \c0.i13744_3_lut_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13744_3_lut_LC_15_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i13744_3_lut_LC_15_14_2  (
            .in0(N__36727),
            .in1(N__33325),
            .in2(_gnd_net_),
            .in3(N__36459),
            .lcout(\c0.n17150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__2__5348_LC_15_14_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__2__5348_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__2__5348_LC_15_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_11__2__5348_LC_15_14_4  (
            .in0(N__33295),
            .in1(N__33642),
            .in2(_gnd_net_),
            .in3(N__46780),
            .lcout(data_out_frame_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71068),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18034_LC_15_14_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18034_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_18034_LC_15_14_5 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_18034_LC_15_14_5  (
            .in0(N__33627),
            .in1(N__40893),
            .in2(N__33613),
            .in3(N__36728),
            .lcout(),
            .ltout(\c0.n21617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n21617_bdd_4_lut_LC_15_14_6 .C_ON=1'b0;
    defparam \c0.n21617_bdd_4_lut_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.n21617_bdd_4_lut_LC_15_14_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n21617_bdd_4_lut_LC_15_14_6  (
            .in0(N__36729),
            .in1(N__33592),
            .in2(N__33577),
            .in3(N__33574),
            .lcout(),
            .ltout(\c0.n21620_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17986_4_lut_LC_15_14_7 .C_ON=1'b0;
    defparam \c0.i17986_4_lut_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17986_4_lut_LC_15_14_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.i17986_4_lut_LC_15_14_7  (
            .in0(N__36376),
            .in1(N__36950),
            .in2(N__33559),
            .in3(N__36730),
            .lcout(\c0.n21574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_271_LC_15_15_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_271_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_271_LC_15_15_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_271_LC_15_15_0  (
            .in0(N__33879),
            .in1(N__33544),
            .in2(_gnd_net_),
            .in3(N__33526),
            .lcout(\c0.n7235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i4_LC_15_15_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i4_LC_15_15_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_15_15_1 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_15_15_1  (
            .in0(N__38674),
            .in1(N__33496),
            .in2(N__40265),
            .in3(N__60687),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71055),
            .ce(),
            .sr(N__46729));
    defparam \c0.select_357_Select_7_i6_2_lut_LC_15_15_7 .C_ON=1'b0;
    defparam \c0.select_357_Select_7_i6_2_lut_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_7_i6_2_lut_LC_15_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_7_i6_2_lut_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__60686),
            .in2(_gnd_net_),
            .in3(N__34441),
            .lcout(\c0.n6_adj_3151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17721_4_lut_LC_15_16_0 .C_ON=1'b0;
    defparam \c0.i17721_4_lut_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17721_4_lut_LC_15_16_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.i17721_4_lut_LC_15_16_0  (
            .in0(N__36696),
            .in1(N__36959),
            .in2(N__33721),
            .in3(N__33892),
            .lcout(\c0.n21308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__5__5377_LC_15_16_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__5__5377_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__5__5377_LC_15_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_7__5__5377_LC_15_16_1  (
            .in0(N__33916),
            .in1(N__33466),
            .in2(_gnd_net_),
            .in3(N__46888),
            .lcout(data_out_frame_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71043),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_15_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_15_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_15_16_2  (
            .in0(N__40846),
            .in1(N__33946),
            .in2(_gnd_net_),
            .in3(N__43441),
            .lcout(\c0.n5_adj_3475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_15_16_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_16_3 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_15_16_3  (
            .in0(N__37531),
            .in1(N__33930),
            .in2(N__33805),
            .in3(N__33881),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71043),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_15_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_15_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_15_16_4  (
            .in0(N__40845),
            .in1(N__33915),
            .in2(_gnd_net_),
            .in3(N__33907),
            .lcout(\c0.n5_adj_3447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_15_16_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_15_16_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_15_16_6  (
            .in0(N__33880),
            .in1(N__33801),
            .in2(N__34119),
            .in3(N__35926),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71043),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17958_4_lut_LC_15_16_7 .C_ON=1'b0;
    defparam \c0.i17958_4_lut_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17958_4_lut_LC_15_16_7 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \c0.i17958_4_lut_LC_15_16_7  (
            .in0(N__36958),
            .in1(N__40844),
            .in2(N__33742),
            .in3(N__36695),
            .lcout(\c0.n21546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_15_i6_2_lut_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.select_357_Select_15_i6_2_lut_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_15_i6_2_lut_LC_15_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_15_i6_2_lut_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__34869),
            .in2(_gnd_net_),
            .in3(N__60653),
            .lcout(\c0.n6_adj_3192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__1__5333_LC_15_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__1__5333_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__1__5333_LC_15_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_13__1__5333_LC_15_17_1  (
            .in0(N__33703),
            .in1(N__33669),
            .in2(_gnd_net_),
            .in3(N__46642),
            .lcout(data_out_frame_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71026),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_16_i6_2_lut_LC_15_17_2 .C_ON=1'b0;
    defparam \c0.select_357_Select_16_i6_2_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_16_i6_2_lut_LC_15_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_16_i6_2_lut_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__60654),
            .in2(_gnd_net_),
            .in3(N__34356),
            .lcout(\c0.n6_adj_3190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11148_4_lut_3_lut_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.rx.i11148_4_lut_3_lut_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11148_4_lut_3_lut_LC_15_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \c0.rx.i11148_4_lut_3_lut_LC_15_17_3  (
            .in0(N__37920),
            .in1(N__56193),
            .in2(_gnd_net_),
            .in3(N__39231),
            .lcout(),
            .ltout(\c0.rx.n14601_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_15_17_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_15_17_4 .LUT_INIT=16'b0001000001010100;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_15_17_4  (
            .in0(N__37800),
            .in1(N__37858),
            .in2(N__34276),
            .in3(N__37537),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71026),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_4_lut_LC_15_17_5.C_ON=1'b0;
    defparam i13_4_lut_4_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam i13_4_lut_4_lut_LC_15_17_5.LUT_INIT=16'b0010010100000101;
    LogicCell40 i13_4_lut_4_lut_LC_15_17_5 (
            .in0(N__37857),
            .in1(N__37799),
            .in2(N__37929),
            .in3(N__37749),
            .lcout(n12301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12241_2_lut_LC_15_17_7 .C_ON=1'b0;
    defparam \c0.i12241_2_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12241_2_lut_LC_15_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i12241_2_lut_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__40826),
            .in2(_gnd_net_),
            .in3(N__36707),
            .lcout(\c0.n15685 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_15_18_0 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_15_18_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \c0.rx.i1_4_lut_LC_15_18_0  (
            .in0(N__37851),
            .in1(N__37805),
            .in2(N__34252),
            .in3(N__37912),
            .lcout(\c0.rx.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_15_18_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_15_18_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__39194),
            .in2(_gnd_net_),
            .in3(N__34633),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71044),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_15_18_2 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \c0.rx.i2_4_lut_LC_15_18_2  (
            .in0(N__37852),
            .in1(N__37806),
            .in2(N__37753),
            .in3(N__37913),
            .lcout(n12492),
            .ltout(n12492_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i9378_3_lut_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.rx.i9378_3_lut_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i9378_3_lut_LC_15_18_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \c0.rx.i9378_3_lut_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__39433),
            .in2(N__34237),
            .in3(N__37853),
            .lcout(n12835),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_o_bdd_4_lut_4_lut_LC_15_18_4 .C_ON=1'b0;
    defparam \c0.tx_o_bdd_4_lut_4_lut_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_o_bdd_4_lut_4_lut_LC_15_18_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.tx_o_bdd_4_lut_4_lut_LC_15_18_4  (
            .in0(N__34234),
            .in1(N__34175),
            .in2(N__34120),
            .in3(N__34099),
            .lcout(\c0.n21611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__7__5375_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__7__5375_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__7__5375_LC_15_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__7__5375_LC_15_18_5  (
            .in0(N__33979),
            .in1(N__33945),
            .in2(_gnd_net_),
            .in3(N__46887),
            .lcout(data_out_frame_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71044),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_15_18_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_15_18_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_15_18_6  (
            .in0(N__39192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34309),
            .lcout(\c0.rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71044),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_15_18_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__39193),
            .in2(_gnd_net_),
            .in3(N__34297),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71044),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_15_19_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_15_19_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_15_19_0  (
            .in0(N__37652),
            .in1(N__37654),
            .in2(N__34683),
            .in3(N__34303),
            .lcout(n13179),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\c0.rx.n17267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_15_19_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_15_19_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_3_lut_LC_15_19_1  (
            .in0(N__37621),
            .in1(N__37617),
            .in2(N__34687),
            .in3(N__34300),
            .lcout(\c0.rx.n9 ),
            .ltout(),
            .carryin(\c0.rx.n17267 ),
            .carryout(\c0.rx.n17268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_15_19_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_15_19_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_4_lut_LC_15_19_2  (
            .in0(N__37687),
            .in1(N__37683),
            .in2(N__34684),
            .in3(N__34291),
            .lcout(n12908),
            .ltout(),
            .carryin(\c0.rx.n17268 ),
            .carryout(\c0.rx.n17269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_15_19_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_15_19_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_5_lut_LC_15_19_3  (
            .in0(N__39151),
            .in1(N__39150),
            .in2(N__34688),
            .in3(N__34288),
            .lcout(n12911),
            .ltout(),
            .carryin(\c0.rx.n17269 ),
            .carryout(\c0.rx.n17270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_15_19_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_15_19_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_6_lut_LC_15_19_4  (
            .in0(N__38107),
            .in1(N__38106),
            .in2(N__34685),
            .in3(N__34285),
            .lcout(n12914),
            .ltout(),
            .carryin(\c0.rx.n17270 ),
            .carryout(\c0.rx.n17271 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_15_19_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_15_19_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_7_lut_LC_15_19_5  (
            .in0(N__38083),
            .in1(N__38082),
            .in2(N__34689),
            .in3(N__34282),
            .lcout(n12917),
            .ltout(),
            .carryin(\c0.rx.n17271 ),
            .carryout(\c0.rx.n17272 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_15_19_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_15_19_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_8_lut_LC_15_19_6  (
            .in0(N__37723),
            .in1(N__37722),
            .in2(N__34686),
            .in3(N__34279),
            .lcout(n12920),
            .ltout(),
            .carryin(\c0.rx.n17272 ),
            .carryout(\c0.rx.n17273 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_15_19_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_15_19_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.rx.add_62_9_lut_LC_15_19_7  (
            .in0(N__39289),
            .in1(N__39290),
            .in2(N__34690),
            .in3(N__34636),
            .lcout(\c0.rx.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_431_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_431_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_431_LC_15_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_adj_431_LC_15_20_0  (
            .in0(N__49672),
            .in1(N__34557),
            .in2(N__34627),
            .in3(N__34590),
            .lcout(\c0.n45_adj_3262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_12_i6_2_lut_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.select_357_Select_12_i6_2_lut_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_12_i6_2_lut_LC_15_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_357_Select_12_i6_2_lut_LC_15_20_1  (
            .in0(N__60618),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34507),
            .lcout(\c0.n6_adj_3161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_25_i6_2_lut_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.select_357_Select_25_i6_2_lut_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_25_i6_2_lut_LC_15_20_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_25_i6_2_lut_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__34558),
            .in2(_gnd_net_),
            .in3(N__60620),
            .lcout(\c0.n6_adj_3172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_14_i6_2_lut_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.select_357_Select_14_i6_2_lut_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_14_i6_2_lut_LC_15_20_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.select_357_Select_14_i6_2_lut_LC_15_20_3  (
            .in0(N__60619),
            .in1(N__34464),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n6_adj_3194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_427_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_427_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_427_LC_15_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_427_LC_15_20_4  (
            .in0(N__34506),
            .in1(N__34481),
            .in2(N__34465),
            .in3(N__34440),
            .lcout(\c0.n43_adj_3257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_11_i6_2_lut_LC_15_20_6 .C_ON=1'b0;
    defparam \c0.select_357_Select_11_i6_2_lut_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_11_i6_2_lut_LC_15_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_11_i6_2_lut_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__60617),
            .in2(_gnd_net_),
            .in3(N__34336),
            .lcout(\c0.n6_adj_3160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_502_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_502_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_502_LC_15_20_7 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_502_LC_15_20_7  (
            .in0(N__40111),
            .in1(N__40286),
            .in2(N__49678),
            .in3(N__40201),
            .lcout(\c0.n12_adj_3361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_428_LC_15_21_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_428_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_428_LC_15_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_428_LC_15_21_0  (
            .in0(N__34386),
            .in1(N__35380),
            .in2(N__34363),
            .in3(N__34335),
            .lcout(),
            .ltout(\c0.n41_adj_3258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_430_LC_15_21_1 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_430_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_430_LC_15_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i24_4_lut_adj_430_LC_15_21_1  (
            .in0(N__35023),
            .in1(N__37966),
            .in2(N__34909),
            .in3(N__34906),
            .lcout(\c0.n50_adj_3261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_429_LC_15_21_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_429_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_429_LC_15_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_429_LC_15_21_2  (
            .in0(N__34900),
            .in1(N__34873),
            .in2(N__35302),
            .in3(N__34849),
            .lcout(\c0.n40_adj_3259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.i13_2_lut_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_LC_15_21_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i13_2_lut_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__35332),
            .in2(_gnd_net_),
            .in3(N__34816),
            .lcout(),
            .ltout(\c0.n39_adj_3260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_LC_15_21_4 .C_ON=1'b0;
    defparam \c0.i25_4_lut_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_LC_15_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i25_4_lut_LC_15_21_4  (
            .in0(N__34783),
            .in1(N__34777),
            .in2(N__34771),
            .in3(N__34768),
            .lcout(\c0.n11440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_930_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_930_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_930_LC_15_22_0 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \c0.i1_4_lut_adj_930_LC_15_22_0  (
            .in0(N__42364),
            .in1(N__35173),
            .in2(N__34969),
            .in3(N__34699),
            .lcout(),
            .ltout(\c0.n14_adj_3080_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_22_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i1_LC_15_22_1 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_15_22_1  (
            .in0(N__38354),
            .in1(N__34762),
            .in2(N__34744),
            .in3(N__34741),
            .lcout(FRAME_MATCHER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71093),
            .ce(),
            .sr(N__46803));
    defparam \c0.i1_3_lut_4_lut_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_15_22_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_15_22_3  (
            .in0(N__34728),
            .in1(N__34950),
            .in2(N__42496),
            .in3(N__42310),
            .lcout(\c0.n19119 ),
            .ltout(\c0.n19119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_463_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_463_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_463_LC_15_22_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \c0.i1_2_lut_adj_463_LC_15_22_4  (
            .in0(N__34965),
            .in1(_gnd_net_),
            .in2(N__34693),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n5_adj_3306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_22_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i0_LC_15_22_5 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_15_22_5  (
            .in0(N__39567),
            .in1(N__34981),
            .in2(N__34972),
            .in3(N__38317),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71093),
            .ce(),
            .sr(N__46803));
    defparam \c0.i1_2_lut_adj_460_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_460_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_460_LC_15_23_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i1_2_lut_adj_460_LC_15_23_0  (
            .in0(N__35123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35154),
            .lcout(\c0.n2_adj_3302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5__5168_LC_15_23_1 .C_ON=1'b0;
    defparam \c0.data_in_3__5__5168_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5__5168_LC_15_23_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__5__5168_LC_15_23_1  (
            .in0(N__67983),
            .in1(N__53176),
            .in2(_gnd_net_),
            .in3(N__39743),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71109),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_423_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_423_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_423_LC_15_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_423_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__38519),
            .in2(_gnd_net_),
            .in3(N__38413),
            .lcout(\c0.n9389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_581_LC_15_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_581_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_581_LC_15_23_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_581_LC_15_23_3  (
            .in0(N__39557),
            .in1(N__42427),
            .in2(N__38989),
            .in3(N__38258),
            .lcout(\c0.n11433 ),
            .ltout(\c0.n11433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_757_LC_15_23_4 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_757_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_757_LC_15_23_4 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_757_LC_15_23_4  (
            .in0(N__42428),
            .in1(N__38211),
            .in2(N__34957),
            .in3(N__42293),
            .lcout(),
            .ltout(\c0.n8_adj_3228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_396_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_396_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_396_LC_15_23_5 .LUT_INIT=16'b1111000000010000;
    LogicCell40 \c0.i4_4_lut_adj_396_LC_15_23_5  (
            .in0(N__38976),
            .in1(N__42429),
            .in2(N__34954),
            .in3(N__35423),
            .lcout(\c0.n2103 ),
            .ltout(\c0.n2103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_15_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_15_23_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_940_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__38520),
            .in2(N__34936),
            .in3(N__38414),
            .lcout(\c0.n1_adj_3002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3__5194_LC_15_23_7 .C_ON=1'b0;
    defparam \c0.data_in_0__3__5194_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3__5194_LC_15_23_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__3__5194_LC_15_23_7  (
            .in0(N__53195),
            .in1(N__39954),
            .in2(_gnd_net_),
            .in3(N__40012),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71109),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_509_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_509_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_509_LC_15_24_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_509_LC_15_24_0  (
            .in0(N__41365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34933),
            .lcout(\c0.n18653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_657_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_657_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_657_LC_15_24_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_657_LC_15_24_1  (
            .in0(N__38266),
            .in1(N__42459),
            .in2(_gnd_net_),
            .in3(N__39569),
            .lcout(n4_adj_3596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_15_24_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_15_24_2 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i1_3_lut_LC_15_24_2  (
            .in0(N__39891),
            .in1(N__38457),
            .in2(_gnd_net_),
            .in3(N__38469),
            .lcout(\c0.FRAME_MATCHER_state_31_N_1736_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_928_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_928_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_928_LC_15_24_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \c0.i1_4_lut_adj_928_LC_15_24_5  (
            .in0(N__38458),
            .in1(N__42460),
            .in2(N__39895),
            .in3(N__38416),
            .lcout(\c0.FRAME_MATCHER_state_31_N_1736_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_23_i6_2_lut_LC_15_24_6 .C_ON=1'b0;
    defparam \c0.select_357_Select_23_i6_2_lut_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_23_i6_2_lut_LC_15_24_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_23_i6_2_lut_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__60633),
            .in2(_gnd_net_),
            .in3(N__38019),
            .lcout(\c0.n6_adj_3176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_939_LC_15_24_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_939_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_939_LC_15_24_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_939_LC_15_24_7  (
            .in0(N__35150),
            .in1(N__38515),
            .in2(N__35133),
            .in3(N__38415),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_424_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_424_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_424_LC_15_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_424_LC_15_25_0  (
            .in0(N__35012),
            .in1(N__35083),
            .in2(N__35059),
            .in3(N__35251),
            .lcout(\c0.n44_adj_3255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5__5176_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.data_in_2__5__5176_LC_15_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5__5176_LC_15_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__5__5176_LC_15_26_0  (
            .in0(N__53215),
            .in1(N__39744),
            .in2(_gnd_net_),
            .in3(N__41877),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71153),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_24_i6_2_lut_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.select_357_Select_24_i6_2_lut_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_24_i6_2_lut_LC_15_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_24_i6_2_lut_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__60583),
            .in2(_gnd_net_),
            .in3(N__35014),
            .lcout(\c0.n6_adj_3174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_854_LC_15_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_854_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_854_LC_15_27_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_854_LC_15_27_1  (
            .in0(_gnd_net_),
            .in1(N__35473),
            .in2(_gnd_net_),
            .in3(N__41429),
            .lcout(\c0.n18675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_4_lut_LC_15_27_2.C_ON=1'b0;
    defparam i2_2_lut_3_lut_4_lut_LC_15_27_2.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_4_lut_LC_15_27_2.LUT_INIT=16'b1000110000000000;
    LogicCell40 i2_2_lut_3_lut_4_lut_LC_15_27_2 (
            .in0(N__42328),
            .in1(N__42368),
            .in2(N__42497),
            .in3(N__35436),
            .lcout(n2108),
            .ltout(n2108_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_26_i6_2_lut_LC_15_27_3 .C_ON=1'b0;
    defparam \c0.select_357_Select_26_i6_2_lut_LC_15_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_26_i6_2_lut_LC_15_27_3 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \c0.select_357_Select_26_i6_2_lut_LC_15_27_3  (
            .in0(_gnd_net_),
            .in1(N__35376),
            .in2(N__35356),
            .in3(_gnd_net_),
            .lcout(\c0.n6_adj_3170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_29_i6_2_lut_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.select_357_Select_29_i6_2_lut_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_29_i6_2_lut_LC_15_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_29_i6_2_lut_LC_15_28_1  (
            .in0(_gnd_net_),
            .in1(N__60585),
            .in2(_gnd_net_),
            .in3(N__37992),
            .lcout(\c0.n6_adj_3165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_27_i6_2_lut_LC_15_28_5 .C_ON=1'b0;
    defparam \c0.select_357_Select_27_i6_2_lut_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_27_i6_2_lut_LC_15_28_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_27_i6_2_lut_LC_15_28_5  (
            .in0(_gnd_net_),
            .in1(N__35328),
            .in2(_gnd_net_),
            .in3(N__60584),
            .lcout(\c0.n6_adj_3168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_28_i6_2_lut_LC_15_29_3 .C_ON=1'b0;
    defparam \c0.select_357_Select_28_i6_2_lut_LC_15_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_28_i6_2_lut_LC_15_29_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_28_i6_2_lut_LC_15_29_3  (
            .in0(_gnd_net_),
            .in1(N__35292),
            .in2(_gnd_net_),
            .in3(N__60632),
            .lcout(\c0.n6_adj_3166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_31_i6_2_lut_LC_15_31_2 .C_ON=1'b0;
    defparam \c0.select_357_Select_31_i6_2_lut_LC_15_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_31_i6_2_lut_LC_15_31_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_357_Select_31_i6_2_lut_LC_15_31_2  (
            .in0(N__60635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38134),
            .lcout(\c0.n6_adj_3159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_30_i6_2_lut_LC_15_31_3 .C_ON=1'b0;
    defparam \c0.select_357_Select_30_i6_2_lut_LC_15_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_30_i6_2_lut_LC_15_31_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_30_i6_2_lut_LC_15_31_3  (
            .in0(_gnd_net_),
            .in1(N__35247),
            .in2(_gnd_net_),
            .in3(N__60634),
            .lcout(\c0.n6_adj_3164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_61_i9_2_lut_3_lut_LC_16_7_0 .C_ON=1'b0;
    defparam \c0.equal_61_i9_2_lut_3_lut_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.equal_61_i9_2_lut_3_lut_LC_16_7_0 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.equal_61_i9_2_lut_3_lut_LC_16_7_0  (
            .in0(N__60204),
            .in1(N__59977),
            .in2(_gnd_net_),
            .in3(N__60108),
            .lcout(\c0.n9_adj_3038 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_6_i6_2_lut_LC_16_8_4 .C_ON=1'b0;
    defparam \c0.select_357_Select_6_i6_2_lut_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_6_i6_2_lut_LC_16_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_6_i6_2_lut_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__60717),
            .in2(_gnd_net_),
            .in3(N__40186),
            .lcout(\c0.n6_adj_3150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_82_i11_2_lut_LC_16_8_6 .C_ON=1'b0;
    defparam \c0.equal_82_i11_2_lut_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_82_i11_2_lut_LC_16_8_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.equal_82_i11_2_lut_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__49665),
            .in2(_gnd_net_),
            .in3(N__40185),
            .lcout(\c0.n11_adj_3093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i12_LC_16_9_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i12_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i12_LC_16_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter1.count_i0_i12_LC_16_9_1  (
            .in0(N__36255),
            .in1(N__37046),
            .in2(_gnd_net_),
            .in3(N__35791),
            .lcout(encoder1_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71156),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17732_4_lut_LC_16_9_6 .C_ON=1'b0;
    defparam \c0.i17732_4_lut_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17732_4_lut_LC_16_9_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.i17732_4_lut_LC_16_9_6  (
            .in0(N__37466),
            .in1(N__38542),
            .in2(N__35999),
            .in3(N__35737),
            .lcout(\c0.n21319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__2__5380_LC_16_10_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__2__5380_LC_16_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__2__5380_LC_16_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_7__2__5380_LC_16_10_1  (
            .in0(N__35767),
            .in1(N__35914),
            .in2(_gnd_net_),
            .in3(N__46859),
            .lcout(data_out_frame_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71140),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17730_4_lut_LC_16_10_5 .C_ON=1'b0;
    defparam \c0.i17730_4_lut_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17730_4_lut_LC_16_10_5 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \c0.i17730_4_lut_LC_16_10_5  (
            .in0(N__35902),
            .in1(N__36759),
            .in2(N__36988),
            .in3(N__35848),
            .lcout(\c0.n21317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i27_LC_16_10_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i27_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i27_LC_16_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \quad_counter0.count_i0_i27_LC_16_10_7  (
            .in0(N__35722),
            .in1(N__35529),
            .in2(_gnd_net_),
            .in3(N__35563),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71140),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_11_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_11_0  (
            .in0(N__35514),
            .in1(N__35503),
            .in2(_gnd_net_),
            .in3(N__40938),
            .lcout(\c0.n5_adj_3380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17735_4_lut_LC_16_11_4 .C_ON=1'b0;
    defparam \c0.i17735_4_lut_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17735_4_lut_LC_16_11_4 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.i17735_4_lut_LC_16_11_4  (
            .in0(N__37467),
            .in1(N__40654),
            .in2(N__36007),
            .in3(N__35479),
            .lcout(),
            .ltout(\c0.n21322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_4_lut_LC_16_11_5 .C_ON=1'b0;
    defparam \c0.i24_3_lut_4_lut_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_4_lut_LC_16_11_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.i24_3_lut_4_lut_LC_16_11_5  (
            .in0(N__37345),
            .in1(N__35941),
            .in2(N__35929),
            .in3(N__37468),
            .lcout(n10_adj_3594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_16_11_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_16_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_16_11_6  (
            .in0(N__35913),
            .in1(N__35871),
            .in2(_gnd_net_),
            .in3(N__40937),
            .lcout(\c0.n5_adj_3106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_62_i9_2_lut_3_lut_LC_16_11_7 .C_ON=1'b0;
    defparam \c0.equal_62_i9_2_lut_3_lut_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.equal_62_i9_2_lut_3_lut_LC_16_11_7 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.equal_62_i9_2_lut_3_lut_LC_16_11_7  (
            .in0(N__60256),
            .in1(N__59978),
            .in2(_gnd_net_),
            .in3(N__60116),
            .lcout(\c0.n9_adj_3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__2__5436_LC_16_12_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__2__5436_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__2__5436_LC_16_12_0 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \c0.data_out_frame_0__2__5436_LC_16_12_0  (
            .in0(N__39490),
            .in1(N__35860),
            .in2(N__37092),
            .in3(N__39003),
            .lcout(\c0.data_out_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71110),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__2__5388_LC_16_12_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__2__5388_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__2__5388_LC_16_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_6__2__5388_LC_16_12_1  (
            .in0(N__46856),
            .in1(N__35896),
            .in2(_gnd_net_),
            .in3(N__35872),
            .lcout(data_out_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71110),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17928_2_lut_LC_16_12_2 .C_ON=1'b0;
    defparam \c0.i17928_2_lut_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17928_2_lut_LC_16_12_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i17928_2_lut_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__36716),
            .in2(_gnd_net_),
            .in3(N__35859),
            .lcout(),
            .ltout(\c0.n21473_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_16_12_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_16_12_3 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_16_12_3  (
            .in0(N__36969),
            .in1(N__40906),
            .in2(N__35851),
            .in3(N__36403),
            .lcout(\c0.n6_adj_3105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__6__5208_LC_16_12_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__6__5208_LC_16_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__6__5208_LC_16_12_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \c0.data_out_frame_28__6__5208_LC_16_12_5  (
            .in0(N__46855),
            .in1(N__50605),
            .in2(N__54481),
            .in3(N__35829),
            .lcout(data_out_frame_28_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71110),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__3__5435_LC_16_12_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__3__5435_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__3__5435_LC_16_12_6 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \c0.data_out_frame_0__3__5435_LC_16_12_6  (
            .in0(N__39491),
            .in1(N__35815),
            .in2(N__37093),
            .in3(N__39004),
            .lcout(\c0.data_out_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71110),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_3_lut_4_lut_LC_16_12_7 .C_ON=1'b0;
    defparam \c0.i16_3_lut_4_lut_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i16_3_lut_4_lut_LC_16_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_3_lut_4_lut_LC_16_12_7  (
            .in0(N__55511),
            .in1(N__51345),
            .in2(N__57379),
            .in3(N__51291),
            .lcout(\c0.n39_adj_3339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i101_LC_16_13_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i101_LC_16_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i101_LC_16_13_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i101_LC_16_13_0  (
            .in0(N__66194),
            .in1(N__67197),
            .in2(N__44624),
            .in3(N__72697),
            .lcout(\c0.data_in_frame_12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71094),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_16_13_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_16_13_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_16_13_1  (
            .in0(N__37183),
            .in1(N__36330),
            .in2(N__40936),
            .in3(_gnd_net_),
            .lcout(\c0.n11_adj_3325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__0__5342_LC_16_13_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__0__5342_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__0__5342_LC_16_13_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame_12__0__5342_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__46848),
            .in2(N__36334),
            .in3(N__36370),
            .lcout(data_out_frame_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71094),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__7__5343_LC_16_13_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__7__5343_LC_16_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__7__5343_LC_16_13_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame_11__7__5343_LC_16_13_3  (
            .in0(N__36318),
            .in1(N__36291),
            .in2(N__46916),
            .in3(_gnd_net_),
            .lcout(data_out_frame_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71094),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i28_LC_16_13_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i28_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i28_LC_16_13_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i28_LC_16_13_4  (
            .in0(N__36277),
            .in1(N__36262),
            .in2(_gnd_net_),
            .in3(N__36074),
            .lcout(encoder1_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71094),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__6__5392_LC_16_13_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__6__5392_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__6__5392_LC_16_13_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.data_out_frame_5__6__5392_LC_16_13_5  (
            .in0(N__36049),
            .in1(N__38632),
            .in2(N__46917),
            .in3(_gnd_net_),
            .lcout(data_out_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71094),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_16_13_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_16_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_16_13_6  (
            .in0(N__36037),
            .in1(N__36018),
            .in2(_gnd_net_),
            .in3(N__40923),
            .lcout(),
            .ltout(\c0.n26_adj_3382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17729_4_lut_LC_16_13_7 .C_ON=1'b0;
    defparam \c0.i17729_4_lut_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17729_4_lut_LC_16_13_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.i17729_4_lut_LC_16_13_7  (
            .in0(N__37464),
            .in1(N__36000),
            .in2(N__35965),
            .in3(N__35962),
            .lcout(\c0.n21316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__4__5394_LC_16_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__4__5394_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__4__5394_LC_16_14_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame_5__4__5394_LC_16_14_0  (
            .in0(N__46865),
            .in1(_gnd_net_),
            .in2(N__36487),
            .in3(N__38752),
            .lcout(data_out_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71081),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17913_2_lut_LC_16_14_1 .C_ON=1'b0;
    defparam \c0.i17913_2_lut_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17913_2_lut_LC_16_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i17913_2_lut_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__36483),
            .in2(_gnd_net_),
            .in3(N__40892),
            .lcout(\c0.n21465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__0__5398_LC_16_14_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__0__5398_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__0__5398_LC_16_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame_5__0__5398_LC_16_14_3  (
            .in0(N__36460),
            .in1(N__39088),
            .in2(_gnd_net_),
            .in3(N__46866),
            .lcout(\c0.data_out_frame_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71081),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i5_LC_16_14_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i5_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i5_LC_16_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i5_LC_16_14_4  (
            .in0(N__36441),
            .in1(N__55384),
            .in2(_gnd_net_),
            .in3(N__41096),
            .lcout(control_mode_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71081),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17980_4_lut_LC_16_14_5 .C_ON=1'b0;
    defparam \c0.i17980_4_lut_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17980_4_lut_LC_16_14_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.i17980_4_lut_LC_16_14_5  (
            .in0(N__36430),
            .in1(N__36949),
            .in2(N__36418),
            .in3(N__36735),
            .lcout(\c0.n21568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__2__5396_LC_16_14_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__2__5396_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__2__5396_LC_16_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame_5__2__5396_LC_16_14_6  (
            .in0(N__46864),
            .in1(N__38620),
            .in2(_gnd_net_),
            .in3(N__36402),
            .lcout(data_out_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71081),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i205_LC_16_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i205_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i205_LC_16_14_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i205_LC_16_14_7  (
            .in0(N__66899),
            .in1(N__63395),
            .in2(N__59669),
            .in3(N__72711),
            .lcout(\c0.data_in_frame_25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71081),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i146_LC_16_15_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i146_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i146_LC_16_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i146_LC_16_15_0  (
            .in0(N__71485),
            .in1(N__63937),
            .in2(_gnd_net_),
            .in3(N__45234),
            .lcout(data_in_frame_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71069),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_16_15_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_16_15_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__39204),
            .in2(_gnd_net_),
            .in3(N__36388),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71069),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_16_15_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_16_15_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_16_15_2  (
            .in0(N__39205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37165),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71069),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__7__5391_LC_16_15_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__7__5391_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__7__5391_LC_16_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_5__7__5391_LC_16_15_3  (
            .in0(N__38722),
            .in1(N__37006),
            .in2(_gnd_net_),
            .in3(N__46764),
            .lcout(data_out_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71069),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_16_15_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_16_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_16_15_6  (
            .in0(N__50863),
            .in1(N__54976),
            .in2(N__50944),
            .in3(N__50829),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_243_LC_16_15_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_243_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_243_LC_16_15_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.i4_4_lut_adj_243_LC_16_15_7  (
            .in0(N__37153),
            .in1(N__37135),
            .in2(N__37111),
            .in3(N__38812),
            .lcout(\c0.n12254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__4__5338_LC_16_16_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__4__5338_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__4__5338_LC_16_16_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame_12__4__5338_LC_16_16_1  (
            .in0(N__37059),
            .in1(N__37023),
            .in2(N__46857),
            .in3(_gnd_net_),
            .lcout(data_out_frame_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71056),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17988_3_lut_LC_16_16_2 .C_ON=1'b0;
    defparam \c0.i17988_3_lut_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17988_3_lut_LC_16_16_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \c0.i17988_3_lut_LC_16_16_2  (
            .in0(N__36960),
            .in1(N__37005),
            .in2(_gnd_net_),
            .in3(N__40886),
            .lcout(),
            .ltout(\c0.n21576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17715_4_lut_LC_16_16_3 .C_ON=1'b0;
    defparam \c0.i17715_4_lut_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17715_4_lut_LC_16_16_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i17715_4_lut_LC_16_16_3  (
            .in0(N__36994),
            .in1(N__36961),
            .in2(N__36769),
            .in3(N__36697),
            .lcout(),
            .ltout(\c0.n21302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17717_4_lut_LC_16_16_4 .C_ON=1'b0;
    defparam \c0.i17717_4_lut_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17717_4_lut_LC_16_16_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.i17717_4_lut_LC_16_16_4  (
            .in0(N__46951),
            .in1(N__37524),
            .in2(N__36508),
            .in3(N__37462),
            .lcout(),
            .ltout(\c0.n21304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_4_lut_LC_16_16_5 .C_ON=1'b0;
    defparam \c0.i23_3_lut_4_lut_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_4_lut_LC_16_16_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.i23_3_lut_4_lut_LC_16_16_5  (
            .in0(N__37463),
            .in1(N__37344),
            .in2(N__36505),
            .in3(N__36502),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17723_4_lut_LC_16_16_6 .C_ON=1'b0;
    defparam \c0.i17723_4_lut_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17723_4_lut_LC_16_16_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.i17723_4_lut_LC_16_16_6  (
            .in0(N__37525),
            .in1(N__37460),
            .in2(N__37498),
            .in3(N__37474),
            .lcout(),
            .ltout(\c0.n21310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_4_lut_adj_620_LC_16_16_7 .C_ON=1'b0;
    defparam \c0.i23_3_lut_4_lut_adj_620_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_4_lut_adj_620_LC_16_16_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.i23_3_lut_4_lut_adj_620_LC_16_16_7  (
            .in0(N__37461),
            .in1(N__37343),
            .in2(N__37255),
            .in3(N__37252),
            .lcout(n9_adj_3590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_16_17_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.rx.i3_4_lut_LC_16_17_0  (
            .in0(N__37849),
            .in1(N__37796),
            .in2(N__37930),
            .in3(N__37744),
            .lcout(\c0.rx.n11302 ),
            .ltout(\c0.rx.n11302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_16_17_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_16_17_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.rx.i1_2_lut_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37219),
            .in3(N__39335),
            .lcout(n11466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__0__5334_LC_16_17_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__0__5334_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__0__5334_LC_16_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame_13__0__5334_LC_16_17_2  (
            .in0(N__37216),
            .in1(N__37182),
            .in2(_gnd_net_),
            .in3(N__46643),
            .lcout(data_out_frame_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71035),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i17914_2_lut_3_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \c0.rx.i17914_2_lut_3_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i17914_2_lut_3_lut_LC_16_17_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.i17914_2_lut_3_lut_LC_16_17_3  (
            .in0(N__56213),
            .in1(N__37927),
            .in2(_gnd_net_),
            .in3(N__39221),
            .lcout(),
            .ltout(\c0.rx.n21451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_16_17_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_16_17_4 .LUT_INIT=16'b0000000001110010;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_16_17_4  (
            .in0(N__37850),
            .in1(N__37570),
            .in2(N__37168),
            .in3(N__37797),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71035),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_516_LC_16_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_516_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_516_LC_16_17_5 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_516_LC_16_17_5  (
            .in0(N__40280),
            .in1(N__49677),
            .in2(N__40126),
            .in3(N__40200),
            .lcout(\c0.n12_adj_3006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i147_LC_16_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i147_LC_16_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i147_LC_16_17_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i147_LC_16_17_6  (
            .in0(N__43116),
            .in1(N__63915),
            .in2(_gnd_net_),
            .in3(N__68622),
            .lcout(data_in_frame_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71035),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_656_LC_16_17_7 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_656_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_656_LC_16_17_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_656_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__63576),
            .in2(_gnd_net_),
            .in3(N__63651),
            .lcout(\c0.n27_adj_3455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_adj_213_LC_16_18_0 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_adj_213_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_adj_213_LC_16_18_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \c0.rx.i2_4_lut_adj_213_LC_16_18_0  (
            .in0(N__39136),
            .in1(N__37715),
            .in2(N__37564),
            .in3(N__39244),
            .lcout(\c0.rx.n15906 ),
            .ltout(\c0.rx.n15906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_208_LC_16_18_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_208_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_208_LC_16_18_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.rx.i2_3_lut_adj_208_LC_16_18_1  (
            .in0(N__39284),
            .in1(_gnd_net_),
            .in2(N__37573),
            .in3(N__37922),
            .lcout(\c0.rx.n20851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_211_LC_16_18_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_211_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_211_LC_16_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_211_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__37682),
            .in2(_gnd_net_),
            .in3(N__37610),
            .lcout(\c0.rx.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_16_18_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_16_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__39285),
            .in2(_gnd_net_),
            .in3(N__37549),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71057),
            .ce(),
            .sr(N__37555));
    defparam \c0.rx.i2_3_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_16_18_5 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.rx.i2_3_lut_LC_16_18_5  (
            .in0(N__37862),
            .in1(N__37921),
            .in2(_gnd_net_),
            .in3(N__37801),
            .lcout(\c0.rx.n20964 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i12463_2_lut_LC_16_18_6 .C_ON=1'b0;
    defparam \c0.rx.i12463_2_lut_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i12463_2_lut_LC_16_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i12463_2_lut_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__39283),
            .in2(_gnd_net_),
            .in3(N__37548),
            .lcout(r_SM_Main_2_N_2473_2),
            .ltout(r_SM_Main_2_N_2473_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_16_18_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_16_18_7 .LUT_INIT=16'b1111000000111111;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__39432),
            .in2(N__37540),
            .in3(N__37923),
            .lcout(\c0.rx.n15926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_215_LC_16_19_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_215_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_215_LC_16_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_215_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__38104),
            .in2(_gnd_net_),
            .in3(N__38080),
            .lcout(\c0.rx.n11455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_214_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_214_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_214_LC_16_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_214_LC_16_19_1  (
            .in0(N__37680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37648),
            .lcout(),
            .ltout(\c0.rx.n35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5_4_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.rx.i5_4_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5_4_lut_LC_16_19_2 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \c0.rx.i5_4_lut_LC_16_19_2  (
            .in0(N__37714),
            .in1(N__38059),
            .in2(N__37933),
            .in3(N__56154),
            .lcout(),
            .ltout(\c0.rx.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i17900_4_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.rx.i17900_4_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i17900_4_lut_LC_16_19_3 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \c0.rx.i17900_4_lut_LC_16_19_3  (
            .in0(N__37585),
            .in1(N__37928),
            .in2(N__37873),
            .in3(N__39142),
            .lcout(),
            .ltout(\c0.rx.n21406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_216_LC_16_19_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_216_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_216_LC_16_19_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \c0.rx.i1_4_lut_adj_216_LC_16_19_4  (
            .in0(N__37863),
            .in1(N__37798),
            .in2(N__37756),
            .in3(N__37748),
            .lcout(n3792),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_4_lut_LC_16_19_5 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_4_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_4_lut_LC_16_19_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.rx.i1_3_lut_4_lut_LC_16_19_5  (
            .in0(N__37679),
            .in1(N__37713),
            .in2(N__37653),
            .in3(N__37608),
            .lcout(\c0.rx.n6_adj_2995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_LC_16_19_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_LC_16_19_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_LC_16_19_7  (
            .in0(N__37681),
            .in1(N__37647),
            .in2(_gnd_net_),
            .in3(N__37609),
            .lcout(\c0.rx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_16_20_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__39190),
            .in2(_gnd_net_),
            .in3(N__37579),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71082),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_925_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_925_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_925_LC_16_20_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_925_LC_16_20_1  (
            .in0(N__44260),
            .in1(N__71623),
            .in2(_gnd_net_),
            .in3(N__59432),
            .lcout(n19129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_16_20_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__39191),
            .in2(_gnd_net_),
            .in3(N__38200),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71082),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_432_LC_16_20_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_432_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_432_LC_16_20_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_432_LC_16_20_3  (
            .in0(N__40110),
            .in1(N__40285),
            .in2(_gnd_net_),
            .in3(N__38186),
            .lcout(),
            .ltout(\c0.n11317_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12193_3_lut_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.i12193_3_lut_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12193_3_lut_LC_16_20_4 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \c0.i12193_3_lut_LC_16_20_4  (
            .in0(N__64340),
            .in1(_gnd_net_),
            .in2(N__38170),
            .in3(N__38160),
            .lcout(\c0.n3632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i119_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i119_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i119_LC_16_20_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i119_LC_16_20_5  (
            .in0(N__69001),
            .in1(N__64136),
            .in2(N__64887),
            .in3(N__62018),
            .lcout(\c0.data_in_frame_14_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71082),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i17680_2_lut_3_lut_LC_16_20_6 .C_ON=1'b0;
    defparam \c0.rx.i17680_2_lut_3_lut_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i17680_2_lut_3_lut_LC_16_20_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.rx.i17680_2_lut_3_lut_LC_16_20_6  (
            .in0(N__39292),
            .in1(N__38105),
            .in2(_gnd_net_),
            .in3(N__38081),
            .lcout(\c0.rx.n21267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_426_LC_16_21_0 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_426_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_426_LC_16_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_426_LC_16_21_0  (
            .in0(N__38050),
            .in1(N__40199),
            .in2(N__38026),
            .in3(N__37999),
            .lcout(\c0.n42_adj_3256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_920_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_920_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_920_LC_16_21_3 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_920_LC_16_21_3  (
            .in0(N__61955),
            .in1(N__71624),
            .in2(_gnd_net_),
            .in3(N__59448),
            .lcout(n19127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_228_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_228_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_228_LC_16_21_4 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \c0.i1_4_lut_adj_228_LC_16_21_4  (
            .in0(N__37959),
            .in1(N__38277),
            .in2(N__42495),
            .in3(N__37942),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12257_2_lut_4_lut_LC_16_21_6 .C_ON=1'b0;
    defparam \c0.i12257_2_lut_4_lut_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i12257_2_lut_4_lut_LC_16_21_6 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \c0.i12257_2_lut_4_lut_LC_16_21_6  (
            .in0(N__53079),
            .in1(N__38373),
            .in2(N__38806),
            .in3(N__42369),
            .lcout(\c0.n15701 ),
            .ltout(\c0.n15701_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_864_LC_16_21_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_864_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_864_LC_16_21_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_864_LC_16_21_7  (
            .in0(N__40287),
            .in1(N__38398),
            .in2(N__38386),
            .in3(N__40125),
            .lcout(\c0.n19098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_16_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_16_22_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_658_LC_16_22_0  (
            .in0(N__38931),
            .in1(N__39552),
            .in2(_gnd_net_),
            .in3(N__38248),
            .lcout(n11421),
            .ltout(n11421_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_483_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_483_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_483_LC_16_22_1 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \c0.i1_2_lut_adj_483_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38383),
            .in3(N__42426),
            .lcout(\c0.n11422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6__5167_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.data_in_3__6__5167_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6__5167_LC_16_22_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__6__5167_LC_16_22_3  (
            .in0(N__69012),
            .in1(N__53174),
            .in2(_gnd_net_),
            .in3(N__52949),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71111),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_662_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_662_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_662_LC_16_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_662_LC_16_22_6  (
            .in0(N__38348),
            .in1(N__38212),
            .in2(N__38964),
            .in3(N__38313),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i117_LC_16_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i117_LC_16_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i117_LC_16_22_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i117_LC_16_22_7  (
            .in0(N__72775),
            .in1(N__64113),
            .in2(N__61987),
            .in3(N__45127),
            .lcout(\c0.data_in_frame_14_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71111),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_885_LC_16_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_885_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_885_LC_16_23_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_885_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__66121),
            .in2(_gnd_net_),
            .in3(N__59439),
            .lcout(\c0.n19140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6__5183_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.data_in_1__6__5183_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6__5183_LC_16_23_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__6__5183_LC_16_23_1  (
            .in0(N__52919),
            .in1(N__53177),
            .in2(_gnd_net_),
            .in3(N__39802),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71124),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_482_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_482_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_482_LC_16_23_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.i1_2_lut_adj_482_LC_16_23_3  (
            .in0(N__39556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38265),
            .lcout(\c0.n15874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_421_LC_16_23_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_421_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_421_LC_16_23_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.i9_4_lut_adj_421_LC_16_23_5  (
            .in0(N__43907),
            .in1(N__49754),
            .in2(N__47014),
            .in3(N__39846),
            .lcout(\c0.n21_adj_3253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1__5180_LC_16_23_6 .C_ON=1'b0;
    defparam \c0.data_in_2__1__5180_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1__5180_LC_16_23_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_2__1__5180_LC_16_23_6  (
            .in0(N__39847),
            .in1(N__53178),
            .in2(_gnd_net_),
            .in3(N__43908),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71124),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i201_LC_16_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i201_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i201_LC_16_23_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i201_LC_16_23_7  (
            .in0(N__63412),
            .in1(N__66849),
            .in2(N__53379),
            .in3(N__65172),
            .lcout(\c0.data_in_frame_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71124),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12187_3_lut_LC_16_24_0 .C_ON=1'b0;
    defparam \c0.i12187_3_lut_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12187_3_lut_LC_16_24_0 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \c0.i12187_3_lut_LC_16_24_0  (
            .in0(N__38425),
            .in1(N__38978),
            .in2(_gnd_net_),
            .in3(N__38449),
            .lcout(\c0.n121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3__5170_LC_16_24_1 .C_ON=1'b0;
    defparam \c0.data_in_3__3__5170_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3__5170_LC_16_24_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__3__5170_LC_16_24_1  (
            .in0(N__69376),
            .in1(N__53175),
            .in2(_gnd_net_),
            .in3(N__39867),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71141),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_417_LC_16_24_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_417_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_417_LC_16_24_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i6_4_lut_adj_417_LC_16_24_2  (
            .in0(N__47034),
            .in1(N__39980),
            .in2(N__47013),
            .in3(N__39751),
            .lcout(\c0.n63_adj_3083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_312_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_312_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_312_LC_16_24_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.i2_3_lut_adj_312_LC_16_24_3  (
            .in0(N__49755),
            .in1(N__38533),
            .in2(_gnd_net_),
            .in3(N__40579),
            .lcout(\c0.n103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_16_24_5 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_16_24_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i11_3_lut_LC_16_24_5  (
            .in0(N__38436),
            .in1(N__38443),
            .in2(_gnd_net_),
            .in3(N__39711),
            .lcout(\c0.n63_adj_3084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_420_LC_16_24_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_420_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_420_LC_16_24_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i7_4_lut_adj_420_LC_16_24_6  (
            .in0(N__39866),
            .in1(N__39666),
            .in2(N__39829),
            .in3(N__41902),
            .lcout(\c0.n19_adj_3252 ),
            .ltout(\c0.n19_adj_3252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4379_2_lut_4_lut_LC_16_24_7 .C_ON=1'b0;
    defparam \c0.i4379_2_lut_4_lut_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4379_2_lut_4_lut_LC_16_24_7 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i4379_2_lut_4_lut_LC_16_24_7  (
            .in0(N__38437),
            .in1(N__39712),
            .in2(N__38428),
            .in3(N__38424),
            .lcout(\c0.n7804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__6__5191_LC_16_25_1 .C_ON=1'b0;
    defparam \c0.data_in_0__6__5191_LC_16_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6__5191_LC_16_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__6__5191_LC_16_25_1  (
            .in0(N__53172),
            .in1(N__39981),
            .in2(_gnd_net_),
            .in3(N__39806),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71155),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2__5195_LC_16_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0__2__5195_LC_16_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2__5195_LC_16_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__2__5195_LC_16_25_2  (
            .in0(N__38494),
            .in1(N__53173),
            .in2(_gnd_net_),
            .in3(N__39667),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71155),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17694_4_lut_LC_16_25_3 .C_ON=1'b0;
    defparam \c0.i17694_4_lut_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17694_4_lut_LC_16_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i17694_4_lut_LC_16_25_3  (
            .in0(N__41876),
            .in1(N__40004),
            .in2(N__42636),
            .in3(N__38493),
            .lcout(),
            .ltout(\c0.n21281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_399_LC_16_25_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_399_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_399_LC_16_25_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i10_4_lut_adj_399_LC_16_25_4  (
            .in0(N__39775),
            .in1(N__42589),
            .in2(N__38536),
            .in3(N__42544),
            .lcout(\c0.n108 ),
            .ltout(\c0.n108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_422_LC_16_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_422_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_422_LC_16_25_5 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i3_4_lut_adj_422_LC_16_25_5  (
            .in0(N__40575),
            .in1(N__39879),
            .in2(N__38527),
            .in3(N__49734),
            .lcout(\c0.n92_adj_3254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i231_LC_16_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i231_LC_16_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i231_LC_16_25_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i231_LC_16_25_7  (
            .in0(N__66933),
            .in1(N__69024),
            .in2(N__39702),
            .in3(N__67199),
            .lcout(\c0.data_in_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71155),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0__5181_LC_16_26_1 .C_ON=1'b0;
    defparam \c0.data_in_2__0__5181_LC_16_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0__5181_LC_16_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__0__5181_LC_16_26_1  (
            .in0(N__53216),
            .in1(N__49756),
            .in2(_gnd_net_),
            .in3(N__42632),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71166),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_411_LC_16_26_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_411_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_411_LC_16_26_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i7_4_lut_adj_411_LC_16_26_3  (
            .in0(N__40003),
            .in1(N__41875),
            .in2(N__39808),
            .in3(N__38491),
            .lcout(\c0.n18_adj_3246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2__5187_LC_16_26_4 .C_ON=1'b0;
    defparam \c0.data_in_1__2__5187_LC_16_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2__5187_LC_16_26_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_1__2__5187_LC_16_26_4  (
            .in0(N__38492),
            .in1(N__53217),
            .in2(_gnd_net_),
            .in3(N__41929),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71166),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_259_LC_16_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_259_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_259_LC_16_27_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_259_LC_16_27_1  (
            .in0(_gnd_net_),
            .in1(N__40316),
            .in2(_gnd_net_),
            .in3(N__41428),
            .lcout(\c0.n18655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_7_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_17_7_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_17_7_7  (
            .in0(N__43762),
            .in1(N__65148),
            .in2(N__56236),
            .in3(N__56084),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71190),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_17_8_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_17_8_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__40590),
            .in2(N__40615),
            .in3(N__40942),
            .lcout(\c0.n26_adj_3107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_725_LC_17_8_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_725_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_725_LC_17_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_725_LC_17_8_1  (
            .in0(N__54706),
            .in1(N__38551),
            .in2(N__55402),
            .in3(N__40597),
            .lcout(\c0.n15499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_17_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_17_8_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i53_LC_17_8_2  (
            .in0(N__72614),
            .in1(N__61677),
            .in2(N__46369),
            .in3(N__61927),
            .lcout(\c0.data_in_frame_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71179),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_adj_358_LC_17_8_3 .C_ON=1'b0;
    defparam \c0.i9_2_lut_adj_358_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_adj_358_LC_17_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i9_2_lut_adj_358_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__54254),
            .in2(_gnd_net_),
            .in3(N__61117),
            .lcout(\c0.n37_adj_3153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_477_LC_17_8_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_477_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_477_LC_17_8_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.i17_4_lut_adj_477_LC_17_8_4  (
            .in0(N__54589),
            .in1(N__54892),
            .in2(N__40639),
            .in3(N__55184),
            .lcout(\c0.n38_adj_3328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i155_LC_17_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i155_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i155_LC_17_9_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_frame_0__i155_LC_17_9_0  (
            .in0(N__69168),
            .in1(_gnd_net_),
            .in2(N__65762),
            .in3(N__68655),
            .lcout(data_in_frame_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71168),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i118_LC_17_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i118_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i118_LC_17_9_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i118_LC_17_9_1  (
            .in0(N__61954),
            .in1(N__64248),
            .in2(N__44712),
            .in3(N__67922),
            .lcout(\c0.data_in_frame_14_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71168),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17692_4_lut_LC_17_9_2 .C_ON=1'b0;
    defparam \c0.i17692_4_lut_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17692_4_lut_LC_17_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17692_4_lut_LC_17_9_2  (
            .in0(N__46302),
            .in1(N__47221),
            .in2(N__42703),
            .in3(N__54468),
            .lcout(),
            .ltout(\c0.n21279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_480_LC_17_9_3 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_480_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_480_LC_17_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.i20_4_lut_adj_480_LC_17_9_3  (
            .in0(N__47311),
            .in1(N__38575),
            .in2(N__38569),
            .in3(N__38563),
            .lcout(FRAME_MATCHER_state_31_N_1800_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17668_2_lut_LC_17_9_4 .C_ON=1'b0;
    defparam \c0.i17668_2_lut_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17668_2_lut_LC_17_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i17668_2_lut_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__47560),
            .in2(_gnd_net_),
            .in3(N__56852),
            .lcout(),
            .ltout(\c0.n21255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_488_LC_17_9_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_488_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_488_LC_17_9_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.i16_4_lut_adj_488_LC_17_9_5  (
            .in0(N__62172),
            .in1(N__50360),
            .in2(N__38566),
            .in3(N__55054),
            .lcout(\c0.n37_adj_3332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_adj_555_LC_17_10_0 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_adj_555_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_adj_555_LC_17_10_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i11_2_lut_3_lut_adj_555_LC_17_10_0  (
            .in0(N__61246),
            .in1(_gnd_net_),
            .in2(N__38607),
            .in3(N__44310),
            .lcout(\c0.n63_adj_3417 ),
            .ltout(\c0.n63_adj_3417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_2_lut_3_lut_4_lut_LC_17_10_1 .C_ON=1'b0;
    defparam \c0.i16_2_lut_3_lut_4_lut_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_2_lut_3_lut_4_lut_LC_17_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_2_lut_3_lut_4_lut_LC_17_10_1  (
            .in0(N__41027),
            .in1(N__44049),
            .in2(N__38557),
            .in3(N__51259),
            .lcout(\c0.n40_adj_3032 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_17_10_2 .C_ON=1'b0;
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_17_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_2_lut_3_lut_4_lut_LC_17_10_2  (
            .in0(N__51260),
            .in1(N__41028),
            .in2(N__44053),
            .in3(N__50500),
            .lcout(\c0.n34_adj_3411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_554_LC_17_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_554_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_554_LC_17_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_554_LC_17_10_3  (
            .in0(N__44311),
            .in1(N__38600),
            .in2(_gnd_net_),
            .in3(N__41029),
            .lcout(\c0.n5_adj_3040 ),
            .ltout(\c0.n5_adj_3040_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_533_LC_17_10_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_533_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_533_LC_17_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_533_LC_17_10_4  (
            .in0(N__51258),
            .in1(_gnd_net_),
            .in2(N__38554),
            .in3(N__44048),
            .lcout(\c0.n11537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_433_LC_17_10_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_433_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_433_LC_17_10_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i13_4_lut_adj_433_LC_17_10_5  (
            .in0(N__41014),
            .in1(N__57289),
            .in2(N__42756),
            .in3(N__50830),
            .lcout(\c0.n30_adj_3264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_17_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_17_10_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i41_LC_17_10_6  (
            .in0(N__65069),
            .in1(N__61795),
            .in2(N__38608),
            .in3(N__60309),
            .lcout(\c0.data_in_frame_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71157),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_17_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_17_10_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i43_LC_17_10_7  (
            .in0(N__61794),
            .in1(N__68656),
            .in2(N__60329),
            .in3(N__61247),
            .lcout(\c0.data_in_frame_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71157),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_17_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_17_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_17_11_1  (
            .in0(N__56846),
            .in1(N__61122),
            .in2(N__54472),
            .in3(N__46303),
            .lcout(\c0.n6_adj_3343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_242_LC_17_11_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_242_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_242_LC_17_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_242_LC_17_11_2  (
            .in0(N__55549),
            .in1(N__49813),
            .in2(N__38589),
            .in3(N__61351),
            .lcout(\c0.n19493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i103_LC_17_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i103_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i103_LC_17_11_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i103_LC_17_11_3  (
            .in0(N__66038),
            .in1(N__67196),
            .in2(N__66286),
            .in3(N__68928),
            .lcout(\c0.data_in_frame_12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71142),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i80_LC_17_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i80_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i80_LC_17_11_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i80_LC_17_11_4  (
            .in0(N__72284),
            .in1(N__63281),
            .in2(N__38590),
            .in3(N__66039),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71142),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_17_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_17_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_17_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i42_LC_17_11_6  (
            .in0(N__60319),
            .in1(N__61797),
            .in2(N__51406),
            .in3(N__71436),
            .lcout(\c0.data_in_frame_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71142),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_17_11_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_17_11_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i19_LC_17_11_7  (
            .in0(N__61796),
            .in1(N__44247),
            .in2(N__68724),
            .in3(N__46333),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71142),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i125_LC_17_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i125_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i125_LC_17_12_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i125_LC_17_12_0  (
            .in0(N__64410),
            .in1(N__64220),
            .in2(N__51582),
            .in3(N__72672),
            .lcout(\c0.data_in_frame_15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71125),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_868_LC_17_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_868_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_868_LC_17_12_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_868_LC_17_12_1  (
            .in0(N__59992),
            .in1(N__60121),
            .in2(N__60264),
            .in3(N__59481),
            .lcout(\c0.n19115 ),
            .ltout(\c0.n19115_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i77_LC_17_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i77_LC_17_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i77_LC_17_12_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i77_LC_17_12_2  (
            .in0(N__41141),
            .in1(N__66046),
            .in2(N__38692),
            .in3(N__72673),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71125),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_17_12_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_17_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_17_12_3  (
            .in0(N__43149),
            .in1(N__38763),
            .in2(N__38689),
            .in3(N__50659),
            .lcout(\c0.n16_adj_3018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_653_LC_17_12_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_653_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_653_LC_17_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_653_LC_17_12_4  (
            .in0(N__49921),
            .in1(N__54893),
            .in2(N__42940),
            .in3(N__42969),
            .lcout(\c0.n12_adj_3477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i82_LC_17_12_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i82_LC_17_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i82_LC_17_12_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i82_LC_17_12_5  (
            .in0(N__66045),
            .in1(N__38688),
            .in2(N__71525),
            .in3(N__62846),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71125),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i74_LC_17_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i74_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i74_LC_17_12_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i74_LC_17_12_7  (
            .in0(N__71492),
            .in1(N__63280),
            .in2(N__66120),
            .in3(N__56707),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71125),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_696_LC_17_13_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_696_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_696_LC_17_13_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_696_LC_17_13_0  (
            .in0(N__44893),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52206),
            .lcout(\c0.n16_adj_3489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_575_LC_17_13_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_575_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_575_LC_17_13_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i9_4_lut_adj_575_LC_17_13_1  (
            .in0(N__42757),
            .in1(N__41566),
            .in2(N__39628),
            .in3(N__41755),
            .lcout(),
            .ltout(\c0.n20_adj_3437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_582_LC_17_13_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_582_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_582_LC_17_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_582_LC_17_13_2  (
            .in0(N__41647),
            .in1(N__38669),
            .in2(N__38638),
            .in3(N__39304),
            .lcout(n21222),
            .ltout(n21222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i6_LC_17_13_3 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i6_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i6_LC_17_13_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.control_mode_i0_i6_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__38631),
            .in2(N__38635),
            .in3(N__54895),
            .lcout(control_mode_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71112),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i2_LC_17_13_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i2_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i2_LC_17_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i2_LC_17_13_4  (
            .in0(N__38619),
            .in1(N__60412),
            .in2(_gnd_net_),
            .in3(N__41086),
            .lcout(control_mode_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71112),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i4_LC_17_13_5 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i4_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i4_LC_17_13_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.control_mode_i0_i4_LC_17_13_5  (
            .in0(N__38751),
            .in1(_gnd_net_),
            .in2(N__41097),
            .in3(N__60931),
            .lcout(control_mode_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71112),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i3_LC_17_13_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i3_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i3_LC_17_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i3_LC_17_13_6  (
            .in0(N__38733),
            .in1(N__61231),
            .in2(_gnd_net_),
            .in3(N__41087),
            .lcout(control_mode_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71112),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i7_LC_17_13_7 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i7_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i7_LC_17_13_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.control_mode_i0_i7_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__38715),
            .in2(N__41098),
            .in3(N__54691),
            .lcout(control_mode_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71112),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i145_LC_17_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i145_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i145_LC_17_14_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i145_LC_17_14_0  (
            .in0(N__51171),
            .in1(N__63944),
            .in2(_gnd_net_),
            .in3(N__65070),
            .lcout(data_in_frame_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71095),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_17_14_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_17_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__45141),
            .in2(_gnd_net_),
            .in3(N__63862),
            .lcout(\c0.n6_adj_3005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_225_LC_17_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_225_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_225_LC_17_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_225_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__41551),
            .in2(_gnd_net_),
            .in3(N__44545),
            .lcout(\c0.n9 ),
            .ltout(\c0.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_908_LC_17_14_3 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_908_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_908_LC_17_14_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_908_LC_17_14_3  (
            .in0(N__52827),
            .in1(N__45459),
            .in2(N__38704),
            .in3(N__45715),
            .lcout(),
            .ltout(\c0.n16_adj_3008_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_233_LC_17_14_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_233_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_233_LC_17_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_233_LC_17_14_4  (
            .in0(N__56313),
            .in1(N__41190),
            .in2(N__38701),
            .in3(N__43023),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_693_LC_17_14_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_693_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_693_LC_17_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_693_LC_17_14_5  (
            .in0(N__43024),
            .in1(N__56314),
            .in2(N__41194),
            .in3(N__38698),
            .lcout(\c0.n19449 ),
            .ltout(\c0.n19449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_694_LC_17_14_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_694_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_694_LC_17_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_694_LC_17_14_6  (
            .in0(N__45460),
            .in1(N__50904),
            .in2(N__39091),
            .in3(N__45640),
            .lcout(\c0.n12218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i0_LC_17_14_7 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i0_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i0_LC_17_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i0_LC_17_14_7  (
            .in0(N__39087),
            .in1(N__55053),
            .in2(_gnd_net_),
            .in3(N__41094),
            .lcout(control_mode_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71095),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_adj_489_LC_17_15_0 .C_ON=1'b0;
    defparam \c0.i24_3_lut_adj_489_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_adj_489_LC_17_15_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \c0.i24_3_lut_adj_489_LC_17_15_0  (
            .in0(N__39060),
            .in1(N__38997),
            .in2(_gnd_net_),
            .in3(N__38837),
            .lcout(\c0.n13_adj_3016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i139_LC_17_15_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i139_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i139_LC_17_15_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i139_LC_17_15_2  (
            .in0(N__68521),
            .in1(N__63357),
            .in2(N__71792),
            .in3(N__68348),
            .lcout(\c0.data_in_frame_17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71083),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_17_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_17_15_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_17_15_3  (
            .in0(N__38802),
            .in1(N__44127),
            .in2(N__53118),
            .in3(N__42132),
            .lcout(\c0.n19111 ),
            .ltout(\c0.n19111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i104_LC_17_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i104_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i104_LC_17_15_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i104_LC_17_15_4  (
            .in0(N__66125),
            .in1(N__57071),
            .in2(N__38770),
            .in3(N__72295),
            .lcout(\c0.data_in_frame_12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71083),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_226_LC_17_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_226_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_226_LC_17_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_226_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__38767),
            .in2(_gnd_net_),
            .in3(N__55618),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_17_15_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_17_15_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_17_15_7  (
            .in0(N__41533),
            .in1(N__68522),
            .in2(N__56080),
            .in3(N__56200),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71083),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_17_16_1 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_17_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_17_16_1  (
            .in0(N__50077),
            .in1(N__47509),
            .in2(N__56359),
            .in3(N__51109),
            .lcout(),
            .ltout(\c0.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_17_16_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_17_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_LC_17_16_2  (
            .in0(N__39112),
            .in1(N__39106),
            .in2(N__39100),
            .in3(N__54467),
            .lcout(\c0.n12026 ),
            .ltout(\c0.n12026_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_230_LC_17_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_230_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_230_LC_17_16_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_230_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39097),
            .in3(N__45137),
            .lcout(\c0.n5_adj_3003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_403_LC_17_16_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_403_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_403_LC_17_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_403_LC_17_16_4  (
            .in0(N__51623),
            .in1(N__48082),
            .in2(N__64723),
            .in3(N__52020),
            .lcout(\c0.n32_adj_3236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i150_LC_17_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i150_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i150_LC_17_16_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i150_LC_17_16_5  (
            .in0(N__67982),
            .in1(N__63948),
            .in2(_gnd_net_),
            .in3(N__44892),
            .lcout(data_in_frame_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71070),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i212_LC_17_16_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i212_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i212_LC_17_16_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i212_LC_17_16_7  (
            .in0(N__69314),
            .in1(N__66754),
            .in2(N__67562),
            .in3(N__62845),
            .lcout(\c0.data_in_frame_26_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71070),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_386_LC_17_17_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_386_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_386_LC_17_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_386_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__64834),
            .in2(_gnd_net_),
            .in3(N__72858),
            .lcout(\c0.n11_adj_3219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_17_17_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_17_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i3_2_lut_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__44717),
            .in2(_gnd_net_),
            .in3(N__48402),
            .lcout(\c0.n10 ),
            .ltout(\c0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_897_LC_17_17_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_897_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_897_LC_17_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_897_LC_17_17_2  (
            .in0(N__41218),
            .in1(N__65849),
            .in2(N__39094),
            .in3(N__47773),
            .lcout(\c0.n12_adj_3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_232_LC_17_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_232_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_232_LC_17_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_232_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__57725),
            .in2(_gnd_net_),
            .in3(N__48650),
            .lcout(\c0.n19551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_adj_685_LC_17_17_5 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_adj_685_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_adj_685_LC_17_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_adj_685_LC_17_17_5  (
            .in0(N__52345),
            .in1(N__44718),
            .in2(N__68364),
            .in3(N__47692),
            .lcout(\c0.n20_adj_3487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_571_LC_17_17_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_571_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_571_LC_17_17_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_571_LC_17_17_6  (
            .in0(N__41518),
            .in1(N__41734),
            .in2(N__45985),
            .in3(N__43348),
            .lcout(\c0.n21104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i112_LC_17_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i112_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i112_LC_17_17_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i112_LC_17_17_7  (
            .in0(N__66060),
            .in1(N__71941),
            .in2(N__56017),
            .in3(N__72283),
            .lcout(\c0.data_in_frame_13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71047),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1998_2_lut_LC_17_18_0 .C_ON=1'b0;
    defparam \c0.rx.i1998_2_lut_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1998_2_lut_LC_17_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i1998_2_lut_LC_17_18_0  (
            .in0(N__43801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39343),
            .lcout(),
            .ltout(n3846_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_17_18_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_17_18_1 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_17_18_1  (
            .in0(N__43849),
            .in1(N__39402),
            .in2(N__39295),
            .in3(N__39375),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71071),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_817_LC_17_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_817_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_817_LC_17_18_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_817_LC_17_18_2  (
            .in0(N__68355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68299),
            .lcout(\c0.n5_adj_3220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_17_18_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_17_18_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_17_18_3  (
            .in0(N__39344),
            .in1(N__39401),
            .in2(_gnd_net_),
            .in3(N__39374),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71071),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4_4_lut_LC_17_18_4 .C_ON=1'b0;
    defparam \c0.rx.i4_4_lut_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4_4_lut_LC_17_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i4_4_lut_LC_17_18_4  (
            .in0(N__39291),
            .in1(N__39250),
            .in2(N__39143),
            .in3(N__39243),
            .lcout(\c0.rx.r_SM_Main_2_N_2479_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_96_i4_2_lut_LC_17_18_5 .C_ON=1'b0;
    defparam \c0.rx.equal_96_i4_2_lut_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_96_i4_2_lut_LC_17_18_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.equal_96_i4_2_lut_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__43840),
            .in2(_gnd_net_),
            .in3(N__43800),
            .lcout(n4_adj_3595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_17_18_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_17_18_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__39195),
            .in2(_gnd_net_),
            .in3(N__39163),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71071),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_207_LC_17_18_7 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_207_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_207_LC_17_18_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_adj_207_LC_17_18_7  (
            .in0(N__39342),
            .in1(N__43839),
            .in2(_gnd_net_),
            .in3(N__43799),
            .lcout(\c0.rx.n15860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i12_LC_17_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_17_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_17_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__41496),
            .in2(_gnd_net_),
            .in3(N__40551),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71084),
            .ce(),
            .sr(N__41284));
    defparam \c0.data_in_frame_0__i229_LC_17_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i229_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i229_LC_17_20_0 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i229_LC_17_20_0  (
            .in0(N__72766),
            .in1(N__41578),
            .in2(N__66850),
            .in3(N__67144),
            .lcout(\c0.data_in_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71096),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_613_LC_17_20_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_613_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_613_LC_17_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_613_LC_17_20_2  (
            .in0(N__65693),
            .in1(N__59115),
            .in2(N__41604),
            .in3(N__39418),
            .lcout(\c0.n13_adj_3463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i49_4_lut_LC_17_20_4 .C_ON=1'b0;
    defparam \c0.i49_4_lut_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i49_4_lut_LC_17_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i49_4_lut_LC_17_20_4  (
            .in0(N__58495),
            .in1(N__58276),
            .in2(N__41275),
            .in3(N__48460),
            .lcout(\c0.n100_adj_3403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i221_LC_17_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i221_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i221_LC_17_20_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i221_LC_17_20_5  (
            .in0(N__66917),
            .in1(N__72767),
            .in2(N__48830),
            .in3(N__64585),
            .lcout(\c0.data_in_frame_27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71096),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_17_20_6 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_17_20_6 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_17_20_6  (
            .in0(N__39406),
            .in1(N__43790),
            .in2(N__39382),
            .in3(N__39345),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71096),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_3_lut_4_lut_adj_587_LC_17_21_0 .C_ON=1'b0;
    defparam \c0.i14_2_lut_3_lut_4_lut_adj_587_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_3_lut_4_lut_adj_587_LC_17_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_2_lut_3_lut_4_lut_adj_587_LC_17_21_0  (
            .in0(N__65527),
            .in1(N__63778),
            .in2(N__63583),
            .in3(N__43093),
            .lcout(\c0.n34_adj_3096 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_439_LC_17_21_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_439_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_439_LC_17_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_439_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__48789),
            .in2(_gnd_net_),
            .in3(N__41721),
            .lcout(),
            .ltout(\c0.n22_adj_3276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_441_LC_17_21_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_441_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_441_LC_17_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_441_LC_17_21_2  (
            .in0(N__41977),
            .in1(N__41706),
            .in2(N__39307),
            .in3(N__45766),
            .lcout(),
            .ltout(\c0.n36_adj_3277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_442_LC_17_21_3 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_442_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_442_LC_17_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_442_LC_17_21_3  (
            .in0(N__49024),
            .in1(N__51760),
            .in2(N__39643),
            .in3(N__45780),
            .lcout(),
            .ltout(\c0.n20415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_537_LC_17_21_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_537_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_537_LC_17_21_4 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i3_4_lut_adj_537_LC_17_21_4  (
            .in0(N__46027),
            .in1(N__59302),
            .in2(N__39640),
            .in3(N__41674),
            .lcout(),
            .ltout(\c0.n14_adj_3407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_544_LC_17_21_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_544_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_544_LC_17_21_5 .LUT_INIT=16'b1111101111110111;
    LogicCell40 \c0.i7_4_lut_adj_544_LC_17_21_5  (
            .in0(N__43315),
            .in1(N__39679),
            .in2(N__39637),
            .in3(N__39634),
            .lcout(\c0.n18_adj_3412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_17_22_0 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_17_22_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_17_22_0  (
            .in0(N__66631),
            .in1(N__53537),
            .in2(N__49303),
            .in3(N__52672),
            .lcout(\c0.n20300 ),
            .ltout(\c0.n20300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_350_LC_17_22_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_350_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_350_LC_17_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_350_LC_17_22_1  (
            .in0(N__49230),
            .in1(N__52567),
            .in2(N__39610),
            .in3(N__57862),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_530_LC_17_22_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_530_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_530_LC_17_22_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_530_LC_17_22_2  (
            .in0(N__59688),
            .in1(N__49231),
            .in2(N__39607),
            .in3(N__45935),
            .lcout(\c0.n20370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i186_LC_17_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i186_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i186_LC_17_22_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i186_LC_17_22_3  (
            .in0(N__66632),
            .in1(N__53702),
            .in2(_gnd_net_),
            .in3(N__71548),
            .lcout(data_in_frame_23_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71126),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1213_2_lut_LC_17_22_4 .C_ON=1'b0;
    defparam \c0.i1213_2_lut_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1213_2_lut_LC_17_22_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.i1213_2_lut_LC_17_22_4  (
            .in0(N__39576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42504),
            .lcout(\c0.n3235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_LC_17_22_5 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_LC_17_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_2_lut_3_lut_LC_17_22_5  (
            .in0(N__64886),
            .in1(N__44897),
            .in2(_gnd_net_),
            .in3(N__48381),
            .lcout(\c0.n40_adj_3374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i133_LC_17_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i133_LC_17_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i133_LC_17_22_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i133_LC_17_22_6  (
            .in0(N__72774),
            .in1(N__65598),
            .in2(_gnd_net_),
            .in3(N__45612),
            .lcout(data_in_frame_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71126),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_850_LC_17_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_850_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_850_LC_17_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_850_LC_17_23_0  (
            .in0(N__41942),
            .in1(N__49458),
            .in2(N__49785),
            .in3(N__53259),
            .lcout(\c0.n17947 ),
            .ltout(\c0.n17947_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_532_LC_17_23_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_532_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_532_LC_17_23_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_3_lut_adj_532_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__39703),
            .in2(N__39682),
            .in3(N__70405),
            .lcout(\c0.n20793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i227_LC_17_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i227_LC_17_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i227_LC_17_23_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i227_LC_17_23_2  (
            .in0(N__68646),
            .in1(N__67178),
            .in2(N__59211),
            .in3(N__66952),
            .lcout(\c0.data_in_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71143),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i213_LC_17_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i213_LC_17_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i213_LC_17_23_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i213_LC_17_23_4  (
            .in0(N__72737),
            .in1(N__66948),
            .in2(N__41949),
            .in3(N__62838),
            .lcout(\c0.data_in_frame_26_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71143),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_407_LC_17_23_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_407_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_407_LC_17_23_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_adj_407_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__39739),
            .in2(_gnd_net_),
            .in3(N__39865),
            .lcout(),
            .ltout(\c0.n10_adj_3242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_410_LC_17_23_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_410_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_410_LC_17_23_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i7_4_lut_adj_410_LC_17_23_6  (
            .in0(N__43906),
            .in1(N__52942),
            .in2(N__39670),
            .in3(N__39649),
            .lcout(\c0.n11446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i214_LC_17_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i214_LC_17_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i214_LC_17_23_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i214_LC_17_23_7  (
            .in0(N__62837),
            .in1(N__67987),
            .in2(N__66977),
            .in3(N__49781),
            .lcout(\c0.data_in_frame_26_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71143),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_408_LC_17_24_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_408_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_408_LC_17_24_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i6_4_lut_adj_408_LC_17_24_0  (
            .in0(N__39844),
            .in1(N__39665),
            .in2(N__39828),
            .in3(N__40025),
            .lcout(\c0.n14_adj_3243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_397_LC_17_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_397_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_397_LC_17_24_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_397_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__47006),
            .in2(_gnd_net_),
            .in3(N__41631),
            .lcout(\c0.n105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3__5178_LC_17_24_3 .C_ON=1'b0;
    defparam \c0.data_in_2__3__5178_LC_17_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3__5178_LC_17_24_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_2__3__5178_LC_17_24_3  (
            .in0(N__40026),
            .in1(_gnd_net_),
            .in2(N__53224),
            .in3(N__39868),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71158),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1__5172_LC_17_24_5 .C_ON=1'b0;
    defparam \c0.data_in_3__1__5172_LC_17_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1__5172_LC_17_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__1__5172_LC_17_24_5  (
            .in0(N__53188),
            .in1(N__71505),
            .in2(_gnd_net_),
            .in3(N__39845),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71158),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_916_LC_17_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_916_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_916_LC_17_24_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_916_LC_17_24_6  (
            .in0(N__71777),
            .in1(N__64393),
            .in2(_gnd_net_),
            .in3(N__59455),
            .lcout(n19126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7__5190_LC_17_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0__7__5190_LC_17_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7__5190_LC_17_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__7__5190_LC_17_24_7  (
            .in0(N__53187),
            .in1(N__39824),
            .in2(_gnd_net_),
            .in3(N__43942),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71158),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_398_LC_17_25_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_398_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_398_LC_17_25_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i7_4_lut_adj_398_LC_17_25_0  (
            .in0(N__39807),
            .in1(N__39914),
            .in2(N__39769),
            .in3(N__41895),
            .lcout(\c0.n18_adj_3229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_415_LC_17_25_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_415_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_415_LC_17_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_415_LC_17_25_1  (
            .in0(N__42605),
            .in1(N__41927),
            .in2(N__49744),
            .in3(N__39961),
            .lcout(),
            .ltout(\c0.n21108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_416_LC_17_25_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_416_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_416_LC_17_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_416_LC_17_25_2  (
            .in0(N__39765),
            .in1(N__41853),
            .in2(N__39754),
            .in3(N__39924),
            .lcout(\c0.n12_adj_3248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_418_LC_17_25_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_418_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_418_LC_17_25_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i8_4_lut_adj_418_LC_17_25_3  (
            .in0(N__39925),
            .in1(N__39745),
            .in2(N__52956),
            .in3(N__40032),
            .lcout(\c0.n20_adj_3250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3__5186_LC_17_25_4 .C_ON=1'b0;
    defparam \c0.data_in_1__3__5186_LC_17_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3__5186_LC_17_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__3__5186_LC_17_25_4  (
            .in0(N__40033),
            .in1(N__53219),
            .in2(_gnd_net_),
            .in3(N__40008),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71167),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4__5177_LC_17_25_5 .C_ON=1'b0;
    defparam \c0.data_in_2__4__5177_LC_17_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4__5177_LC_17_25_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_2__4__5177_LC_17_25_5  (
            .in0(N__53218),
            .in1(N__47033),
            .in2(_gnd_net_),
            .in3(N__43981),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71167),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2__5179_LC_17_25_6 .C_ON=1'b0;
    defparam \c0.data_in_2__2__5179_LC_17_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2__5179_LC_17_25_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_2__2__5179_LC_17_25_6  (
            .in0(N__41928),
            .in1(N__53220),
            .in2(_gnd_net_),
            .in3(N__39915),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71167),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_404_LC_17_25_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_404_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_404_LC_17_25_7 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i4_4_lut_adj_404_LC_17_25_7  (
            .in0(N__42604),
            .in1(N__47032),
            .in2(N__39982),
            .in3(N__39960),
            .lcout(\c0.n10_adj_3238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_412_LC_17_26_0 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_412_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_412_LC_17_26_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i5_2_lut_adj_412_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__40573),
            .in2(_gnd_net_),
            .in3(N__42536),
            .lcout(\c0.n16_adj_3247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_413_LC_17_26_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_413_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_413_LC_17_26_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_413_LC_17_26_2  (
            .in0(N__52920),
            .in1(N__39940),
            .in2(N__39916),
            .in3(N__42550),
            .lcout(),
            .ltout(\c0.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_414_LC_17_26_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_414_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_414_LC_17_26_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i10_4_lut_adj_414_LC_17_26_3  (
            .in0(N__41623),
            .in1(N__42628),
            .in2(N__39934),
            .in3(N__39931),
            .lcout(\c0.n11311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7__5166_LC_17_26_4 .C_ON=1'b0;
    defparam \c0.data_in_3__7__5166_LC_17_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7__5166_LC_17_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__7__5166_LC_17_26_4  (
            .in0(N__53222),
            .in1(N__72292),
            .in2(_gnd_net_),
            .in3(N__41624),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71178),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2__5171_LC_17_26_5 .C_ON=1'b0;
    defparam \c0.data_in_3__2__5171_LC_17_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2__5171_LC_17_26_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__2__5171_LC_17_26_5  (
            .in0(N__68644),
            .in1(N__53223),
            .in2(_gnd_net_),
            .in3(N__39913),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71178),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5__5192_LC_17_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0__5__5192_LC_17_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5__5192_LC_17_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__5__5192_LC_17_26_6  (
            .in0(N__53221),
            .in1(N__41854),
            .in2(_gnd_net_),
            .in3(N__40574),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71178),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i18_LC_17_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_17_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_17_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__40317),
            .in2(_gnd_net_),
            .in3(N__40552),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71189),
            .ce(),
            .sr(N__40297));
    defparam \c0.rx.equal_94_i4_2_lut_LC_18_5_6 .C_ON=1'b0;
    defparam \c0.rx.equal_94_i4_2_lut_LC_18_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_94_i4_2_lut_LC_18_5_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.equal_94_i4_2_lut_LC_18_5_6  (
            .in0(_gnd_net_),
            .in1(N__43870),
            .in2(_gnd_net_),
            .in3(N__43818),
            .lcout(n4_adj_3579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_65_i9_2_lut_3_lut_LC_18_7_2 .C_ON=1'b0;
    defparam \c0.equal_65_i9_2_lut_3_lut_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.equal_65_i9_2_lut_3_lut_LC_18_7_2 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.equal_65_i9_2_lut_3_lut_LC_18_7_2  (
            .in0(N__60252),
            .in1(N__59985),
            .in2(_gnd_net_),
            .in3(N__60104),
            .lcout(\c0.n9_adj_3025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_18_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_18_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_18_7_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i25_LC_18_7_4  (
            .in0(N__65147),
            .in1(N__61688),
            .in2(N__61449),
            .in3(N__47598),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71200),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_525_LC_18_7_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_525_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_525_LC_18_7_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_525_LC_18_7_7  (
            .in0(N__40288),
            .in1(N__40175),
            .in2(N__40118),
            .in3(N__49655),
            .lcout(\c0.n12_adj_3265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_703_LC_18_8_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_703_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_703_LC_18_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_703_LC_18_8_0  (
            .in0(N__54058),
            .in1(N__47596),
            .in2(N__47344),
            .in3(N__55183),
            .lcout(\c0.n20224 ),
            .ltout(\c0.n20224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_274_LC_18_8_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_274_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_274_LC_18_8_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i3_2_lut_adj_274_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40039),
            .in3(N__41143),
            .lcout(),
            .ltout(\c0.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_277_LC_18_8_2 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_277_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_277_LC_18_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_277_LC_18_8_2  (
            .in0(N__42649),
            .in1(N__40621),
            .in2(N__40036),
            .in3(N__50076),
            .lcout(\c0.n20246 ),
            .ltout(\c0.n20246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_286_LC_18_8_3 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_286_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_286_LC_18_8_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i4_2_lut_adj_286_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40642),
            .in3(N__47259),
            .lcout(\c0.n12_adj_3049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_810_LC_18_8_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_810_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_810_LC_18_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i3_2_lut_adj_810_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__61226),
            .in2(_gnd_net_),
            .in3(N__60411),
            .lcout(\c0.n24_adj_3327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_LC_18_8_5 .C_ON=1'b0;
    defparam \c0.i7_2_lut_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_LC_18_8_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i7_2_lut_LC_18_8_5  (
            .in0(N__47597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50604),
            .lcout(\c0.n23_adj_3039 ),
            .ltout(\c0.n23_adj_3039_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_941_LC_18_8_6 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_941_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_941_LC_18_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_941_LC_18_8_6  (
            .in0(N__41002),
            .in1(N__42717),
            .in2(N__40630),
            .in3(N__42690),
            .lcout(\c0.n42_adj_3560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_275_LC_18_8_7 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_275_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_275_LC_18_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_275_LC_18_8_7  (
            .in0(N__40627),
            .in1(N__43230),
            .in2(N__42718),
            .in3(N__41001),
            .lcout(\c0.n30_adj_3042 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i37_LC_18_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i37_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i37_LC_18_9_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i37_LC_18_9_0  (
            .in0(N__44117),
            .in1(N__61596),
            .in2(N__54266),
            .in3(N__72612),
            .lcout(\c0.data_in_frame_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71181),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__2__5204_LC_18_9_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__2__5204_LC_18_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__2__5204_LC_18_9_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \c0.data_out_frame_29__2__5204_LC_18_9_1  (
            .in0(N__55185),
            .in1(N__46907),
            .in2(_gnd_net_),
            .in3(N__40614),
            .lcout(data_out_frame_29_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71181),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_550_LC_18_9_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_550_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_550_LC_18_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_550_LC_18_9_2  (
            .in0(N__49917),
            .in1(N__54876),
            .in2(_gnd_net_),
            .in3(N__42970),
            .lcout(),
            .ltout(\c0.n18428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_593_LC_18_9_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_593_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_593_LC_18_9_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i12_4_lut_adj_593_LC_18_9_3  (
            .in0(N__49828),
            .in1(N__44506),
            .in2(N__40600),
            .in3(N__47911),
            .lcout(\c0.n29_adj_3446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__2__5212_LC_18_9_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__2__5212_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__2__5212_LC_18_9_4 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \c0.data_out_frame_28__2__5212_LC_18_9_4  (
            .in0(N__46905),
            .in1(N__40591),
            .in2(N__46300),
            .in3(N__56853),
            .lcout(data_out_frame_28_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71181),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__1__5213_LC_18_9_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__1__5213_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__1__5213_LC_18_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_frame_28__1__5213_LC_18_9_5  (
            .in0(N__40957),
            .in1(N__46906),
            .in2(_gnd_net_),
            .in3(N__46287),
            .lcout(data_out_frame_28_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71181),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i40_LC_18_9_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i40_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i40_LC_18_9_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i40_LC_18_9_6  (
            .in0(N__44118),
            .in1(N__72231),
            .in2(N__51282),
            .in3(N__61597),
            .lcout(\c0.data_in_frame_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71181),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_704_LC_18_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_704_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_704_LC_18_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_704_LC_18_9_7  (
            .in0(N__51399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51266),
            .lcout(\c0.n5_adj_3044 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_922_LC_18_10_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_922_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_922_LC_18_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_922_LC_18_10_0  (
            .in0(N__46283),
            .in1(N__42817),
            .in2(N__42868),
            .in3(N__42823),
            .lcout(\c0.data_out_frame_28__0__N_708 ),
            .ltout(\c0.data_out_frame_28__0__N_708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__1__5205_LC_18_10_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__1__5205_LC_18_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__1__5205_LC_18_10_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.data_out_frame_29__1__5205_LC_18_10_1  (
            .in0(N__50348),
            .in1(_gnd_net_),
            .in2(N__40984),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71169),
            .ce(N__46858),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__0__5206_LC_18_10_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__0__5206_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__0__5206_LC_18_10_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.data_out_frame_29__0__5206_LC_18_10_2  (
            .in0(N__55165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40981),
            .lcout(\c0.data_out_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71169),
            .ce(N__46858),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_18_10_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_18_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_18_10_4  (
            .in0(N__40963),
            .in1(N__40956),
            .in2(_gnd_net_),
            .in3(N__40926),
            .lcout(\c0.n26_adj_3103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_794_LC_18_10_5 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_794_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_794_LC_18_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_794_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__55163),
            .in2(_gnd_net_),
            .in3(N__62127),
            .lcout(\c0.n14_adj_3525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_808_LC_18_10_6 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_808_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_808_LC_18_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3_2_lut_adj_808_LC_18_10_6  (
            .in0(N__62126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54383),
            .lcout(\c0.n11_adj_3507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_241_LC_18_10_7 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_241_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_241_LC_18_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_241_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__55164),
            .in2(_gnd_net_),
            .in3(N__54134),
            .lcout(\c0.n12_adj_3015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_747_LC_18_11_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_747_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_747_LC_18_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_747_LC_18_11_0  (
            .in0(N__47545),
            .in1(N__54410),
            .in2(_gnd_net_),
            .in3(N__50554),
            .lcout(\c0.n20209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_781_LC_18_11_1 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_781_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_781_LC_18_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_781_LC_18_11_1  (
            .in0(N__50496),
            .in1(N__54560),
            .in2(N__50086),
            .in3(N__54423),
            .lcout(\c0.n20204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_adj_304_LC_18_11_2 .C_ON=1'b0;
    defparam \c0.i8_2_lut_adj_304_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_adj_304_LC_18_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i8_2_lut_adj_304_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__41124),
            .in2(_gnd_net_),
            .in3(N__51386),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_18_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_18_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_18_11_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i6_LC_18_11_3  (
            .in0(N__61723),
            .in1(N__67979),
            .in2(N__50582),
            .in3(N__55888),
            .lcout(data_in_frame_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71159),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_600_LC_18_11_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_600_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_600_LC_18_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_600_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__50641),
            .in2(_gnd_net_),
            .in3(N__55179),
            .lcout(\c0.n19217 ),
            .ltout(\c0.n19217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_3_lut_LC_18_11_5 .C_ON=1'b0;
    defparam \c0.i33_3_lut_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i33_3_lut_LC_18_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i33_3_lut_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__40995),
            .in2(N__41005),
            .in3(N__47615),
            .lcout(\c0.n85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_18_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_18_11_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i5_LC_18_11_6  (
            .in0(N__72649),
            .in1(N__55887),
            .in2(N__54459),
            .in3(N__61724),
            .lcout(data_in_frame_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71159),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_LC_18_11_7 .C_ON=1'b0;
    defparam \c0.i14_2_lut_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_LC_18_11_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i14_2_lut_LC_18_11_7  (
            .in0(N__54411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47546),
            .lcout(\c0.n66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_601_LC_18_12_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_601_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_601_LC_18_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_601_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__47614),
            .in2(_gnd_net_),
            .in3(N__47547),
            .lcout(\c0.n23_adj_3076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i1_LC_18_12_1 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i1_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i1_LC_18_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i1_LC_18_12_1  (
            .in0(N__41049),
            .in1(N__54135),
            .in2(_gnd_net_),
            .in3(N__41095),
            .lcout(control_mode_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71144),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_18_12_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_18_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_18_12_3  (
            .in0(N__41038),
            .in1(N__55510),
            .in2(N__43179),
            .in3(N__54733),
            .lcout(\c0.n20321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_18_12_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_18_12_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_18_12_4  (
            .in0(N__61779),
            .in1(N__61448),
            .in2(N__50679),
            .in3(N__71496),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71144),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_829_LC_18_12_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_829_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_829_LC_18_12_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_829_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__50550),
            .in2(_gnd_net_),
            .in3(N__54395),
            .lcout(\c0.n15_adj_3543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i93_LC_18_12_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i93_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i93_LC_18_12_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i93_LC_18_12_6  (
            .in0(N__72677),
            .in1(N__64551),
            .in2(N__50984),
            .in3(N__66050),
            .lcout(\c0.data_in_frame_11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71144),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_18_12_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_18_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_18_12_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i23_LC_18_12_7  (
            .in0(N__47548),
            .in1(N__68980),
            .in2(N__44253),
            .in3(N__61780),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71144),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_18_13_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_18_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_18_13_0  (
            .in0(N__62255),
            .in1(N__47921),
            .in2(_gnd_net_),
            .in3(N__56650),
            .lcout(\c0.n19176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_4_lut_adj_714_LC_18_13_1 .C_ON=1'b0;
    defparam \c0.i12_3_lut_4_lut_adj_714_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_4_lut_adj_714_LC_18_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_3_lut_4_lut_adj_714_LC_18_13_1  (
            .in0(N__56651),
            .in1(N__41131),
            .in2(N__56452),
            .in3(N__42672),
            .lcout(),
            .ltout(\c0.n32_adj_3493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_849_LC_18_13_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_849_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_849_LC_18_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_849_LC_18_13_2  (
            .in0(N__42901),
            .in1(N__61284),
            .in2(N__41032),
            .in3(N__42933),
            .lcout(),
            .ltout(\c0.n36_adj_3547_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_856_LC_18_13_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_856_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_856_LC_18_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_856_LC_18_13_3  (
            .in0(N__56703),
            .in1(N__54556),
            .in2(N__41182),
            .in3(N__54442),
            .lcout(),
            .ltout(\c0.n38_adj_3548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_861_LC_18_13_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_861_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_861_LC_18_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_861_LC_18_13_4  (
            .in0(N__41179),
            .in1(N__41149),
            .in2(N__41167),
            .in3(N__41164),
            .lcout(\c0.n18443 ),
            .ltout(\c0.n18443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_LC_18_13_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_LC_18_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_2_lut_3_lut_LC_18_13_5  (
            .in0(N__44734),
            .in1(_gnd_net_),
            .in2(N__41152),
            .in3(N__64633),
            .lcout(\c0.n24_adj_3335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_298_LC_18_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_298_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_298_LC_18_14_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_298_LC_18_14_0  (
            .in0(N__50157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50182),
            .lcout(\c0.n4_adj_3071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_adj_784_LC_18_14_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_adj_784_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_adj_784_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_2_lut_3_lut_adj_784_LC_18_14_1  (
            .in0(N__51338),
            .in1(N__50349),
            .in2(_gnd_net_),
            .in3(N__55052),
            .lcout(\c0.n25_adj_3495 ),
            .ltout(\c0.n25_adj_3495_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_4_lut_LC_18_14_2 .C_ON=1'b0;
    defparam \c0.i20_3_lut_4_lut_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_4_lut_LC_18_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_3_lut_4_lut_LC_18_14_2  (
            .in0(N__41142),
            .in1(N__42671),
            .in2(N__41101),
            .in3(N__47428),
            .lcout(\c0.n44_adj_3117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i222_LC_18_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i222_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i222_LC_18_14_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i222_LC_18_14_3  (
            .in0(N__67920),
            .in1(N__64577),
            .in2(N__48785),
            .in3(N__66962),
            .lcout(\c0.data_in_frame_27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71113),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i137_LC_18_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i137_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i137_LC_18_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i137_LC_18_14_4  (
            .in0(N__71786),
            .in1(N__63354),
            .in2(N__48366),
            .in3(N__65239),
            .lcout(\c0.data_in_frame_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71113),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i140_LC_18_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i140_LC_18_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i140_LC_18_14_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i140_LC_18_14_5  (
            .in0(N__63353),
            .in1(N__71787),
            .in2(N__69444),
            .in3(N__68274),
            .lcout(\c0.data_in_frame_17_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71113),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i206_LC_18_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i206_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i206_LC_18_14_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i206_LC_18_14_6  (
            .in0(N__59719),
            .in1(N__63355),
            .in2(N__66978),
            .in3(N__67919),
            .lcout(\c0.data_in_frame_25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71113),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_588_LC_18_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_588_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_588_LC_18_14_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_588_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__44220),
            .in2(_gnd_net_),
            .in3(N__59480),
            .lcout(\c0.n19134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_819_LC_18_15_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_819_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_819_LC_18_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_819_LC_18_15_0  (
            .in0(N__43275),
            .in1(N__44472),
            .in2(N__63575),
            .in3(N__58466),
            .lcout(\c0.n20_adj_3539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_744_LC_18_15_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_744_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_744_LC_18_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_744_LC_18_15_1  (
            .in0(N__44631),
            .in1(N__62418),
            .in2(N__44480),
            .in3(N__43274),
            .lcout(\c0.n10_adj_3514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_18_15_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_18_15_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_LC_18_15_2  (
            .in0(N__57412),
            .in1(N__43126),
            .in2(N__47653),
            .in3(N__41200),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_602_LC_18_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_602_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_602_LC_18_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_602_LC_18_15_3  (
            .in0(N__62968),
            .in1(N__47802),
            .in2(_gnd_net_),
            .in3(N__61879),
            .lcout(\c0.n6_adj_3453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i129_LC_18_15_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i129_LC_18_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i129_LC_18_15_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i129_LC_18_15_4  (
            .in0(N__65238),
            .in1(N__65595),
            .in2(_gnd_net_),
            .in3(N__62969),
            .lcout(data_in_frame_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71097),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i130_LC_18_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i130_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i130_LC_18_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i130_LC_18_15_5  (
            .in0(N__65594),
            .in1(N__71486),
            .in2(_gnd_net_),
            .in3(N__47803),
            .lcout(data_in_frame_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71097),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_18_15_6 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_18_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_18_15_6  (
            .in0(N__62890),
            .in1(N__47925),
            .in2(N__49582),
            .in3(N__57045),
            .lcout(\c0.n18_adj_3369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_LC_18_15_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_LC_18_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__55669),
            .in2(_gnd_net_),
            .in3(N__52092),
            .lcout(\c0.n17849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_821_LC_18_16_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_821_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_821_LC_18_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_821_LC_18_16_0  (
            .in0(N__41254),
            .in1(N__44584),
            .in2(N__56878),
            .in3(N__50113),
            .lcout(\c0.n19474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_927_LC_18_16_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_927_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_927_LC_18_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_927_LC_18_16_1  (
            .in0(N__43276),
            .in1(N__44479),
            .in2(N__41233),
            .in3(N__62419),
            .lcout(),
            .ltout(\c0.n12_adj_3001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_227_LC_18_16_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_227_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_227_LC_18_16_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_227_LC_18_16_2  (
            .in0(N__57152),
            .in1(N__44632),
            .in2(N__41248),
            .in3(N__52275),
            .lcout(\c0.n20403 ),
            .ltout(\c0.n20403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_745_LC_18_16_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_745_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_745_LC_18_16_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_745_LC_18_16_3  (
            .in0(N__43277),
            .in1(N__48429),
            .in2(N__41245),
            .in3(N__41216),
            .lcout(),
            .ltout(\c0.n20398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_746_LC_18_16_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_746_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_746_LC_18_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_746_LC_18_16_4  (
            .in0(N__57153),
            .in1(N__41242),
            .in2(N__41236),
            .in3(N__41232),
            .lcout(\c0.n10_adj_3445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_639_LC_18_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_639_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_639_LC_18_16_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_639_LC_18_16_5  (
            .in0(N__64769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68289),
            .lcout(\c0.n12134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_596_LC_18_16_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_596_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_596_LC_18_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_596_LC_18_16_6  (
            .in0(N__41217),
            .in1(N__45637),
            .in2(N__45458),
            .in3(N__44633),
            .lcout(\c0.n20_adj_3448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_2_lut_3_lut_adj_678_LC_18_17_0 .C_ON=1'b0;
    defparam \c0.i19_2_lut_3_lut_adj_678_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_2_lut_3_lut_adj_678_LC_18_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i19_2_lut_3_lut_adj_678_LC_18_17_0  (
            .in0(N__68374),
            .in1(N__52346),
            .in2(_gnd_net_),
            .in3(N__52171),
            .lcout(\c0.n36_adj_3267 ),
            .ltout(\c0.n36_adj_3267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i35_2_lut_LC_18_17_1 .C_ON=1'b0;
    defparam \c0.i35_2_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i35_2_lut_LC_18_17_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i35_2_lut_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41203),
            .in3(N__49068),
            .lcout(\c0.n86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i167_LC_18_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i167_LC_18_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i167_LC_18_17_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i167_LC_18_17_2  (
            .in0(N__69002),
            .in1(N__71776),
            .in2(N__70125),
            .in3(N__67130),
            .lcout(\c0.data_in_frame_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71059),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i43_4_lut_LC_18_17_3 .C_ON=1'b0;
    defparam \c0.i43_4_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i43_4_lut_LC_18_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i43_4_lut_LC_18_17_3  (
            .in0(N__49069),
            .in1(N__43087),
            .in2(N__45051),
            .in3(N__44945),
            .lcout(\c0.n94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i143_LC_18_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i143_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i143_LC_18_17_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i143_LC_18_17_4  (
            .in0(N__63356),
            .in1(N__71775),
            .in2(N__69025),
            .in3(N__51200),
            .lcout(\c0.data_in_frame_17_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71059),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_938_LC_18_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_938_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_938_LC_18_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_938_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__47830),
            .in2(_gnd_net_),
            .in3(N__62981),
            .lcout(\c0.n19427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_944_LC_18_17_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_944_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_944_LC_18_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_944_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__65525),
            .in2(_gnd_net_),
            .in3(N__63774),
            .lcout(\c0.n19187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_231_LC_18_17_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_231_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_231_LC_18_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_231_LC_18_17_7  (
            .in0(N__48373),
            .in1(N__41260),
            .in2(N__41605),
            .in3(N__43278),
            .lcout(\c0.n19514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_356_LC_18_18_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_356_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_356_LC_18_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_356_LC_18_18_0  (
            .in0(N__67566),
            .in1(N__48595),
            .in2(N__47068),
            .in3(N__52491),
            .lcout(\c0.n29_adj_3148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_adj_905_LC_18_18_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_adj_905_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_adj_905_LC_18_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_2_lut_3_lut_adj_905_LC_18_18_1  (
            .in0(N__44716),
            .in1(N__65868),
            .in2(_gnd_net_),
            .in3(N__47772),
            .lcout(\c0.n17_adj_3451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i220_LC_18_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i220_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i220_LC_18_18_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i220_LC_18_18_2  (
            .in0(N__69216),
            .in1(N__66881),
            .in2(N__48617),
            .in3(N__64584),
            .lcout(\c0.data_in_frame_27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71085),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i215_LC_18_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i215_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i215_LC_18_18_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i215_LC_18_18_4  (
            .in0(N__62801),
            .in1(N__66880),
            .in2(N__69023),
            .in3(N__43668),
            .lcout(\c0.data_in_frame_26_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71085),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i211_LC_18_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i211_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i211_LC_18_18_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i211_LC_18_18_5  (
            .in0(N__66879),
            .in1(N__68553),
            .in2(N__58708),
            .in3(N__62802),
            .lcout(\c0.data_in_frame_26_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71085),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i151_LC_18_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i151_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i151_LC_18_18_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i151_LC_18_18_6  (
            .in0(N__68994),
            .in1(N__63939),
            .in2(_gnd_net_),
            .in3(N__41547),
            .lcout(data_in_frame_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71085),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_18_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_18_18_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_18_18_7  (
            .in0(N__41529),
            .in1(N__69215),
            .in2(N__56224),
            .in3(N__55467),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71085),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i152_LC_18_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i152_LC_18_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i152_LC_18_19_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i152_LC_18_19_1  (
            .in0(N__72260),
            .in1(N__63938),
            .in2(_gnd_net_),
            .in3(N__59116),
            .lcout(data_in_frame_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71098),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i134_LC_18_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i134_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i134_LC_18_19_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i134_LC_18_19_2  (
            .in0(N__65597),
            .in1(N__67939),
            .in2(_gnd_net_),
            .in3(N__45433),
            .lcout(data_in_frame_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71098),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_642_LC_18_19_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_642_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_642_LC_18_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_642_LC_18_19_3  (
            .in0(N__42003),
            .in1(N__66500),
            .in2(N__59794),
            .in3(N__66469),
            .lcout(\c0.n14_adj_3434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i43_4_lut_adj_515_LC_18_19_4 .C_ON=1'b0;
    defparam \c0.i43_4_lut_adj_515_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i43_4_lut_adj_515_LC_18_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i43_4_lut_adj_515_LC_18_19_4  (
            .in0(N__45052),
            .in1(N__49081),
            .in2(N__58552),
            .in3(N__44946),
            .lcout(\c0.n94_adj_3375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_327_LC_18_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_327_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_327_LC_18_19_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_327_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__60346),
            .in2(_gnd_net_),
            .in3(N__59459),
            .lcout(\c0.n19107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_855_LC_18_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_855_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_855_LC_18_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_855_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__41495),
            .in2(_gnd_net_),
            .in3(N__41433),
            .lcout(\c0.n18667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_2_lut_3_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \c0.i28_2_lut_3_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i28_2_lut_3_lut_LC_18_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i28_2_lut_3_lut_LC_18_20_0  (
            .in0(N__49079),
            .in1(N__43089),
            .in2(_gnd_net_),
            .in3(N__51808),
            .lcout(\c0.n61 ),
            .ltout(\c0.n61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_4_lut_adj_303_LC_18_20_1 .C_ON=1'b0;
    defparam \c0.i31_4_lut_adj_303_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i31_4_lut_adj_303_LC_18_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_4_lut_adj_303_LC_18_20_1  (
            .in0(N__41665),
            .in1(N__45211),
            .in2(N__41668),
            .in3(N__45345),
            .lcout(\c0.n64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_300_LC_18_20_2 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_300_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_300_LC_18_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i17_4_lut_adj_300_LC_18_20_2  (
            .in0(N__45189),
            .in1(N__41973),
            .in2(N__48778),
            .in3(N__42002),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i37_4_lut_LC_18_20_3 .C_ON=1'b0;
    defparam \c0.i37_4_lut_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i37_4_lut_LC_18_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i37_4_lut_LC_18_20_3  (
            .in0(N__48538),
            .in1(N__45346),
            .in2(N__45870),
            .in3(N__45190),
            .lcout(),
            .ltout(\c0.n86_adj_3393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i46_4_lut_adj_558_LC_18_20_4 .C_ON=1'b0;
    defparam \c0.i46_4_lut_adj_558_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i46_4_lut_adj_558_LC_18_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i46_4_lut_adj_558_LC_18_20_4  (
            .in0(N__43303),
            .in1(N__41659),
            .in2(N__41653),
            .in3(N__45306),
            .lcout(),
            .ltout(\c0.n95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_580_LC_18_20_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_580_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_580_LC_18_20_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i4_4_lut_adj_580_LC_18_20_5  (
            .in0(N__58159),
            .in1(N__43060),
            .in2(N__41650),
            .in3(N__43483),
            .lcout(\c0.n15_adj_3441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7__5174_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.data_in_2__7__5174_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7__5174_LC_18_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__7__5174_LC_18_21_0  (
            .in0(N__42574),
            .in1(N__41635),
            .in2(_gnd_net_),
            .in3(N__53179),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71127),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i135_LC_18_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i135_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i135_LC_18_21_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i135_LC_18_21_1  (
            .in0(N__41600),
            .in1(N__65590),
            .in2(_gnd_net_),
            .in3(N__69015),
            .lcout(data_in_frame_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71127),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i216_LC_18_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i216_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i216_LC_18_21_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i216_LC_18_21_2  (
            .in0(N__66896),
            .in1(N__62803),
            .in2(N__45868),
            .in3(N__72287),
            .lcout(\c0.data_in_frame_26_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71127),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_546_LC_18_21_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_546_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_546_LC_18_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_546_LC_18_21_4  (
            .in0(N__41577),
            .in1(N__70456),
            .in2(_gnd_net_),
            .in3(N__70180),
            .lcout(\c0.n20931 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i232_LC_18_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i232_LC_18_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i232_LC_18_21_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i232_LC_18_21_5  (
            .in0(N__72286),
            .in1(N__66897),
            .in2(N__52794),
            .in3(N__67166),
            .lcout(\c0.data_in_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71127),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i191_LC_18_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i191_LC_18_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i191_LC_18_21_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i191_LC_18_21_6  (
            .in0(N__69014),
            .in1(N__53714),
            .in2(_gnd_net_),
            .in3(N__66496),
            .lcout(data_in_frame_23_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71127),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_389_LC_18_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_389_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_389_LC_18_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_389_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__59332),
            .in2(_gnd_net_),
            .in3(N__59512),
            .lcout(\c0.n18537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_470_LC_18_22_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_470_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_470_LC_18_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_470_LC_18_22_0  (
            .in0(N__48829),
            .in1(N__52563),
            .in2(N__41694),
            .in3(N__41722),
            .lcout(\c0.n18_adj_3314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i233_LC_18_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i233_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i233_LC_18_22_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i233_LC_18_22_1  (
            .in0(N__41800),
            .in1(N__65260),
            .in2(N__66976),
            .in3(N__71869),
            .lcout(\c0.data_in_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71145),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i240_LC_18_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i240_LC_18_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i240_LC_18_22_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i240_LC_18_22_2  (
            .in0(N__71868),
            .in1(N__72285),
            .in2(N__41710),
            .in3(N__66947),
            .lcout(\c0.data_in_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71145),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i239_LC_18_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i239_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i239_LC_18_22_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i239_LC_18_22_3  (
            .in0(N__66943),
            .in1(N__69022),
            .in2(N__41695),
            .in3(N__71870),
            .lcout(\c0.data_in_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71145),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_357_LC_18_22_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_357_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_357_LC_18_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_357_LC_18_22_4  (
            .in0(N__53263),
            .in1(N__53512),
            .in2(N__43687),
            .in3(N__46095),
            .lcout(),
            .ltout(\c0.n10_adj_3152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_768_LC_18_22_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_768_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_768_LC_18_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_768_LC_18_22_5  (
            .in0(N__43389),
            .in1(N__49507),
            .in2(N__41677),
            .in3(N__49459),
            .lcout(\c0.n21117 ),
            .ltout(\c0.n21117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_446_LC_18_22_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_446_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_446_LC_18_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_446_LC_18_22_6  (
            .in0(N__41782),
            .in1(N__41799),
            .in2(N__41791),
            .in3(N__43522),
            .lcout(\c0.n40_adj_3282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_351_LC_18_23_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_351_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_351_LC_18_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i10_4_lut_adj_351_LC_18_23_0  (
            .in0(N__41788),
            .in1(N__52423),
            .in2(N__49522),
            .in3(N__45937),
            .lcout(\c0.n5_adj_3142 ),
            .ltout(\c0.n5_adj_3142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_462_LC_18_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_462_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_462_LC_18_23_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_462_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41776),
            .in3(N__46003),
            .lcout(),
            .ltout(\c0.n22_adj_3305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_467_LC_18_23_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_467_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_467_LC_18_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_467_LC_18_23_2  (
            .in0(N__59595),
            .in1(N__49346),
            .in2(N__41773),
            .in3(N__49375),
            .lcout(),
            .ltout(\c0.n37_adj_3309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_479_LC_18_23_3 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_479_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_479_LC_18_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_479_LC_18_23_3  (
            .in0(N__46066),
            .in1(N__53560),
            .in2(N__41770),
            .in3(N__43528),
            .lcout(),
            .ltout(\c0.n21099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_492_LC_18_23_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_492_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_492_LC_18_23_4 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i2_4_lut_adj_492_LC_18_23_4  (
            .in0(N__52519),
            .in1(N__48736),
            .in2(N__41767),
            .in3(N__41764),
            .lcout(),
            .ltout(\c0.n10_adj_3353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_542_LC_18_23_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_542_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_542_LC_18_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_542_LC_18_23_5  (
            .in0(N__41740),
            .in1(N__43561),
            .in2(N__41758),
            .in3(N__43702),
            .lcout(\c0.n21111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_490_LC_18_24_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_490_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_490_LC_18_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_490_LC_18_24_0  (
            .in0(N__41971),
            .in1(N__41998),
            .in2(_gnd_net_),
            .in3(N__49543),
            .lcout(),
            .ltout(\c0.n9_adj_3352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_491_LC_18_24_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_491_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_491_LC_18_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_491_LC_18_24_1  (
            .in0(N__59700),
            .in1(N__43555),
            .in2(N__41743),
            .in3(N__45889),
            .lcout(\c0.n21051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i224_LC_18_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i224_LC_18_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i224_LC_18_24_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i224_LC_18_24_3  (
            .in0(N__72241),
            .in1(N__64565),
            .in2(N__42004),
            .in3(N__66912),
            .lcout(\c0.data_in_frame_27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71170),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i223_LC_18_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i223_LC_18_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i223_LC_18_24_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i223_LC_18_24_4  (
            .in0(N__41972),
            .in1(N__69031),
            .in2(N__64578),
            .in3(N__66916),
            .lcout(\c0.data_in_frame_27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71170),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i217_LC_18_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i217_LC_18_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i217_LC_18_24_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i217_LC_18_24_5  (
            .in0(N__65242),
            .in1(N__64564),
            .in2(N__66958),
            .in3(N__43385),
            .lcout(\c0.data_in_frame_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71170),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_454_LC_18_24_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_454_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_454_LC_18_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_454_LC_18_24_6  (
            .in0(N__70382),
            .in1(N__70337),
            .in2(N__41950),
            .in3(N__51862),
            .lcout(\c0.n21003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i138_LC_18_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i138_LC_18_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i138_LC_18_24_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i138_LC_18_24_7  (
            .in0(N__71734),
            .in1(N__63377),
            .in2(N__52331),
            .in3(N__71506),
            .lcout(\c0.data_in_frame_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71170),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_405_LC_18_25_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_405_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_405_LC_18_25_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i5_3_lut_adj_405_LC_18_25_0  (
            .in0(N__41851),
            .in1(N__41926),
            .in2(_gnd_net_),
            .in3(N__41908),
            .lcout(\c0.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7__5182_LC_18_25_1 .C_ON=1'b0;
    defparam \c0.data_in_1__7__5182_LC_18_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7__5182_LC_18_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__7__5182_LC_18_25_1  (
            .in0(N__53209),
            .in1(N__42577),
            .in2(_gnd_net_),
            .in3(N__43941),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71180),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5__5184_LC_18_25_2 .C_ON=1'b0;
    defparam \c0.data_in_1__5__5184_LC_18_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5__5184_LC_18_25_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_1__5__5184_LC_18_25_2  (
            .in0(N__41852),
            .in1(N__53211),
            .in2(_gnd_net_),
            .in3(N__41884),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71180),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_902_LC_18_25_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_902_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_902_LC_18_25_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_902_LC_18_25_4  (
            .in0(N__66924),
            .in1(N__41833),
            .in2(N__55886),
            .in3(N__42071),
            .lcout(n20896),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__0__5189_LC_18_25_5 .C_ON=1'b0;
    defparam \c0.data_in_1__0__5189_LC_18_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0__5189_LC_18_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__0__5189_LC_18_25_5  (
            .in0(N__53208),
            .in1(N__42640),
            .in2(_gnd_net_),
            .in3(N__42606),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71180),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__0__5197_LC_18_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0__0__5197_LC_18_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0__5197_LC_18_25_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__0__5197_LC_18_25_6  (
            .in0(N__42607),
            .in1(N__53210),
            .in2(_gnd_net_),
            .in3(N__43954),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71180),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i187_LC_18_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i187_LC_18_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i187_LC_18_25_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i187_LC_18_25_7  (
            .in0(N__68645),
            .in1(N__53693),
            .in2(_gnd_net_),
            .in3(N__43410),
            .lcout(data_in_frame_23_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71180),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_752_LC_18_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_752_LC_18_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_752_LC_18_26_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_752_LC_18_26_0  (
            .in0(N__43924),
            .in1(N__43973),
            .in2(N__52921),
            .in3(N__42576),
            .lcout(\c0.n12_adj_3230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_402_LC_18_26_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_402_LC_18_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_402_LC_18_26_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i5_3_lut_adj_402_LC_18_26_1  (
            .in0(N__43972),
            .in1(N__42575),
            .in2(_gnd_net_),
            .in3(N__43923),
            .lcout(\c0.n11443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i194_LC_18_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i194_LC_18_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i194_LC_18_26_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i194_LC_18_26_4  (
            .in0(N__46134),
            .in1(N__71536),
            .in2(_gnd_net_),
            .in3(N__70374),
            .lcout(data_in_frame_24_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71191),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1__5196_LC_18_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0__1__5196_LC_18_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1__5196_LC_18_26_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__1__5196_LC_18_26_7  (
            .in0(N__53225),
            .in1(N__42540),
            .in2(_gnd_net_),
            .in3(N__43888),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71191),
            .ce(),
            .sr(_gnd_net_));
    defparam i16083_1_lut_2_lut_3_lut_LC_18_27_5.C_ON=1'b0;
    defparam i16083_1_lut_2_lut_3_lut_LC_18_27_5.SEQ_MODE=4'b0000;
    defparam i16083_1_lut_2_lut_3_lut_LC_18_27_5.LUT_INIT=16'b0011001110111011;
    LogicCell40 i16083_1_lut_2_lut_3_lut_LC_18_27_5 (
            .in0(N__42517),
            .in1(N__42370),
            .in2(_gnd_net_),
            .in3(N__42331),
            .lcout(n1295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i12201_2_lut_LC_19_7_0 .C_ON=1'b0;
    defparam \c0.rx.i12201_2_lut_LC_19_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i12201_2_lut_LC_19_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i12201_2_lut_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(N__43859),
            .in2(_gnd_net_),
            .in3(N__43817),
            .lcout(n15645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_566_LC_19_7_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_566_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_566_LC_19_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_566_LC_19_7_1  (
            .in0(N__51410),
            .in1(N__51331),
            .in2(_gnd_net_),
            .in3(N__51283),
            .lcout(\c0.n11549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_322_LC_19_7_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_322_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_322_LC_19_7_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_322_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(N__61874),
            .in2(_gnd_net_),
            .in3(N__47255),
            .lcout(\c0.n5_adj_3099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_19_7_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_19_7_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_19_7_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i60_LC_19_7_3  (
            .in0(N__69436),
            .in1(N__64345),
            .in2(N__47269),
            .in3(N__61685),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71214),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_19_7_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_19_7_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_19_7_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_19_7_4  (
            .in0(N__71374),
            .in1(N__61684),
            .in2(N__62002),
            .in3(N__49906),
            .lcout(\c0.data_in_frame_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71214),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_19_7_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_19_7_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_19_7_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i58_LC_19_7_5  (
            .in0(N__61683),
            .in1(N__64344),
            .in2(N__63149),
            .in3(N__71375),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71214),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_3_lut_LC_19_7_6 .C_ON=1'b0;
    defparam \c0.i13_3_lut_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_3_lut_LC_19_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i13_3_lut_LC_19_7_6  (
            .in0(N__63135),
            .in1(N__42691),
            .in2(_gnd_net_),
            .in3(N__63180),
            .lcout(\c0.n31_adj_3121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_276_LC_19_7_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_276_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_276_LC_19_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_276_LC_19_7_7  (
            .in0(N__63181),
            .in1(N__42673),
            .in2(N__63148),
            .in3(N__56642),
            .lcout(\c0.n25_adj_3045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_19_8_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_19_8_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_19_8_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i18_LC_19_8_0  (
            .in0(N__44215),
            .in1(N__61759),
            .in2(N__54627),
            .in3(N__71348),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71202),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_302_LC_19_8_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_302_LC_19_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_302_LC_19_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_302_LC_19_8_1  (
            .in0(N__44028),
            .in1(N__46390),
            .in2(N__47153),
            .in3(N__51255),
            .lcout(),
            .ltout(\c0.n14_adj_3073_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_595_LC_19_8_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_595_LC_19_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_595_LC_19_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_595_LC_19_8_2  (
            .in0(N__46414),
            .in1(N__42724),
            .in2(N__42643),
            .in3(N__42783),
            .lcout(\c0.n4_adj_3009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_LC_19_8_3 .C_ON=1'b0;
    defparam \c0.i9_2_lut_LC_19_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_LC_19_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i9_2_lut_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__51330),
            .in2(_gnd_net_),
            .in3(N__51257),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_294_LC_19_8_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_294_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_294_LC_19_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_294_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(N__55213),
            .in2(_gnd_net_),
            .in3(N__54242),
            .lcout(\c0.n10_adj_3068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_19_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_19_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_19_8_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i24_LC_19_8_5  (
            .in0(N__61758),
            .in1(N__44216),
            .in2(N__72270),
            .in3(N__44157),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71202),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i34_LC_19_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i34_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i34_LC_19_8_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i34_LC_19_8_6  (
            .in0(N__44119),
            .in1(N__61760),
            .in2(N__55234),
            .in3(N__71349),
            .lcout(\c0.data_in_frame_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71202),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_4_lut_LC_19_8_7 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_4_lut_LC_19_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_4_lut_LC_19_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_2_lut_3_lut_4_lut_LC_19_8_7  (
            .in0(N__44029),
            .in1(N__51256),
            .in2(N__50680),
            .in3(N__55180),
            .lcout(\c0.n22_adj_3041 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_476_LC_19_9_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_476_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_476_LC_19_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_476_LC_19_9_0  (
            .in0(N__54297),
            .in1(N__44156),
            .in2(N__46345),
            .in3(N__42784),
            .lcout(\c0.n21079 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i67_LC_19_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i67_LC_19_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i67_LC_19_9_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i67_LC_19_9_1  (
            .in0(N__55795),
            .in1(N__64198),
            .in2(N__50149),
            .in3(N__68648),
            .lcout(\c0.data_in_frame_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71193),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_19_9_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_19_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_2_lut_3_lut_4_lut_LC_19_9_2  (
            .in0(N__50407),
            .in1(N__44155),
            .in2(N__50359),
            .in3(N__50592),
            .lcout(\c0.n13_adj_3017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_730_LC_19_9_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_730_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_730_LC_19_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_730_LC_19_9_3  (
            .in0(N__44382),
            .in1(N__54296),
            .in2(N__47152),
            .in3(N__61073),
            .lcout(\c0.n13_adj_3504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_726_LC_19_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_726_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_726_LC_19_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_726_LC_19_9_4  (
            .in0(_gnd_net_),
            .in1(N__47715),
            .in2(_gnd_net_),
            .in3(N__49851),
            .lcout(\c0.n6_adj_3501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_19_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_19_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_19_9_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i4_LC_19_9_5  (
            .in0(N__61686),
            .in1(N__69435),
            .in2(N__55819),
            .in3(N__62129),
            .lcout(data_in_frame_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71193),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_19_9_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_19_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_19_9_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i3_LC_19_9_6  (
            .in0(N__68647),
            .in1(N__55796),
            .in2(N__61099),
            .in3(N__61687),
            .lcout(data_in_frame_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71193),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_282_LC_19_9_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_282_LC_19_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_282_LC_19_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_282_LC_19_9_7  (
            .in0(N__44383),
            .in1(N__62128),
            .in2(_gnd_net_),
            .in3(N__54427),
            .lcout(\c0.n11516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_663_LC_19_10_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_663_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_663_LC_19_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_663_LC_19_10_0  (
            .in0(N__50347),
            .in1(N__54422),
            .in2(N__50599),
            .in3(N__55181),
            .lcout(\c0.n14_adj_3480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_844_LC_19_10_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_844_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_844_LC_19_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_844_LC_19_10_1  (
            .in0(N__61080),
            .in1(N__56810),
            .in2(N__46292),
            .in3(N__62163),
            .lcout(\c0.n13_adj_3546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_702_LC_19_10_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_702_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_702_LC_19_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i5_4_lut_adj_702_LC_19_10_2  (
            .in0(N__62164),
            .in1(N__55182),
            .in2(N__50600),
            .in3(N__46273),
            .lcout(),
            .ltout(\c0.n13_adj_3490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12053_4_lut_LC_19_10_3 .C_ON=1'b0;
    defparam \c0.i12053_4_lut_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12053_4_lut_LC_19_10_3 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \c0.i12053_4_lut_LC_19_10_3  (
            .in0(N__42733),
            .in1(N__42772),
            .in2(N__42766),
            .in3(N__42763),
            .lcout(\c0.n15497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_608_LC_19_10_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_608_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_608_LC_19_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_608_LC_19_10_4  (
            .in0(N__50346),
            .in1(N__54421),
            .in2(N__56830),
            .in3(N__61079),
            .lcout(\c0.n14_adj_3459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_19_10_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_19_10_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_19_10_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i1_LC_19_10_5  (
            .in0(N__55800),
            .in1(N__65240),
            .in2(N__46293),
            .in3(N__61730),
            .lcout(data_in_frame_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71182),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_524_LC_19_10_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_524_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_524_LC_19_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_524_LC_19_10_6  (
            .in0(N__54298),
            .in1(N__61078),
            .in2(N__56829),
            .in3(N__55364),
            .lcout(\c0.n11_adj_3394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_635_LC_19_10_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_635_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_635_LC_19_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_635_LC_19_10_7  (
            .in0(N__56032),
            .in1(N__45093),
            .in2(N__42844),
            .in3(N__47270),
            .lcout(\c0.n10_adj_3207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_743_LC_19_11_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_743_LC_19_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_743_LC_19_11_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i6_2_lut_adj_743_LC_19_11_0  (
            .in0(N__44355),
            .in1(_gnd_net_),
            .in2(N__42796),
            .in3(_gnd_net_),
            .lcout(\c0.n39_adj_3398 ),
            .ltout(\c0.n39_adj_3398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_761_LC_19_11_1 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_761_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_761_LC_19_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_761_LC_19_11_1  (
            .in0(N__44292),
            .in1(N__44280),
            .in2(N__42826),
            .in3(N__50553),
            .lcout(\c0.n28_adj_3519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_795_LC_19_11_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_795_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_795_LC_19_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_adj_795_LC_19_11_2  (
            .in0(N__50551),
            .in1(N__56800),
            .in2(_gnd_net_),
            .in3(N__50317),
            .lcout(\c0.n13_adj_3526 ),
            .ltout(\c0.n13_adj_3526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_830_LC_19_11_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_830_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_830_LC_19_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_830_LC_19_11_3  (
            .in0(N__42816),
            .in1(N__42805),
            .in2(N__42799),
            .in3(N__42874),
            .lcout(\c0.n13_adj_3513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_19_11_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_19_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_19_11_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i45_LC_19_11_4  (
            .in0(N__61726),
            .in1(N__60336),
            .in2(N__50023),
            .in3(N__72611),
            .lcout(\c0.data_in_frame_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71171),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_790_LC_19_11_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_790_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_790_LC_19_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_790_LC_19_11_5  (
            .in0(_gnd_net_),
            .in1(N__42792),
            .in2(_gnd_net_),
            .in3(N__50552),
            .lcout(\c0.n24_adj_3011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_19_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_19_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_19_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i21_LC_19_11_6  (
            .in0(N__61725),
            .in1(N__44240),
            .in2(N__60983),
            .in3(N__72610),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71171),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_adj_727_LC_19_11_7 .C_ON=1'b0;
    defparam \c0.i27_4_lut_adj_727_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_adj_727_LC_19_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_adj_727_LC_19_11_7  (
            .in0(N__44293),
            .in1(N__44281),
            .in2(N__47278),
            .in3(N__44272),
            .lcout(\c0.n60_adj_3503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_552_LC_19_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_552_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_552_LC_19_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_552_LC_19_12_0  (
            .in0(N__55588),
            .in1(N__56299),
            .in2(_gnd_net_),
            .in3(N__55378),
            .lcout(),
            .ltout(\c0.n16_adj_3416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_762_LC_19_12_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_762_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_762_LC_19_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_762_LC_19_12_1  (
            .in0(N__42883),
            .in1(N__61225),
            .in2(N__42877),
            .in3(N__50691),
            .lcout(\c0.n20088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_826_LC_19_12_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_826_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_826_LC_19_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_826_LC_19_12_2  (
            .in0(N__42861),
            .in1(N__47217),
            .in2(N__47559),
            .in3(N__54623),
            .lcout(\c0.n16_adj_3542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_799_LC_19_12_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_799_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_799_LC_19_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_799_LC_19_12_3  (
            .in0(_gnd_net_),
            .in1(N__61092),
            .in2(_gnd_net_),
            .in3(N__54384),
            .lcout(\c0.n5_adj_3528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_2_lut_3_lut_LC_19_12_4 .C_ON=1'b0;
    defparam \c0.i26_2_lut_3_lut_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i26_2_lut_3_lut_LC_19_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i26_2_lut_3_lut_LC_19_12_4  (
            .in0(N__50639),
            .in1(N__44158),
            .in2(_gnd_net_),
            .in3(N__50566),
            .lcout(\c0.n78 ),
            .ltout(\c0.n78_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_567_LC_19_12_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_567_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_567_LC_19_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_567_LC_19_12_5  (
            .in0(N__55509),
            .in1(N__50239),
            .in2(N__42850),
            .in3(N__54130),
            .lcout(\c0.n11800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_496_LC_19_12_6 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_496_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_496_LC_19_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_496_LC_19_12_6  (
            .in0(N__50640),
            .in1(N__55585),
            .in2(_gnd_net_),
            .in3(N__47391),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_19_13_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_19_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_19_13_0  (
            .in0(N__62256),
            .in1(N__63105),
            .in2(N__44634),
            .in3(N__56911),
            .lcout(),
            .ltout(\c0.n30_adj_3119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_334_LC_19_13_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_334_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_334_LC_19_13_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_334_LC_19_13_1  (
            .in0(N__56719),
            .in1(N__50108),
            .in2(N__42847),
            .in3(N__57142),
            .lcout(\c0.n33_adj_3122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_801_LC_19_13_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_801_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_801_LC_19_13_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_801_LC_19_13_2  (
            .in0(N__49879),
            .in1(N__62682),
            .in2(N__42968),
            .in3(N__57307),
            .lcout(\c0.n20055 ),
            .ltout(\c0.n20055_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_329_LC_19_13_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_329_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_329_LC_19_13_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i13_4_lut_adj_329_LC_19_13_3  (
            .in0(N__63843),
            .in1(N__62411),
            .in2(N__42943),
            .in3(N__42926),
            .lcout(),
            .ltout(\c0.n37_adj_3110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_19_13_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_19_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_LC_19_13_4  (
            .in0(N__63155),
            .in1(N__42900),
            .in2(N__42904),
            .in3(N__56646),
            .lcout(\c0.n43_adj_3116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_807_LC_19_13_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_807_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_807_LC_19_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_807_LC_19_13_5  (
            .in0(N__63202),
            .in1(_gnd_net_),
            .in2(N__63070),
            .in3(N__63231),
            .lcout(\c0.n22_adj_3115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i83_LC_19_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i83_LC_19_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i83_LC_19_14_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i83_LC_19_14_0  (
            .in0(N__68593),
            .in1(N__66012),
            .in2(N__43042),
            .in3(N__62793),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71128),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_813_LC_19_14_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_813_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_813_LC_19_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_813_LC_19_14_1  (
            .in0(N__44499),
            .in1(N__62587),
            .in2(N__45022),
            .in3(N__57330),
            .lcout(\c0.n23_adj_3534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i84_LC_19_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i84_LC_19_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i84_LC_19_14_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i84_LC_19_14_2  (
            .in0(N__66011),
            .in1(N__62794),
            .in2(N__44481),
            .in3(N__69408),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71128),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_886_LC_19_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_886_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_886_LC_19_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_886_LC_19_14_3  (
            .in0(N__62465),
            .in1(N__43034),
            .in2(_gnd_net_),
            .in3(N__44538),
            .lcout(),
            .ltout(\c0.n6_adj_3024_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_245_LC_19_14_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_245_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_245_LC_19_14_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_245_LC_19_14_4  (
            .in0(N__56352),
            .in1(N__57328),
            .in2(N__42889),
            .in3(N__62683),
            .lcout(\c0.n18435 ),
            .ltout(\c0.n18435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_LC_19_14_5 .C_ON=1'b0;
    defparam \c0.i8_2_lut_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_LC_19_14_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i8_2_lut_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42886),
            .in3(N__47684),
            .lcout(\c0.n25_adj_3035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_887_LC_19_14_6 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_887_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_887_LC_19_14_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_887_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(N__57329),
            .in2(N__43041),
            .in3(N__62466),
            .lcout(\c0.n14_adj_3007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_929_LC_19_14_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_929_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_929_LC_19_14_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_929_LC_19_14_7  (
            .in0(N__65864),
            .in1(N__52093),
            .in2(N__55671),
            .in3(N__43273),
            .lcout(\c0.n17871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_19_15_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_19_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_19_15_0  (
            .in0(N__57075),
            .in1(N__62467),
            .in2(N__44482),
            .in3(N__62911),
            .lcout(),
            .ltout(\c0.n28_adj_3120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_335_LC_19_15_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_335_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_335_LC_19_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_335_LC_19_15_1  (
            .in0(N__43012),
            .in1(N__43000),
            .in2(N__42991),
            .in3(N__42988),
            .lcout(\c0.n20052 ),
            .ltout(\c0.n20052_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_342_LC_19_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_342_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_342_LC_19_15_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_342_LC_19_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42979),
            .in3(N__44804),
            .lcout(),
            .ltout(\c0.n10_adj_3129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_345_LC_19_15_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_345_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_345_LC_19_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_345_LC_19_15_3  (
            .in0(N__51617),
            .in1(N__48068),
            .in2(N__42976),
            .in3(N__51991),
            .lcout(),
            .ltout(\c0.n18400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_349_LC_19_15_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_349_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_349_LC_19_15_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_349_LC_19_15_4  (
            .in0(N__45565),
            .in1(N__61878),
            .in2(N__42973),
            .in3(N__57646),
            .lcout(\c0.n13_adj_3139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_LC_19_15_5 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_LC_19_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_LC_19_15_5  (
            .in0(N__55516),
            .in1(N__57371),
            .in2(N__51846),
            .in3(N__54136),
            .lcout(\c0.n37_adj_3215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_4_lut_LC_19_16_1 .C_ON=1'b0;
    defparam \c0.i12_3_lut_4_lut_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_4_lut_LC_19_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_3_lut_4_lut_LC_19_16_1  (
            .in0(N__55921),
            .in1(N__51108),
            .in2(N__51847),
            .in3(N__50678),
            .lcout(),
            .ltout(\c0.n35_adj_3342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_942_LC_19_16_2 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_942_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_942_LC_19_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_adj_942_LC_19_16_2  (
            .in0(N__43237),
            .in1(N__43213),
            .in2(N__43198),
            .in3(N__50082),
            .lcout(),
            .ltout(\c0.n44_adj_3561_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_943_LC_19_16_3 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_943_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_943_LC_19_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_adj_943_LC_19_16_3  (
            .in0(N__43195),
            .in1(N__43180),
            .in2(N__43156),
            .in3(N__43153),
            .lcout(\c0.n21118 ),
            .ltout(\c0.n21118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_638_LC_19_16_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_638_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_638_LC_19_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_638_LC_19_16_4  (
            .in0(N__43120),
            .in1(N__57454),
            .in2(N__43102),
            .in3(N__45182),
            .lcout(\c0.n11_adj_3206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_352_LC_19_16_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_352_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_352_LC_19_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_352_LC_19_16_5  (
            .in0(N__57572),
            .in1(N__48489),
            .in2(N__48032),
            .in3(N__43099),
            .lcout(\c0.n20826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i45_4_lut_adj_556_LC_19_17_0 .C_ON=1'b0;
    defparam \c0.i45_4_lut_adj_556_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i45_4_lut_adj_556_LC_19_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i45_4_lut_adj_556_LC_19_17_0  (
            .in0(N__45339),
            .in1(N__43048),
            .in2(N__66532),
            .in3(N__45316),
            .lcout(),
            .ltout(\c0.n96_adj_3418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_adj_562_LC_19_17_1 .C_ON=1'b0;
    defparam \c0.i48_4_lut_adj_562_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_adj_562_LC_19_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i48_4_lut_adj_562_LC_19_17_1  (
            .in0(N__58009),
            .in1(N__43088),
            .in2(N__43063),
            .in3(N__57532),
            .lcout(\c0.n99_adj_3424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_3_lut_LC_19_17_2 .C_ON=1'b0;
    defparam \c0.i26_3_lut_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i26_3_lut_LC_19_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i26_3_lut_LC_19_17_2  (
            .in0(N__70390),
            .in1(N__70264),
            .in2(_gnd_net_),
            .in3(N__45188),
            .lcout(\c0.n77_adj_3415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_646_LC_19_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_646_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_646_LC_19_17_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_646_LC_19_17_3  (
            .in0(N__64003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58053),
            .lcout(\c0.n10_adj_3474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_867_LC_19_17_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_867_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_867_LC_19_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_867_LC_19_17_4  (
            .in0(N__51133),
            .in1(N__48260),
            .in2(N__51718),
            .in3(N__51674),
            .lcout(\c0.n20801 ),
            .ltout(\c0.n20801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i45_4_lut_LC_19_17_5 .C_ON=1'b0;
    defparam \c0.i45_4_lut_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i45_4_lut_LC_19_17_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i45_4_lut_LC_19_17_5  (
            .in0(N__43554),
            .in1(N__59809),
            .in2(N__43321),
            .in3(N__45338),
            .lcout(),
            .ltout(\c0.n96_adj_3401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_adj_538_LC_19_17_6 .C_ON=1'b0;
    defparam \c0.i48_4_lut_adj_538_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_adj_538_LC_19_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i48_4_lut_adj_538_LC_19_17_6  (
            .in0(N__43299),
            .in1(N__51807),
            .in2(N__43318),
            .in3(N__45315),
            .lcout(\c0.n99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i204_LC_19_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i204_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i204_LC_19_18_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i204_LC_19_18_0  (
            .in0(N__66923),
            .in1(N__63394),
            .in2(N__49213),
            .in3(N__69218),
            .lcout(\c0.data_in_frame_25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71099),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i148_LC_19_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i148_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i148_LC_19_18_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i148_LC_19_18_1  (
            .in0(N__69217),
            .in1(N__63943),
            .in2(_gnd_net_),
            .in3(N__64002),
            .lcout(data_in_frame_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71099),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_adj_641_LC_19_18_3 .C_ON=1'b0;
    defparam \c0.i14_2_lut_adj_641_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_adj_641_LC_19_18_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i14_2_lut_adj_641_LC_19_18_3  (
            .in0(_gnd_net_),
            .in1(N__67666),
            .in2(_gnd_net_),
            .in3(N__58037),
            .lcout(\c0.n47_adj_3408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_3_lut_LC_19_18_4 .C_ON=1'b0;
    defparam \c0.i28_3_lut_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i28_3_lut_LC_19_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i28_3_lut_LC_19_18_4  (
            .in0(N__48177),
            .in1(N__44944),
            .in2(_gnd_net_),
            .in3(N__48860),
            .lcout(\c0.n61_adj_3387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_2_lut_3_lut_LC_19_18_5 .C_ON=1'b0;
    defparam \c0.i10_2_lut_3_lut_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_2_lut_3_lut_LC_19_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i10_2_lut_3_lut_LC_19_18_5  (
            .in0(N__55670),
            .in1(N__52103),
            .in2(_gnd_net_),
            .in3(N__43282),
            .lcout(\c0.n43_adj_3386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_adj_734_LC_19_18_6 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_adj_734_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_adj_734_LC_19_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i9_2_lut_3_lut_adj_734_LC_19_18_6  (
            .in0(N__57723),
            .in1(N__48133),
            .in2(_gnd_net_),
            .in3(N__48654),
            .lcout(\c0.n42_adj_3064 ),
            .ltout(\c0.n42_adj_3064_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_3_lut_LC_19_18_7 .C_ON=1'b0;
    defparam \c0.i27_3_lut_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i27_3_lut_LC_19_18_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i27_3_lut_LC_19_18_7  (
            .in0(N__48103),
            .in1(N__45038),
            .in2(N__43240),
            .in3(_gnd_net_),
            .lcout(\c0.n60_adj_3065 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i178_LC_19_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i178_LC_19_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i178_LC_19_19_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i178_LC_19_19_0  (
            .in0(N__71464),
            .in1(N__67522),
            .in2(_gnd_net_),
            .in3(N__70438),
            .lcout(data_in_frame_22_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71114),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i98_LC_19_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i98_LC_19_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i98_LC_19_19_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i98_LC_19_19_1  (
            .in0(N__66209),
            .in1(N__67187),
            .in2(N__63853),
            .in3(N__71466),
            .lcout(\c0.data_in_frame_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71114),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12045_2_lut_3_lut_LC_19_19_2 .C_ON=1'b0;
    defparam \c0.i12045_2_lut_3_lut_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12045_2_lut_3_lut_LC_19_19_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i12045_2_lut_3_lut_LC_19_19_2  (
            .in0(N__60274),
            .in1(N__60000),
            .in2(_gnd_net_),
            .in3(N__60132),
            .lcout(\c0.n15489 ),
            .ltout(\c0.n15489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i123_LC_19_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i123_LC_19_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i123_LC_19_19_3 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \c0.data_in_frame_0__i123_LC_19_19_3  (
            .in0(N__68691),
            .in1(N__43333),
            .in2(N__43336),
            .in3(N__64221),
            .lcout(\c0.data_in_frame_15_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71114),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_234_LC_19_19_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_234_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_234_LC_19_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_234_LC_19_19_4  (
            .in0(N__45564),
            .in1(N__43332),
            .in2(_gnd_net_),
            .in3(N__48325),
            .lcout(\c0.n19505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i106_LC_19_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i106_LC_19_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i106_LC_19_19_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i106_LC_19_19_6  (
            .in0(N__71465),
            .in1(N__48326),
            .in2(N__71898),
            .in3(N__66210),
            .lcout(\c0.data_in_frame_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71114),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i144_LC_19_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i144_LC_19_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i144_LC_19_19_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i144_LC_19_19_7  (
            .in0(N__71766),
            .in1(N__63413),
            .in2(N__56524),
            .in3(N__72261),
            .lcout(\c0.data_in_frame_17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71114),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_559_LC_19_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_559_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_559_LC_19_20_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_559_LC_19_20_0  (
            .in0(N__65694),
            .in1(N__65797),
            .in2(_gnd_net_),
            .in3(N__53869),
            .lcout(\c0.n12035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i181_LC_19_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i181_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i181_LC_19_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i181_LC_19_20_1  (
            .in0(N__53326),
            .in1(N__72748),
            .in2(_gnd_net_),
            .in3(N__67504),
            .lcout(data_in_frame_22_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71129),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_716_LC_19_20_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_716_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_716_LC_19_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_716_LC_19_20_2  (
            .in0(N__70428),
            .in1(N__45509),
            .in2(N__43420),
            .in3(N__53325),
            .lcout(\c0.n12_adj_3494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__7__5383_LC_19_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__7__5383_LC_19_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__7__5383_LC_19_20_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame_6__7__5383_LC_19_20_3  (
            .in0(N__46886),
            .in1(_gnd_net_),
            .in2(N__43465),
            .in3(N__43434),
            .lcout(data_out_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71129),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i188_LC_19_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i188_LC_19_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i188_LC_19_20_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i188_LC_19_20_4  (
            .in0(N__69247),
            .in1(N__53720),
            .in2(_gnd_net_),
            .in3(N__45510),
            .lcout(data_in_frame_23_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71129),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_534_LC_19_20_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_534_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_534_LC_19_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_534_LC_19_20_6  (
            .in0(N__43419),
            .in1(N__70123),
            .in2(N__71284),
            .in3(N__53868),
            .lcout(),
            .ltout(\c0.n13_adj_3405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_535_LC_19_20_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_535_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_535_LC_19_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_535_LC_19_20_7  (
            .in0(N__50908),
            .in1(N__45490),
            .in2(N__43396),
            .in3(N__47980),
            .lcout(\c0.n24_adj_3134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_adj_497_LC_19_21_0 .C_ON=1'b0;
    defparam \c0.i29_4_lut_adj_497_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_adj_497_LC_19_21_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i29_4_lut_adj_497_LC_19_21_0  (
            .in0(N__53333),
            .in1(N__43641),
            .in2(N__43393),
            .in3(N__45929),
            .lcout(\c0.n78_adj_3357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_547_LC_19_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_547_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_547_LC_19_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_547_LC_19_21_1  (
            .in0(N__65695),
            .in1(N__65782),
            .in2(N__69607),
            .in3(N__53870),
            .lcout(\c0.n17880 ),
            .ltout(\c0.n17880_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_531_LC_19_21_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_531_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_531_LC_19_21_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_531_LC_19_21_2  (
            .in0(N__53755),
            .in1(N__69903),
            .in2(N__43363),
            .in3(N__52130),
            .lcout(\c0.n19342 ),
            .ltout(\c0.n19342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_539_LC_19_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_539_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_539_LC_19_21_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_539_LC_19_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43360),
            .in3(N__59738),
            .lcout(\c0.n19496 ),
            .ltout(\c0.n19496_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_527_LC_19_21_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_527_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_527_LC_19_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_527_LC_19_21_4  (
            .in0(N__69517),
            .in1(N__43357),
            .in2(N__43351),
            .in3(N__45930),
            .lcout(\c0.n15_adj_3395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_3_lut_4_lut_adj_627_LC_19_21_5 .C_ON=1'b0;
    defparam \c0.i12_3_lut_4_lut_adj_627_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_3_lut_4_lut_adj_627_LC_19_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_3_lut_4_lut_adj_627_LC_19_21_5  (
            .in0(N__59742),
            .in1(N__43547),
            .in2(N__59692),
            .in3(N__48894),
            .lcout(\c0.n32_adj_3095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_778_LC_19_21_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_778_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_778_LC_19_21_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_4_lut_adj_778_LC_19_21_6  (
            .in0(N__66382),
            .in1(N__66465),
            .in2(N__58760),
            .in3(N__45825),
            .lcout(\c0.n25_adj_3524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_465_LC_19_22_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_465_LC_19_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_465_LC_19_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_465_LC_19_22_0  (
            .in0(N__58726),
            .in1(N__45745),
            .in2(N__49183),
            .in3(N__43695),
            .lcout(),
            .ltout(\c0.n36_adj_3307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_468_LC_19_22_1 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_468_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_468_LC_19_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i18_4_lut_adj_468_LC_19_22_1  (
            .in0(N__43520),
            .in1(N__52671),
            .in2(N__43531),
            .in3(N__49302),
            .lcout(\c0.n39_adj_3312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_adj_500_LC_19_22_2 .C_ON=1'b0;
    defparam \c0.i26_4_lut_adj_500_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_adj_500_LC_19_22_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i26_4_lut_adj_500_LC_19_22_2  (
            .in0(N__43521),
            .in1(N__46094),
            .in2(N__70338),
            .in3(N__43696),
            .lcout(),
            .ltout(\c0.n75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i44_4_lut_LC_19_22_3 .C_ON=1'b0;
    defparam \c0.i44_4_lut_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i44_4_lut_LC_19_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i44_4_lut_LC_19_22_3  (
            .in0(N__43471),
            .in1(N__43495),
            .in2(N__43489),
            .in3(N__45790),
            .lcout(),
            .ltout(\c0.n93_adj_3373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i47_4_lut_LC_19_22_4 .C_ON=1'b0;
    defparam \c0.i47_4_lut_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i47_4_lut_LC_19_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i47_4_lut_LC_19_22_4  (
            .in0(N__52774),
            .in1(N__43618),
            .in2(N__43486),
            .in3(N__57790),
            .lcout(\c0.n96_adj_3419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_390_LC_19_22_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_390_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_390_LC_19_22_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i5_2_lut_adj_390_LC_19_22_5  (
            .in0(N__48838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49397),
            .lcout(\c0.n23_adj_3222 ),
            .ltout(\c0.n23_adj_3222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_adj_498_LC_19_22_6 .C_ON=1'b0;
    defparam \c0.i27_4_lut_adj_498_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_adj_498_LC_19_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_adj_498_LC_19_22_6  (
            .in0(N__58725),
            .in1(N__59596),
            .in2(N__43474),
            .in3(N__49178),
            .lcout(\c0.n76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_287_LC_19_23_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_287_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_287_LC_19_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_287_LC_19_23_0  (
            .in0(N__53986),
            .in1(N__45270),
            .in2(N__43654),
            .in3(N__43584),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_337_LC_19_23_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_337_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_337_LC_19_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_337_LC_19_23_1  (
            .in0(N__45877),
            .in1(N__43677),
            .in2(_gnd_net_),
            .in3(N__52863),
            .lcout(\c0.n19403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_4_lut_LC_19_23_2 .C_ON=1'b0;
    defparam \c0.i12_2_lut_4_lut_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_4_lut_LC_19_23_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_2_lut_4_lut_LC_19_23_2  (
            .in0(N__52862),
            .in1(N__45876),
            .in2(N__43678),
            .in3(N__49396),
            .lcout(\c0.n38_adj_3051 ),
            .ltout(\c0.n38_adj_3051_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_3_lut_adj_448_LC_19_23_3 .C_ON=1'b0;
    defparam \c0.i19_3_lut_adj_448_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i19_3_lut_adj_448_LC_19_23_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i19_3_lut_adj_448_LC_19_23_3  (
            .in0(N__43585),
            .in1(_gnd_net_),
            .in2(N__43645),
            .in3(N__49347),
            .lcout(\c0.n45_adj_3284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_19_23_4 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_19_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_19_23_4  (
            .in0(N__43642),
            .in1(N__70279),
            .in2(N__45931),
            .in3(N__43627),
            .lcout(),
            .ltout(\c0.n51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_LC_19_23_5 .C_ON=1'b0;
    defparam \c0.i32_4_lut_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_LC_19_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_4_lut_LC_19_23_5  (
            .in0(N__43617),
            .in1(N__43600),
            .in2(N__43588),
            .in3(N__57789),
            .lcout(\c0.n32_adj_3052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_495_LC_19_23_6 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_495_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_495_LC_19_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_495_LC_19_23_6  (
            .in0(N__45271),
            .in1(N__43576),
            .in2(N__43570),
            .in3(N__45724),
            .lcout(\c0.n20930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_461_LC_19_24_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_461_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_461_LC_19_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_461_LC_19_24_0  (
            .in0(N__57255),
            .in1(N__52690),
            .in2(N__67021),
            .in3(N__44788),
            .lcout(\c0.n23_adj_3304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_458_LC_19_24_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_458_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_458_LC_19_24_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_458_LC_19_24_1  (
            .in0(N__46096),
            .in1(N__59301),
            .in2(_gnd_net_),
            .in3(N__59250),
            .lcout(),
            .ltout(\c0.n15_adj_3297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_19_24_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_19_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_19_24_2  (
            .in0(N__46207),
            .in1(N__49498),
            .in2(N__43729),
            .in3(N__52843),
            .lcout(\c0.n24_adj_3298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_4_lut_LC_19_24_3 .C_ON=1'b0;
    defparam \c0.i9_3_lut_4_lut_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_4_lut_LC_19_24_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_3_lut_4_lut_LC_19_24_3  (
            .in0(N__67618),
            .in1(N__53473),
            .in2(N__59254),
            .in3(N__49301),
            .lcout(),
            .ltout(\c0.n21_adj_3300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17661_4_lut_LC_19_24_4 .C_ON=1'b0;
    defparam \c0.i17661_4_lut_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17661_4_lut_LC_19_24_4 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.i17661_4_lut_LC_19_24_4  (
            .in0(N__53556),
            .in1(N__43726),
            .in2(N__43720),
            .in3(N__46042),
            .lcout(),
            .ltout(\c0.n21247_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_494_LC_19_24_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_494_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_494_LC_19_24_5 .LUT_INIT=16'b1101111111101111;
    LogicCell40 \c0.i6_4_lut_adj_494_LC_19_24_5  (
            .in0(N__43717),
            .in1(N__52579),
            .in2(N__43711),
            .in3(N__43708),
            .lcout(\c0.n14_adj_3354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i195_LC_19_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i195_LC_19_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i195_LC_19_25_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i195_LC_19_25_0  (
            .in0(N__46135),
            .in1(_gnd_net_),
            .in2(N__68751),
            .in3(N__70209),
            .lcout(data_in_frame_24_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71192),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i199_LC_19_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i199_LC_19_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i199_LC_19_25_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i199_LC_19_25_1  (
            .in0(N__69013),
            .in1(N__46138),
            .in2(_gnd_net_),
            .in3(N__49505),
            .lcout(data_in_frame_24_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71192),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i198_LC_19_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i198_LC_19_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i198_LC_19_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i198_LC_19_25_4  (
            .in0(N__46137),
            .in1(N__67972),
            .in2(_gnd_net_),
            .in3(N__59616),
            .lcout(data_in_frame_24_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71192),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i197_LC_19_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i197_LC_19_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i197_LC_19_25_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0__i197_LC_19_25_6  (
            .in0(N__46136),
            .in1(_gnd_net_),
            .in2(N__72755),
            .in3(N__49444),
            .lcout(data_in_frame_24_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71192),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i153_LC_19_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i153_LC_19_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i153_LC_19_25_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i153_LC_19_25_7  (
            .in0(N__69146),
            .in1(N__65217),
            .in2(_gnd_net_),
            .in3(N__45408),
            .lcout(data_in_frame_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71192),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4__5169_LC_19_26_2 .C_ON=1'b0;
    defparam \c0.data_in_3__4__5169_LC_19_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4__5169_LC_19_26_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__4__5169_LC_19_26_2  (
            .in0(N__72710),
            .in1(N__53226),
            .in2(_gnd_net_),
            .in3(N__43974),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71201),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_400_LC_19_26_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_400_LC_19_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_400_LC_19_26_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i4_4_lut_adj_400_LC_19_26_4  (
            .in0(N__43953),
            .in1(N__43886),
            .in2(N__46168),
            .in3(N__43940),
            .lcout(\c0.n10_adj_3231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i196_LC_19_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i196_LC_19_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i196_LC_19_26_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i196_LC_19_26_6  (
            .in0(N__69421),
            .in1(N__46139),
            .in2(_gnd_net_),
            .in3(N__70324),
            .lcout(data_in_frame_24_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71201),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1__5188_LC_19_27_6 .C_ON=1'b0;
    defparam \c0.data_in_1__1__5188_LC_19_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1__5188_LC_19_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__1__5188_LC_19_27_6  (
            .in0(N__53227),
            .in1(N__43915),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71213),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_98_i4_2_lut_LC_20_6_6 .C_ON=1'b0;
    defparam \c0.rx.equal_98_i4_2_lut_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_98_i4_2_lut_LC_20_6_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.equal_98_i4_2_lut_LC_20_6_6  (
            .in0(_gnd_net_),
            .in1(N__43869),
            .in2(_gnd_net_),
            .in3(N__43819),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_20_7_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_20_7_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_20_7_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i17_LC_20_7_0  (
            .in0(N__44233),
            .in1(N__61731),
            .in2(N__47216),
            .in3(N__65094),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71224),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_20_7_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_20_7_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_20_7_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_20_7_3  (
            .in0(N__43744),
            .in1(N__67777),
            .in2(N__56239),
            .in3(N__55466),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71224),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_7_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_7_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_20_7_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_20_7_5  (
            .in0(N__43755),
            .in1(N__71347),
            .in2(N__56237),
            .in3(N__55465),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71224),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_20_7_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_20_7_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_20_7_7  (
            .in0(N__43743),
            .in1(N__72531),
            .in2(N__56238),
            .in3(N__56086),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71224),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_526_LC_20_8_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_526_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_526_LC_20_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_526_LC_20_8_0  (
            .in0(N__60927),
            .in1(N__49975),
            .in2(N__44423),
            .in3(N__55382),
            .lcout(\c0.n19424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_529_LC_20_8_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_529_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_529_LC_20_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_529_LC_20_8_1  (
            .in0(N__49974),
            .in1(N__44413),
            .in2(_gnd_net_),
            .in3(N__60926),
            .lcout(\c0.n8_adj_3397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_20_8_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_20_8_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_20_8_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i31_LC_20_8_2  (
            .in0(N__69035),
            .in1(N__61430),
            .in2(N__44424),
            .in3(N__61673),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71216),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_773_LC_20_8_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_773_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_773_LC_20_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_773_LC_20_8_3  (
            .in0(_gnd_net_),
            .in1(N__56825),
            .in2(_gnd_net_),
            .in3(N__61081),
            .lcout(\c0.n9_adj_3346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_20_8_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_20_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_20_8_4  (
            .in0(N__63854),
            .in1(N__47768),
            .in2(N__64453),
            .in3(N__52107),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i39_LC_20_8_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i39_LC_20_8_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i39_LC_20_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i39_LC_20_8_5  (
            .in0(N__61671),
            .in1(N__44126),
            .in2(N__44047),
            .in3(N__69036),
            .lcout(\c0.data_in_frame_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71216),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_20_8_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_20_8_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_20_8_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i22_LC_20_8_6  (
            .in0(N__67776),
            .in1(N__61672),
            .in2(N__44395),
            .in3(N__44252),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71216),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i35_LC_20_8_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i35_LC_20_8_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i35_LC_20_8_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i35_LC_20_8_7  (
            .in0(N__61670),
            .in1(N__44125),
            .in2(N__68758),
            .in3(N__46393),
            .lcout(\c0.data_in_frame_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71216),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_705_LC_20_9_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_705_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_705_LC_20_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_705_LC_20_9_0  (
            .in0(N__46391),
            .in1(N__55212),
            .in2(N__46288),
            .in3(N__54612),
            .lcout(\c0.n7_adj_3491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_772_LC_20_9_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_772_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_772_LC_20_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_772_LC_20_9_1  (
            .in0(N__54613),
            .in1(N__46416),
            .in2(_gnd_net_),
            .in3(N__46265),
            .lcout(\c0.n9_adj_3027 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i33_LC_20_9_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i33_LC_20_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i33_LC_20_9_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i33_LC_20_9_2  (
            .in0(N__65198),
            .in1(N__61691),
            .in2(N__44128),
            .in3(N__49980),
            .lcout(\c0.data_in_frame_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71204),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i36_LC_20_9_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i36_LC_20_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i36_LC_20_9_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i36_LC_20_9_3  (
            .in0(N__61689),
            .in1(N__69424),
            .in2(N__46420),
            .in3(N__44124),
            .lcout(\c0.data_in_frame_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71204),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_20_9_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_20_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_20_9_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i20_LC_20_9_4  (
            .in0(N__69423),
            .in1(N__61690),
            .in2(N__54316),
            .in3(N__44248),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71204),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_545_LC_20_9_5 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_545_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_545_LC_20_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_545_LC_20_9_5  (
            .in0(N__44151),
            .in1(N__62131),
            .in2(N__44393),
            .in3(N__54466),
            .lcout(\c0.n4_adj_3406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i38_LC_20_9_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i38_LC_20_9_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i38_LC_20_9_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i38_LC_20_9_6  (
            .in0(N__44120),
            .in1(N__67802),
            .in2(N__47155),
            .in3(N__61692),
            .lcout(\c0.data_in_frame_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71204),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_733_LC_20_9_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_733_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_733_LC_20_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_733_LC_20_9_7  (
            .in0(N__44030),
            .in1(N__44005),
            .in2(N__43993),
            .in3(N__56801),
            .lcout(\c0.data_out_frame_0__7__N_1537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_785_LC_20_10_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_785_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_785_LC_20_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_785_LC_20_10_0  (
            .in0(N__60956),
            .in1(N__62130),
            .in2(_gnd_net_),
            .in3(N__61077),
            .lcout(\c0.n12131 ),
            .ltout(\c0.n12131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_536_LC_20_10_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_536_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_536_LC_20_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_536_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__47297),
            .in2(N__43984),
            .in3(N__62197),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_20_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_20_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_20_10_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i2_LC_20_10_2  (
            .in0(N__56823),
            .in1(N__61801),
            .in2(N__55868),
            .in3(N__71393),
            .lcout(data_in_frame_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71194),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_786_LC_20_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_786_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_786_LC_20_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_786_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(N__44304),
            .in2(_gnd_net_),
            .in3(N__62198),
            .lcout(\c0.n19415 ),
            .ltout(\c0.n19415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i36_2_lut_4_lut_LC_20_10_4 .C_ON=1'b0;
    defparam \c0.i36_2_lut_4_lut_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i36_2_lut_4_lut_LC_20_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i36_2_lut_4_lut_LC_20_10_4  (
            .in0(N__47298),
            .in1(N__55032),
            .in2(N__44284),
            .in3(N__55308),
            .lcout(\c0.n88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_736_LC_20_10_5 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_736_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_736_LC_20_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_adj_736_LC_20_10_5  (
            .in0(N__55033),
            .in1(N__54122),
            .in2(N__55309),
            .in3(N__47299),
            .lcout(\c0.n54_adj_3502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_361_LC_20_10_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_361_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_361_LC_20_10_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i4_4_lut_adj_361_LC_20_10_6  (
            .in0(N__61860),
            .in1(N__56629),
            .in2(N__62698),
            .in3(N__55732),
            .lcout(\c0.n21_adj_3205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i38_4_lut_LC_20_10_7 .C_ON=1'b0;
    defparam \c0.i38_4_lut_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i38_4_lut_LC_20_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i38_4_lut_LC_20_10_7  (
            .in0(N__47336),
            .in1(N__60957),
            .in2(N__62080),
            .in3(N__62199),
            .lcout(\c0.n90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i44_3_lut_4_lut_LC_20_11_0 .C_ON=1'b0;
    defparam \c0.i44_3_lut_4_lut_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i44_3_lut_4_lut_LC_20_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i44_3_lut_4_lut_LC_20_11_0  (
            .in0(N__54888),
            .in1(N__44271),
            .in2(N__44571),
            .in3(N__44658),
            .lcout(\c0.n96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_791_LC_20_11_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_791_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_791_LC_20_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_791_LC_20_11_2  (
            .in0(N__46334),
            .in1(N__46269),
            .in2(_gnd_net_),
            .in3(N__56802),
            .lcout(\c0.n20095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_4_lut_LC_20_11_3 .C_ON=1'b0;
    defparam \c0.i31_4_lut_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i31_4_lut_LC_20_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_4_lut_LC_20_11_3  (
            .in0(N__56803),
            .in1(N__54492),
            .in2(N__55178),
            .in3(N__54267),
            .lcout(\c0.n83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_20_11_4 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_20_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_20_11_4  (
            .in0(N__54452),
            .in1(N__62156),
            .in2(N__50406),
            .in3(N__55147),
            .lcout(\c0.n14_adj_3371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_818_LC_20_11_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_818_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_818_LC_20_11_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_818_LC_20_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47619),
            .in3(N__54054),
            .lcout(\c0.n10_adj_3538 ),
            .ltout(\c0.n10_adj_3538_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_822_LC_20_11_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_822_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_822_LC_20_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_822_LC_20_11_6  (
            .in0(N__44431),
            .in1(N__44425),
            .in2(N__44398),
            .in3(N__44394),
            .lcout(\c0.n22_adj_3356 ),
            .ltout(\c0.n22_adj_3356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_2_lut_3_lut_LC_20_11_7 .C_ON=1'b0;
    defparam \c0.i19_2_lut_3_lut_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i19_2_lut_3_lut_LC_20_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i19_2_lut_3_lut_LC_20_11_7  (
            .in0(_gnd_net_),
            .in1(N__54887),
            .in2(N__44359),
            .in3(N__47454),
            .lcout(\c0.n52_adj_3402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_20_12_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_20_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_20_12_0  (
            .in0(N__47370),
            .in1(N__44329),
            .in2(N__44344),
            .in3(N__44641),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_832_LC_20_12_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_832_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_832_LC_20_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_832_LC_20_12_1  (
            .in0(_gnd_net_),
            .in1(N__54880),
            .in2(_gnd_net_),
            .in3(N__44356),
            .lcout(\c0.n23_adj_3021 ),
            .ltout(\c0.n23_adj_3021_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_2_lut_4_lut_LC_20_12_2 .C_ON=1'b0;
    defparam \c0.i10_2_lut_4_lut_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_2_lut_4_lut_LC_20_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_2_lut_4_lut_LC_20_12_2  (
            .in0(N__50673),
            .in1(N__55587),
            .in2(N__44335),
            .in3(N__44654),
            .lcout(\c0.n26_adj_3114 ),
            .ltout(\c0.n26_adj_3114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_332_LC_20_12_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_332_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_332_LC_20_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_332_LC_20_12_3  (
            .in0(N__49951),
            .in1(N__47369),
            .in2(N__44332),
            .in3(N__44517),
            .lcout(\c0.n20981 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_758_LC_20_12_4 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_758_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_758_LC_20_12_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i4_2_lut_adj_758_LC_20_12_4  (
            .in0(N__57655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57571),
            .lcout(\c0.n12_adj_3518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_270_LC_20_12_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_270_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_270_LC_20_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_270_LC_20_12_5  (
            .in0(N__55263),
            .in1(N__60451),
            .in2(N__50158),
            .in3(N__55239),
            .lcout(\c0.n20490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_237_LC_20_12_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_237_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_237_LC_20_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_237_LC_20_12_6  (
            .in0(N__50457),
            .in1(N__44328),
            .in2(N__55291),
            .in3(N__44320),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_LC_20_12_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_LC_20_12_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i4_2_lut_3_lut_LC_20_12_7  (
            .in0(N__55586),
            .in1(_gnd_net_),
            .in2(N__44659),
            .in3(N__50672),
            .lcout(\c0.n22_adj_3022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_879_LC_20_13_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_879_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_879_LC_20_13_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_879_LC_20_13_0  (
            .in0(N__44972),
            .in1(_gnd_net_),
            .in2(N__51519),
            .in3(N__60778),
            .lcout(\c0.n11_adj_3340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_514_LC_20_13_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_514_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_514_LC_20_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_514_LC_20_13_1  (
            .in0(N__45015),
            .in1(_gnd_net_),
            .in2(N__44635),
            .in3(N__44970),
            .lcout(\c0.n18_adj_3372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_adj_616_LC_20_13_2 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_adj_616_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_adj_616_LC_20_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i9_2_lut_3_lut_adj_616_LC_20_13_2  (
            .in0(N__44971),
            .in1(_gnd_net_),
            .in2(N__44904),
            .in3(N__45016),
            .lcout(\c0.n33_adj_3289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_20_13_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_20_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_20_13_3  (
            .in0(N__44572),
            .in1(N__47356),
            .in2(N__44554),
            .in3(N__50461),
            .lcout(\c0.n20029 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_766_LC_20_13_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_766_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_766_LC_20_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_766_LC_20_13_4  (
            .in0(N__47350),
            .in1(N__44527),
            .in2(N__44521),
            .in3(N__47374),
            .lcout(\c0.n18422 ),
            .ltout(\c0.n18422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_272_LC_20_13_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_272_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_272_LC_20_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_272_LC_20_13_5  (
            .in0(N__62583),
            .in1(_gnd_net_),
            .in2(N__44488),
            .in3(N__57308),
            .lcout(\c0.n19433 ),
            .ltout(\c0.n19433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_273_LC_20_13_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_273_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_273_LC_20_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_273_LC_20_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44485),
            .in3(N__45014),
            .lcout(),
            .ltout(\c0.n11891_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_288_LC_20_13_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_288_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_288_LC_20_13_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_288_LC_20_13_7  (
            .in0(N__44465),
            .in1(N__50109),
            .in2(N__44434),
            .in3(N__57143),
            .lcout(\c0.n20151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_20_14_0 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_20_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_LC_20_14_0  (
            .in0(N__44752),
            .in1(N__44743),
            .in2(N__47508),
            .in3(N__47629),
            .lcout(\c0.n27_adj_3118 ),
            .ltout(\c0.n27_adj_3118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_2_lut_3_lut_LC_20_14_1 .C_ON=1'b0;
    defparam \c0.i11_2_lut_3_lut_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_2_lut_3_lut_LC_20_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_2_lut_3_lut_LC_20_14_1  (
            .in0(_gnd_net_),
            .in1(N__48279),
            .in2(N__44737),
            .in3(N__51942),
            .lcout(\c0.n28_adj_3245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_505_LC_20_14_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_505_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_505_LC_20_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_505_LC_20_14_2  (
            .in0(N__48033),
            .in1(N__44730),
            .in2(_gnd_net_),
            .in3(N__56561),
            .lcout(\c0.n19_adj_3336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i87_LC_20_14_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i87_LC_20_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i87_LC_20_14_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i87_LC_20_14_3  (
            .in0(N__66156),
            .in1(N__62812),
            .in2(N__66336),
            .in3(N__68903),
            .lcout(\c0.data_in_frame_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71146),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_4_lut_adj_898_LC_20_14_4 .C_ON=1'b0;
    defparam \c0.i12_2_lut_4_lut_adj_898_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_4_lut_adj_898_LC_20_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_2_lut_4_lut_adj_898_LC_20_14_4  (
            .in0(N__52040),
            .in1(N__60771),
            .in2(N__51518),
            .in3(N__44969),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_611_LC_20_14_5 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_611_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_611_LC_20_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_611_LC_20_14_5  (
            .in0(N__56562),
            .in1(N__44719),
            .in2(_gnd_net_),
            .in3(N__48034),
            .lcout(\c0.n23_adj_3364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_315_LC_20_14_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_315_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_315_LC_20_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_315_LC_20_14_7  (
            .in0(N__57191),
            .in1(_gnd_net_),
            .in2(N__65863),
            .in3(N__47745),
            .lcout(\c0.n19372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_20_15_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_20_15_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_20_15_0  (
            .in0(N__51154),
            .in1(N__56451),
            .in2(N__65350),
            .in3(N__51673),
            .lcout(\c0.n19916 ),
            .ltout(\c0.n19916_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_LC_20_15_1 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_LC_20_15_1 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i9_2_lut_3_lut_LC_20_15_1  (
            .in0(N__44671),
            .in1(N__44805),
            .in2(N__44662),
            .in3(_gnd_net_),
            .lcout(\c0.n22_adj_3341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_LC_20_15_2 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_LC_20_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_LC_20_15_2  (
            .in0(N__64628),
            .in1(N__65853),
            .in2(N__48219),
            .in3(N__48261),
            .lcout(\c0.n21_adj_3337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_831_LC_20_15_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_831_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_831_LC_20_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_831_LC_20_15_3  (
            .in0(N__50739),
            .in1(N__56743),
            .in2(N__50784),
            .in3(N__44827),
            .lcout(\c0.n19477 ),
            .ltout(\c0.n19477_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_20_15_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_20_15_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_20_15_4  (
            .in0(N__63049),
            .in1(N__56450),
            .in2(N__44818),
            .in3(N__51672),
            .lcout(),
            .ltout(\c0.n12_adj_3348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_659_LC_20_15_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_659_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_659_LC_20_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_659_LC_20_15_5  (
            .in0(N__65343),
            .in1(N__57443),
            .in2(N__44815),
            .in3(N__47887),
            .lcout(\c0.n21045 ),
            .ltout(\c0.n21045_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_640_LC_20_15_6 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_640_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_640_LC_20_15_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i6_2_lut_adj_640_LC_20_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44812),
            .in3(N__52758),
            .lcout(\c0.n19_adj_3303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_adj_875_LC_20_16_0 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_adj_875_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_adj_875_LC_20_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_2_lut_3_lut_adj_875_LC_20_16_0  (
            .in0(N__60793),
            .in1(N__44979),
            .in2(_gnd_net_),
            .in3(N__44809),
            .lcout(\c0.n40_adj_3366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i177_LC_20_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i177_LC_20_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i177_LC_20_16_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i177_LC_20_16_1  (
            .in0(N__65262),
            .in1(N__67530),
            .in2(_gnd_net_),
            .in3(N__70037),
            .lcout(data_in_frame_22_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71115),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_645_LC_20_16_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_645_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_645_LC_20_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_645_LC_20_16_2  (
            .in0(N__49136),
            .in1(N__44775),
            .in2(N__57235),
            .in3(N__52722),
            .lcout(\c0.n20085 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_20_16_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_20_16_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_LC_20_16_3  (
            .in0(N__44764),
            .in1(N__55668),
            .in2(N__45069),
            .in3(N__48510),
            .lcout(\c0.n21110 ),
            .ltout(\c0.n21110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_654_LC_20_16_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_654_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_654_LC_20_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_654_LC_20_16_4  (
            .in0(N__45154),
            .in1(N__45142),
            .in2(N__45100),
            .in3(N__45097),
            .lcout(\c0.n40_adj_3413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i113_LC_20_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i113_LC_20_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i113_LC_20_16_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i113_LC_20_16_5  (
            .in0(N__65263),
            .in1(N__64238),
            .in2(N__62048),
            .in3(N__57225),
            .lcout(\c0.data_in_frame_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71115),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i116_LC_20_16_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i116_LC_20_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i116_LC_20_16_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i116_LC_20_16_6  (
            .in0(N__64237),
            .in1(N__62035),
            .in2(N__45070),
            .in3(N__69315),
            .lcout(\c0.data_in_frame_14_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71115),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_2_lut_3_lut_LC_20_17_0 .C_ON=1'b0;
    defparam \c0.i16_2_lut_3_lut_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_2_lut_3_lut_LC_20_17_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i16_2_lut_3_lut_LC_20_17_0  (
            .in0(N__44986),
            .in1(_gnd_net_),
            .in2(N__64014),
            .in3(N__45021),
            .lcout(\c0.n67_adj_3063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_3_lut_4_lut_LC_20_17_1 .C_ON=1'b0;
    defparam \c0.i17_3_lut_4_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_3_lut_4_lut_LC_20_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_3_lut_4_lut_LC_20_17_1  (
            .in0(N__45020),
            .in1(N__44985),
            .in2(N__44947),
            .in3(N__48933),
            .lcout(\c0.n43_adj_3330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_755_LC_20_17_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_755_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_755_LC_20_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_755_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__64833),
            .in2(_gnd_net_),
            .in3(N__67378),
            .lcout(),
            .ltout(\c0.n12_adj_3517_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_765_LC_20_17_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_765_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_765_LC_20_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_765_LC_20_17_3  (
            .in0(N__57709),
            .in1(N__44920),
            .in2(N__44908),
            .in3(N__69082),
            .lcout(\c0.n20512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_665_LC_20_17_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_665_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_665_LC_20_17_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_665_LC_20_17_4  (
            .in0(N__45702),
            .in1(N__53414),
            .in2(N__44905),
            .in3(N__45577),
            .lcout(\c0.n20840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_847_LC_20_17_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_847_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_847_LC_20_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_847_LC_20_17_5  (
            .in0(N__44848),
            .in1(N__51912),
            .in2(N__44839),
            .in3(N__52053),
            .lcout(\c0.n20451 ),
            .ltout(\c0.n20451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_569_LC_20_17_6 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_569_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_569_LC_20_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_569_LC_20_17_6  (
            .in0(N__69080),
            .in1(N__64832),
            .in2(N__45253),
            .in3(N__45810),
            .lcout(\c0.n15_adj_3432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_387_LC_20_17_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_387_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_387_LC_20_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_387_LC_20_17_7  (
            .in0(N__67379),
            .in1(N__45250),
            .in2(N__45814),
            .in3(N__69081),
            .lcout(\c0.n13_adj_3221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_4_lut_adj_738_LC_20_18_0 .C_ON=1'b0;
    defparam \c0.i31_4_lut_adj_738_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i31_4_lut_adj_738_LC_20_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_4_lut_adj_738_LC_20_18_0  (
            .in0(N__48869),
            .in1(N__49098),
            .in2(N__48102),
            .in3(N__57511),
            .lcout(\c0.n64_adj_3512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_870_LC_20_18_1 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_870_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_870_LC_20_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i4_2_lut_adj_870_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(N__57455),
            .in2(_gnd_net_),
            .in3(N__45179),
            .lcout(),
            .ltout(\c0.n27_adj_3529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_802_LC_20_18_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_802_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_802_LC_20_18_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_802_LC_20_18_2  (
            .in0(N__45238),
            .in1(N__62950),
            .in2(N__45220),
            .in3(N__51685),
            .lcout(),
            .ltout(\c0.n32_adj_3530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_811_LC_20_18_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_811_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_811_LC_20_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_811_LC_20_18_3  (
            .in0(N__47941),
            .in1(N__47704),
            .in2(N__45217),
            .in3(N__56470),
            .lcout(\c0.n19244 ),
            .ltout(\c0.n19244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_2_lut_3_lut_LC_20_18_4 .C_ON=1'b0;
    defparam \c0.i24_2_lut_3_lut_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i24_2_lut_3_lut_LC_20_18_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i24_2_lut_3_lut_LC_20_18_4  (
            .in0(N__45290),
            .in1(_gnd_net_),
            .in2(N__45214),
            .in3(N__67657),
            .lcout(\c0.n85_adj_3074 ),
            .ltout(\c0.n85_adj_3074_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_650_LC_20_18_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_650_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_650_LC_20_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_650_LC_20_18_5  (
            .in0(N__45334),
            .in1(N__45180),
            .in2(N__45199),
            .in3(N__45196),
            .lcout(\c0.n13_adj_3244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_3_lut_4_lut_LC_20_18_6 .C_ON=1'b0;
    defparam \c0.i21_3_lut_4_lut_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i21_3_lut_4_lut_LC_20_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_3_lut_4_lut_LC_20_18_6  (
            .in0(N__45181),
            .in1(N__47834),
            .in2(N__57460),
            .in3(N__51687),
            .lcout(\c0.n49_adj_3358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_2_lut_adj_644_LC_20_18_7 .C_ON=1'b0;
    defparam \c0.i16_2_lut_adj_644_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i16_2_lut_adj_644_LC_20_18_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i16_2_lut_adj_644_LC_20_18_7  (
            .in0(N__51686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57456),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_788_LC_20_19_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_788_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_788_LC_20_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_788_LC_20_19_0  (
            .in0(N__63994),
            .in1(N__67288),
            .in2(N__67434),
            .in3(N__51885),
            .lcout(\c0.n30_adj_3392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_3_lut_LC_20_19_1 .C_ON=1'b0;
    defparam \c0.i15_2_lut_3_lut_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_3_lut_LC_20_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i15_2_lut_3_lut_LC_20_19_1  (
            .in0(N__65520),
            .in1(N__47835),
            .in2(_gnd_net_),
            .in3(N__59074),
            .lcout(\c0.n48_adj_3409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_775_LC_20_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_775_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_775_LC_20_19_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_775_LC_20_19_2  (
            .in0(N__72474),
            .in1(_gnd_net_),
            .in2(N__66421),
            .in3(_gnd_net_),
            .lcout(\c0.n4_adj_3522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i168_LC_20_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i168_LC_20_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i168_LC_20_19_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i168_LC_20_19_3  (
            .in0(N__71791),
            .in1(N__70147),
            .in2(N__67219),
            .in3(N__72221),
            .lcout(\c0.data_in_frame_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71130),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_20_19_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_20_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_20_19_4  (
            .in0(N__59075),
            .in1(N__65521),
            .in2(_gnd_net_),
            .in3(N__58024),
            .lcout(\c0.n22_adj_3287 ),
            .ltout(\c0.n22_adj_3287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_895_LC_20_19_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_895_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_895_LC_20_19_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_895_LC_20_19_5  (
            .in0(N__67289),
            .in1(N__63995),
            .in2(N__45274),
            .in3(N__57547),
            .lcout(\c0.n10_adj_3555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_672_LC_20_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_672_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_672_LC_20_19_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_672_LC_20_19_6  (
            .in0(N__70126),
            .in1(_gnd_net_),
            .in2(N__70154),
            .in3(_gnd_net_),
            .lcout(\c0.n19223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_3_lut_adj_869_LC_20_19_7 .C_ON=1'b0;
    defparam \c0.i13_2_lut_3_lut_adj_869_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_3_lut_adj_869_LC_20_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i13_2_lut_3_lut_adj_869_LC_20_19_7  (
            .in0(N__68165),
            .in1(N__66417),
            .in2(_gnd_net_),
            .in3(N__72475),
            .lcout(\c0.n39_adj_3050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_adj_560_LC_20_20_0 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_adj_560_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_adj_560_LC_20_20_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_3_lut_4_lut_adj_560_LC_20_20_0  (
            .in0(N__57656),
            .in1(N__59126),
            .in2(N__57724),
            .in3(N__57581),
            .lcout(\c0.n14_adj_3421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_591_LC_20_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_591_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_591_LC_20_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_591_LC_20_20_1  (
            .in0(_gnd_net_),
            .in1(N__45638),
            .in2(_gnd_net_),
            .in3(N__45704),
            .lcout(\c0.n19384 ),
            .ltout(\c0.n19384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_621_LC_20_20_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_621_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_621_LC_20_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_621_LC_20_20_2  (
            .in0(N__45484),
            .in1(N__45475),
            .in2(N__45463),
            .in3(N__45661),
            .lcout(\c0.n17819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_20_20_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_4_lut_LC_20_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_2_lut_3_lut_4_lut_LC_20_20_3  (
            .in0(N__64892),
            .in1(N__48377),
            .in2(N__45452),
            .in3(N__45703),
            .lcout(\c0.n9_adj_3430 ),
            .ltout(\c0.n9_adj_3430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_590_LC_20_20_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_590_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_590_LC_20_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_590_LC_20_20_4  (
            .in0(N__45412),
            .in1(N__45366),
            .in2(N__45394),
            .in3(N__45390),
            .lcout(\c0.n20431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_751_LC_20_20_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_751_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_751_LC_20_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_751_LC_20_20_5  (
            .in0(N__45391),
            .in1(N__45376),
            .in2(N__45370),
            .in3(N__59345),
            .lcout(\c0.n18433 ),
            .ltout(\c0.n18433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_474_LC_20_20_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_474_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_474_LC_20_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_474_LC_20_20_6  (
            .in0(N__53907),
            .in1(N__66381),
            .in2(N__45358),
            .in3(N__67639),
            .lcout(\c0.n40_adj_3323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_710_LC_20_20_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_710_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_710_LC_20_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_710_LC_20_20_7  (
            .in0(N__57582),
            .in1(N__57713),
            .in2(_gnd_net_),
            .in3(N__57657),
            .lcout(\c0.n20479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_632_LC_20_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_632_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_632_LC_20_21_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_632_LC_20_21_0  (
            .in0(N__45355),
            .in1(N__53963),
            .in2(N__45639),
            .in3(N__45713),
            .lcout(\c0.n4_adj_3123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_661_LC_20_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_661_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_661_LC_20_21_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_661_LC_20_21_1  (
            .in0(N__59073),
            .in1(_gnd_net_),
            .in2(N__63777),
            .in3(_gnd_net_),
            .lcout(\c0.n19511 ),
            .ltout(\c0.n19511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_633_LC_20_21_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_633_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_633_LC_20_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_633_LC_20_21_2  (
            .in0(N__45633),
            .in1(N__58839),
            .in2(N__45718),
            .in3(N__45714),
            .lcout(\c0.n7_adj_3054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i193_LC_20_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i193_LC_20_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i193_LC_20_21_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i193_LC_20_21_3  (
            .in0(N__65248),
            .in1(N__46153),
            .in2(_gnd_net_),
            .in3(N__58756),
            .lcout(data_in_frame_24_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71160),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_597_LC_20_21_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_597_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_597_LC_20_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i10_4_lut_adj_597_LC_20_21_4  (
            .in0(N__57658),
            .in1(N__45673),
            .in2(N__65281),
            .in3(N__45660),
            .lcout(\c0.n22_adj_3450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_adj_740_LC_20_21_5 .C_ON=1'b0;
    defparam \c0.i32_4_lut_adj_740_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_adj_740_LC_20_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_4_lut_adj_740_LC_20_21_5  (
            .in0(N__45649),
            .in1(N__58084),
            .in2(N__59149),
            .in3(N__48544),
            .lcout(\c0.n21071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_579_LC_20_21_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_579_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_579_LC_20_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_579_LC_20_21_6  (
            .in0(N__45629),
            .in1(N__63767),
            .in2(_gnd_net_),
            .in3(N__59072),
            .lcout(\c0.n7_adj_3440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i105_LC_20_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i105_LC_20_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i105_LC_20_21_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i105_LC_20_21_7  (
            .in0(N__65249),
            .in1(N__71965),
            .in2(N__66211),
            .in3(N__45560),
            .lcout(\c0.data_in_frame_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71160),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_388_LC_20_22_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_388_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_388_LC_20_22_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_388_LC_20_22_0  (
            .in0(N__68434),
            .in1(N__69835),
            .in2(N__45541),
            .in3(N__45523),
            .lcout(\c0.n18431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_637_LC_20_22_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_637_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_637_LC_20_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_637_LC_20_22_1  (
            .in0(N__71283),
            .in1(N__45514),
            .in2(N__69907),
            .in3(N__52444),
            .lcout(\c0.n20324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_3_lut_LC_20_22_2 .C_ON=1'b0;
    defparam \c0.i15_3_lut_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_3_lut_LC_20_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i15_3_lut_LC_20_22_2  (
            .in0(N__46177),
            .in1(N__48534),
            .in2(_gnd_net_),
            .in3(N__45496),
            .lcout(\c0.n21044 ),
            .ltout(\c0.n21044_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_328_LC_20_22_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_328_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_328_LC_20_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_328_LC_20_22_3  (
            .in0(N__53602),
            .in1(N__47098),
            .in2(N__45880),
            .in3(N__58761),
            .lcout(),
            .ltout(\c0.n16_adj_3109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_333_LC_20_22_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_333_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_333_LC_20_22_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_4_lut_adj_333_LC_20_22_4  (
            .in0(N__45869),
            .in1(N__49411),
            .in2(N__45829),
            .in3(N__45826),
            .lcout(\c0.n21076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_585_LC_20_22_5 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_585_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_585_LC_20_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_585_LC_20_22_5  (
            .in0(_gnd_net_),
            .in1(N__64830),
            .in2(_gnd_net_),
            .in3(N__45804),
            .lcout(\c0.n9_adj_3069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_adj_499_LC_20_23_0 .C_ON=1'b0;
    defparam \c0.i28_4_lut_adj_499_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_adj_499_LC_20_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i28_4_lut_adj_499_LC_20_23_0  (
            .in0(N__49765),
            .in1(N__47086),
            .in2(N__49348),
            .in3(N__49371),
            .lcout(\c0.n77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_320_LC_20_23_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_320_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_320_LC_20_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_320_LC_20_23_1  (
            .in0(N__45784),
            .in1(N__45765),
            .in2(N__51759),
            .in3(N__49017),
            .lcout(\c0.n18457 ),
            .ltout(\c0.n18457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_445_LC_20_23_2 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_445_LC_20_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_445_LC_20_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_445_LC_20_23_2  (
            .in0(N__52646),
            .in1(N__53586),
            .in2(N__45748),
            .in3(N__46053),
            .lcout(\c0.n41_adj_3281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_444_LC_20_23_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_444_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_444_LC_20_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_444_LC_20_23_3  (
            .in0(N__59833),
            .in1(N__52599),
            .in2(N__53824),
            .in3(N__45744),
            .lcout(),
            .ltout(\c0.n43_adj_3280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_447_LC_20_23_4 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_447_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_447_LC_20_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_447_LC_20_23_4  (
            .in0(N__53442),
            .in1(N__49354),
            .in2(N__45733),
            .in3(N__45730),
            .lcout(\c0.n50_adj_3283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_466_LC_20_23_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_466_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_466_LC_20_23_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_4_lut_adj_466_LC_20_23_5  (
            .in0(N__46102),
            .in1(N__46093),
            .in2(N__46057),
            .in3(N__52647),
            .lcout(\c0.n33_adj_3308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_318_LC_20_24_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_318_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_318_LC_20_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_318_LC_20_24_0  (
            .in0(N__49491),
            .in1(N__52864),
            .in2(N__46206),
            .in3(N__52689),
            .lcout(\c0.n18417 ),
            .ltout(\c0.n18417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_453_LC_20_24_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_453_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_453_LC_20_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_453_LC_20_24_1  (
            .in0(N__46035),
            .in1(N__48619),
            .in2(N__46045),
            .in3(N__52651),
            .lcout(\c0.n19_adj_3292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i237_LC_20_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i237_LC_20_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i237_LC_20_24_2 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i237_LC_20_24_2  (
            .in0(N__72744),
            .in1(N__46036),
            .in2(N__66975),
            .in3(N__71934),
            .lcout(\c0.data_in_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71195),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i235_LC_20_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i235_LC_20_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i235_LC_20_24_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i235_LC_20_24_3  (
            .in0(N__71932),
            .in1(N__68744),
            .in2(N__46023),
            .in3(N__66942),
            .lcout(\c0.data_in_frame_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71195),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i234_LC_20_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i234_LC_20_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i234_LC_20_24_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i234_LC_20_24_4  (
            .in0(N__71534),
            .in1(N__45999),
            .in2(N__66974),
            .in3(N__71933),
            .lcout(\c0.data_in_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71195),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i226_LC_20_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i226_LC_20_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i226_LC_20_24_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i226_LC_20_24_5  (
            .in0(N__45975),
            .in1(N__71535),
            .in2(N__67222),
            .in3(N__66941),
            .lcout(\c0.data_in_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71195),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i225_LC_20_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i225_LC_20_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i225_LC_20_24_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i225_LC_20_24_6  (
            .in0(N__66934),
            .in1(N__67200),
            .in2(N__45955),
            .in3(N__65261),
            .lcout(\c0.data_in_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71195),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_486_LC_20_24_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_486_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_486_LC_20_24_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_486_LC_20_24_7  (
            .in0(N__59560),
            .in1(N__53842),
            .in2(N__45954),
            .in3(N__45936),
            .lcout(\c0.n14_adj_3349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_308_LC_20_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_308_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_308_LC_20_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_308_LC_20_25_0  (
            .in0(_gnd_net_),
            .in1(N__49326),
            .in2(_gnd_net_),
            .in3(N__53383),
            .lcout(\c0.n7_adj_3078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i136_LC_20_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i136_LC_20_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i136_LC_20_25_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i136_LC_20_25_1  (
            .in0(N__72294),
            .in1(N__65596),
            .in2(_gnd_net_),
            .in3(N__57692),
            .lcout(data_in_frame_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71203),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i141_LC_20_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i141_LC_20_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i141_LC_20_25_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i141_LC_20_25_2  (
            .in0(N__71762),
            .in1(N__63358),
            .in2(N__64760),
            .in3(N__72729),
            .lcout(\c0.data_in_frame_17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71203),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i203_LC_20_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i203_LC_20_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i203_LC_20_25_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i203_LC_20_25_3  (
            .in0(N__68740),
            .in1(N__49259),
            .in2(N__63389),
            .in3(N__66973),
            .lcout(\c0.data_in_frame_25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71203),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_776_LC_20_25_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_776_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_776_LC_20_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_776_LC_20_25_4  (
            .in0(N__46189),
            .in1(N__53942),
            .in2(N__72397),
            .in3(N__53974),
            .lcout(\c0.n26_adj_3523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i202_LC_20_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i202_LC_20_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i202_LC_20_25_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i202_LC_20_25_5  (
            .in0(N__49327),
            .in1(N__71543),
            .in2(N__63390),
            .in3(N__66972),
            .lcout(\c0.data_in_frame_25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71203),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_540_LC_20_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_540_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_540_LC_20_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_540_LC_20_25_7  (
            .in0(_gnd_net_),
            .in1(N__59612),
            .in2(_gnd_net_),
            .in3(N__49435),
            .lcout(\c0.n11865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4__5193_LC_20_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0__4__5193_LC_20_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4__5193_LC_20_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__4__5193_LC_20_26_1  (
            .in0(N__53229),
            .in1(N__46993),
            .in2(_gnd_net_),
            .in3(N__46167),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71215),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3848_2_lut_LC_20_26_2 .C_ON=1'b0;
    defparam \c0.i3848_2_lut_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3848_2_lut_LC_20_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3848_2_lut_LC_20_26_2  (
            .in0(_gnd_net_),
            .in1(N__49487),
            .in2(_gnd_net_),
            .in3(N__53618),
            .lcout(\c0.n6495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i200_LC_20_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i200_LC_20_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i200_LC_20_26_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i200_LC_20_26_4  (
            .in0(N__53622),
            .in1(N__46152),
            .in2(_gnd_net_),
            .in3(N__72291),
            .lcout(data_in_frame_24_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71215),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_543_LC_20_26_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_543_LC_20_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_543_LC_20_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_543_LC_20_26_6  (
            .in0(N__70375),
            .in1(N__70314),
            .in2(_gnd_net_),
            .in3(N__70208),
            .lcout(\c0.n12085 ),
            .ltout(\c0.n12085_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_787_LC_20_26_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_787_LC_20_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_787_LC_20_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_787_LC_20_26_7  (
            .in0(_gnd_net_),
            .in1(N__47082),
            .in2(N__47071),
            .in3(N__47052),
            .lcout(\c0.n19274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4__5185_LC_20_27_1 .C_ON=1'b0;
    defparam \c0.data_in_1__4__5185_LC_20_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4__5185_LC_20_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__4__5185_LC_20_27_1  (
            .in0(N__53228),
            .in1(N__46992),
            .in2(_gnd_net_),
            .in3(N__47041),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71223),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_223_LC_21_7_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_223_LC_21_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_223_LC_21_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_223_LC_21_7_6  (
            .in0(N__51015),
            .in1(N__54750),
            .in2(_gnd_net_),
            .in3(N__50989),
            .lcout(\c0.n19291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__7__5207_LC_21_8_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__7__5207_LC_21_8_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__7__5207_LC_21_8_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__7__5207_LC_21_8_1  (
            .in0(N__46963),
            .in1(N__62176),
            .in2(N__55186),
            .in3(N__50339),
            .lcout(\c0.data_out_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71225),
            .ce(N__46936),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_717_LC_21_8_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_717_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_717_LC_21_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_717_LC_21_8_2  (
            .in0(N__46415),
            .in1(N__46392),
            .in2(N__46368),
            .in3(N__47205),
            .lcout(),
            .ltout(\c0.n13_adj_3496_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_721_LC_21_8_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_721_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_721_LC_21_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_721_LC_21_8_3  (
            .in0(N__46213),
            .in1(N__49692),
            .in2(N__46348),
            .in3(N__46341),
            .lcout(\c0.n5_adj_3031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_713_LC_21_8_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_713_LC_21_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_713_LC_21_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_713_LC_21_8_4  (
            .in0(_gnd_net_),
            .in1(N__46301),
            .in2(_gnd_net_),
            .in3(N__56824),
            .lcout(\c0.n19277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_777_LC_21_8_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_777_LC_21_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_777_LC_21_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_777_LC_21_8_6  (
            .in0(N__49691),
            .in1(N__47206),
            .in2(N__47182),
            .in3(N__55383),
            .lcout(\c0.n20391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_780_LC_21_9_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_780_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_780_LC_21_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_780_LC_21_9_0  (
            .in0(N__60450),
            .in1(N__51054),
            .in2(_gnd_net_),
            .in3(N__55235),
            .lcout(\c0.n11833 ),
            .ltout(\c0.n11833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i40_4_lut_LC_21_9_1 .C_ON=1'b0;
    defparam \c0.i40_4_lut_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i40_4_lut_LC_21_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i40_4_lut_LC_21_9_1  (
            .in0(N__66287),
            .in1(N__47167),
            .in2(N__47173),
            .in3(N__47116),
            .lcout(),
            .ltout(\c0.n92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i46_4_lut_LC_21_9_2 .C_ON=1'b0;
    defparam \c0.i46_4_lut_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i46_4_lut_LC_21_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i46_4_lut_LC_21_9_2  (
            .in0(N__47161),
            .in1(N__50230),
            .in2(N__47170),
            .in3(N__62165),
            .lcout(\c0.n98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_21_9_3 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_21_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i28_4_lut_LC_21_9_3  (
            .in0(N__49847),
            .in1(N__56378),
            .in2(N__49875),
            .in3(N__54518),
            .lcout(\c0.n80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_692_LC_21_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_692_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_692_LC_21_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_692_LC_21_9_4  (
            .in0(_gnd_net_),
            .in1(N__50332),
            .in2(_gnd_net_),
            .in3(N__50405),
            .lcout(\c0.n19196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_836_LC_21_9_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_836_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_836_LC_21_9_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_836_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(N__49979),
            .in2(_gnd_net_),
            .in3(N__61197),
            .lcout(\c0.n5_adj_3030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_792_LC_21_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_792_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_792_LC_21_9_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_792_LC_21_9_6  (
            .in0(N__54262),
            .in1(_gnd_net_),
            .in2(N__47154),
            .in3(_gnd_net_),
            .lcout(\c0.n19241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_900_LC_21_9_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_900_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_900_LC_21_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_900_LC_21_9_7  (
            .in0(N__62582),
            .in1(N__47145),
            .in2(_gnd_net_),
            .in3(N__54261),
            .lcout(\c0.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i51_4_lut_LC_21_10_0 .C_ON=1'b0;
    defparam \c0.i51_4_lut_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i51_4_lut_LC_21_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i51_4_lut_LC_21_10_0  (
            .in0(N__47110),
            .in1(N__49990),
            .in2(N__47404),
            .in3(N__47104),
            .lcout(\c0.n12_adj_3034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_adj_840_LC_21_10_1 .C_ON=1'b0;
    defparam \c0.i8_2_lut_adj_840_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_adj_840_LC_21_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i8_2_lut_adj_840_LC_21_10_1  (
            .in0(N__54094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61194),
            .lcout(\c0.n24_adj_3013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i66_LC_21_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i66_LC_21_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i66_LC_21_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i66_LC_21_10_2  (
            .in0(N__64255),
            .in1(N__55883),
            .in2(N__51520),
            .in3(N__71376),
            .lcout(\c0.data_in_frame_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71205),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_604_LC_21_10_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_604_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_604_LC_21_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i2_2_lut_adj_604_LC_21_10_3  (
            .in0(N__50301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55034),
            .lcout(\c0.n7_adj_3029 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_551_LC_21_10_4 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_551_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_551_LC_21_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_551_LC_21_10_4  (
            .in0(N__61196),
            .in1(N__54096),
            .in2(N__50434),
            .in3(N__50300),
            .lcout(\c0.n20313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17690_4_lut_LC_21_10_5 .C_ON=1'b0;
    defparam \c0.i17690_4_lut_LC_21_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17690_4_lut_LC_21_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17690_4_lut_LC_21_10_5  (
            .in0(N__54097),
            .in1(N__50602),
            .in2(N__60988),
            .in3(N__61118),
            .lcout(\c0.n21277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_652_LC_21_10_6 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_652_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_652_LC_21_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_2_lut_3_lut_4_lut_adj_652_LC_21_10_6  (
            .in0(N__61195),
            .in1(N__54095),
            .in2(N__54894),
            .in3(N__54674),
            .lcout(),
            .ltout(\c0.n14_adj_3476_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_701_LC_21_10_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_701_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_701_LC_21_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_701_LC_21_10_7  (
            .in0(N__50601),
            .in1(N__47296),
            .in2(N__47281),
            .in3(N__55284),
            .lcout(\c0.n19966 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_306_LC_21_11_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_306_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_306_LC_21_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_306_LC_21_11_0  (
            .in0(N__55610),
            .in1(N__47227),
            .in2(N__50005),
            .in3(N__47274),
            .lcout(\c0.n30_adj_3075 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_305_LC_21_11_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_305_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_305_LC_21_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_305_LC_21_11_1  (
            .in0(_gnd_net_),
            .in1(N__55919),
            .in2(_gnd_net_),
            .in3(N__51097),
            .lcout(\c0.n19508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_833_LC_21_11_2 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_833_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_833_LC_21_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_833_LC_21_11_2  (
            .in0(N__51287),
            .in1(N__55127),
            .in2(N__51414),
            .in3(N__47476),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_LC_21_11_3 .C_ON=1'b0;
    defparam \c0.i15_2_lut_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_LC_21_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i15_2_lut_LC_21_11_3  (
            .in0(_gnd_net_),
            .in1(N__60488),
            .in2(_gnd_net_),
            .in3(N__56291),
            .lcout(),
            .ltout(\c0.n67_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i48_4_lut_LC_21_11_4 .C_ON=1'b0;
    defparam \c0.i48_4_lut_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i48_4_lut_LC_21_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i48_4_lut_LC_21_11_4  (
            .in0(N__47470),
            .in1(N__47461),
            .in2(N__47443),
            .in3(N__47440),
            .lcout(),
            .ltout(\c0.n100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i50_4_lut_LC_21_11_5 .C_ON=1'b0;
    defparam \c0.i50_4_lut_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i50_4_lut_LC_21_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i50_4_lut_LC_21_11_5  (
            .in0(N__47434),
            .in1(N__47424),
            .in2(N__47407),
            .in3(N__49930),
            .lcout(\c0.n102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_236_LC_21_11_7 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_236_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_236_LC_21_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_236_LC_21_11_7  (
            .in0(_gnd_net_),
            .in1(N__56290),
            .in2(_gnd_net_),
            .in3(N__47395),
            .lcout(\c0.n21_adj_3010 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_4_lut_adj_624_LC_21_12_0 .C_ON=1'b0;
    defparam \c0.i10_3_lut_4_lut_adj_624_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_4_lut_adj_624_LC_21_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_3_lut_4_lut_adj_624_LC_21_12_0  (
            .in0(N__50175),
            .in1(N__54531),
            .in2(N__60493),
            .in3(N__54727),
            .lcout(\c0.n28_adj_3023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_735_LC_21_12_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_735_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_735_LC_21_12_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_735_LC_21_12_1  (
            .in0(N__54532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60492),
            .lcout(\c0.n17_adj_3508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i89_LC_21_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i89_LC_21_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i89_LC_21_12_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i89_LC_21_12_2  (
            .in0(N__64502),
            .in1(N__66154),
            .in2(N__53657),
            .in3(N__65202),
            .lcout(\c0.data_in_frame_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71183),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_307_LC_21_12_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_307_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_307_LC_21_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_307_LC_21_12_4  (
            .in0(N__47340),
            .in1(N__54461),
            .in2(N__54567),
            .in3(N__47317),
            .lcout(),
            .ltout(\c0.n32_adj_3077_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_314_LC_21_12_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_314_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_314_LC_21_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_314_LC_21_12_5  (
            .in0(N__50486),
            .in1(N__50063),
            .in2(N__47656),
            .in3(N__50836),
            .lcout(\c0.n21047 ),
            .ltout(\c0.n21047_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_330_LC_21_12_6 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_330_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_330_LC_21_12_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i18_4_lut_adj_330_LC_21_12_6  (
            .in0(N__64449),
            .in1(N__47646),
            .in2(N__47632),
            .in3(N__54462),
            .lcout(\c0.n42_adj_3111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_2_lut_3_lut_LC_21_12_7 .C_ON=1'b0;
    defparam \c0.i17_2_lut_3_lut_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17_2_lut_3_lut_LC_21_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i17_2_lut_3_lut_LC_21_12_7  (
            .in0(N__50485),
            .in1(N__47620),
            .in2(_gnd_net_),
            .in3(N__47555),
            .lcout(\c0.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_239_LC_21_13_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_239_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_239_LC_21_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_239_LC_21_13_0  (
            .in0(N__66326),
            .in1(N__54155),
            .in2(N__53658),
            .in3(N__57091),
            .lcout(),
            .ltout(\c0.n10_adj_3014_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_240_LC_21_13_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_240_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_240_LC_21_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_240_LC_21_13_1  (
            .in0(_gnd_net_),
            .in1(N__49558),
            .in2(N__47512),
            .in3(N__56957),
            .lcout(\c0.n19456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i127_LC_21_13_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i127_LC_21_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i127_LC_21_13_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i127_LC_21_13_2  (
            .in0(N__64411),
            .in1(N__64247),
            .in2(N__47886),
            .in3(N__68927),
            .lcout(\c0.data_in_frame_15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71172),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_21_13_3 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_21_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_LC_21_13_3  (
            .in0(N__47490),
            .in1(N__50191),
            .in2(N__50081),
            .in3(N__50797),
            .lcout(\c0.n16_adj_3218 ),
            .ltout(\c0.n16_adj_3218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_873_LC_21_13_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_873_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_873_LC_21_13_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_873_LC_21_13_4  (
            .in0(N__51540),
            .in1(_gnd_net_),
            .in2(N__47479),
            .in3(N__58432),
            .lcout(\c0.n12_adj_3469 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i71_LC_21_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i71_LC_21_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i71_LC_21_13_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i71_LC_21_13_5  (
            .in0(N__64246),
            .in1(N__55876),
            .in2(N__68973),
            .in3(N__49559),
            .lcout(\c0.data_in_frame_8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71172),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_21_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_21_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_LC_21_13_6  (
            .in0(_gnd_net_),
            .in1(N__63232),
            .in2(_gnd_net_),
            .in3(N__57372),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i69_LC_21_13_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i69_LC_21_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i69_LC_21_13_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i69_LC_21_13_7  (
            .in0(N__64245),
            .in1(N__55875),
            .in2(N__56971),
            .in3(N__72659),
            .lcout(\c0.data_in_frame_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71172),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i72_LC_21_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i72_LC_21_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i72_LC_21_14_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i72_LC_21_14_0  (
            .in0(N__64243),
            .in1(N__55873),
            .in2(N__54162),
            .in3(N__72255),
            .lcout(\c0.data_in_frame_8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71161),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i99_LC_21_14_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i99_LC_21_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i99_LC_21_14_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i99_LC_21_14_1  (
            .in0(N__68594),
            .in1(N__67118),
            .in2(N__47767),
            .in3(N__66155),
            .lcout(\c0.data_in_frame_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71161),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i70_LC_21_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i70_LC_21_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i70_LC_21_14_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i70_LC_21_14_2  (
            .in0(N__64242),
            .in1(N__67854),
            .in2(N__57114),
            .in3(N__55874),
            .lcout(\c0.data_in_frame_8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71161),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_874_LC_21_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_874_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_874_LC_21_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_874_LC_21_14_3  (
            .in0(_gnd_net_),
            .in1(N__65515),
            .in2(_gnd_net_),
            .in3(N__59085),
            .lcout(\c0.n5_adj_3549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_804_LC_21_14_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_804_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_804_LC_21_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_804_LC_21_14_4  (
            .in0(N__57107),
            .in1(N__57024),
            .in2(N__56731),
            .in3(N__47722),
            .lcout(\c0.n30_adj_3531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i68_LC_21_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i68_LC_21_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i68_LC_21_14_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i68_LC_21_14_5  (
            .in0(N__55872),
            .in1(N__64244),
            .in2(N__58467),
            .in3(N__69409),
            .lcout(\c0.data_in_frame_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71161),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_adj_563_LC_21_14_6 .C_ON=1'b0;
    defparam \c0.i9_2_lut_adj_563_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_adj_563_LC_21_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i9_2_lut_adj_563_LC_21_14_6  (
            .in0(_gnd_net_),
            .in1(N__51436),
            .in2(_gnd_net_),
            .in3(N__47688),
            .lcout(\c0.n42_adj_3367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_3_lut_adj_806_LC_21_14_7 .C_ON=1'b0;
    defparam \c0.i13_3_lut_adj_806_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_3_lut_adj_806_LC_21_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i13_3_lut_adj_806_LC_21_14_7  (
            .in0(N__54021),
            .in1(N__49699),
            .in2(_gnd_net_),
            .in3(N__49858),
            .lcout(\c0.n31_adj_3532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_487_LC_21_15_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_487_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_487_LC_21_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_487_LC_21_15_0  (
            .in0(N__62257),
            .in1(N__47926),
            .in2(N__62313),
            .in3(N__56652),
            .lcout(\c0.n9_adj_3350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_281_LC_21_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_281_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_281_LC_21_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_281_LC_21_15_1  (
            .in0(_gnd_net_),
            .in1(N__48334),
            .in2(_gnd_net_),
            .in3(N__55952),
            .lcout(\c0.n11942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_668_LC_21_15_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_668_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_668_LC_21_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_668_LC_21_15_3  (
            .in0(N__47885),
            .in1(N__56726),
            .in2(N__56533),
            .in3(N__65292),
            .lcout(),
            .ltout(\c0.n16_adj_3481_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_670_LC_21_15_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_670_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_670_LC_21_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_670_LC_21_15_4  (
            .in0(N__51139),
            .in1(N__47850),
            .in2(N__47857),
            .in3(N__63109),
            .lcout(\c0.n11815 ),
            .ltout(\c0.n11815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_673_LC_21_15_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_673_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_673_LC_21_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_673_LC_21_15_5  (
            .in0(N__58353),
            .in1(N__66244),
            .in2(N__47854),
            .in3(N__58131),
            .lcout(\c0.n10_adj_3483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_21_15_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_21_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_21_15_6  (
            .in0(N__51043),
            .in1(N__51033),
            .in2(N__63700),
            .in3(N__47851),
            .lcout(\c0.n11632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_2_lut_3_lut_adj_720_LC_21_16_0 .C_ON=1'b0;
    defparam \c0.i18_2_lut_3_lut_adj_720_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_2_lut_3_lut_adj_720_LC_21_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i18_2_lut_3_lut_adj_720_LC_21_16_0  (
            .in0(N__62992),
            .in1(_gnd_net_),
            .in2(N__47836),
            .in3(N__47779),
            .lcout(\c0.n35_adj_3266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_933_LC_21_16_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_933_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_933_LC_21_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_933_LC_21_16_1  (
            .in0(N__56668),
            .in1(N__56484),
            .in2(N__63013),
            .in3(N__65434),
            .lcout(\c0.n12056 ),
            .ltout(\c0.n12056_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_21_16_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_21_16_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_21_16_2  (
            .in0(N__58931),
            .in1(N__59133),
            .in2(N__47782),
            .in3(N__56528),
            .lcout(\c0.n12_adj_3249 ),
            .ltout(\c0.n12_adj_3249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_681_LC_21_16_3 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_681_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_681_LC_21_16_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_681_LC_21_16_3  (
            .in0(N__68383),
            .in1(_gnd_net_),
            .in2(N__48043),
            .in3(N__52351),
            .lcout(\c0.n36_adj_3452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_667_LC_21_16_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_667_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_667_LC_21_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_667_LC_21_16_4  (
            .in0(N__51208),
            .in1(N__48040),
            .in2(N__69475),
            .in3(N__65325),
            .lcout(\c0.n19524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_285_LC_21_16_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_285_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_285_LC_21_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_285_LC_21_16_5  (
            .in0(N__51214),
            .in1(N__58130),
            .in2(N__62314),
            .in3(N__57267),
            .lcout(\c0.n19301 ),
            .ltout(\c0.n19301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_828_LC_21_16_6 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_828_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_828_LC_21_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i3_2_lut_adj_828_LC_21_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48007),
            .in3(N__56566),
            .lcout(\c0.n9_adj_3240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_3_lut_4_lut_LC_21_17_0 .C_ON=1'b0;
    defparam \c0.i12_2_lut_3_lut_4_lut_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_3_lut_4_lut_LC_21_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_2_lut_3_lut_4_lut_LC_21_17_0  (
            .in0(N__48130),
            .in1(N__47975),
            .in2(N__48000),
            .in3(N__48930),
            .lcout(\c0.n31_adj_3126 ),
            .ltout(\c0.n31_adj_3126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_2_lut_4_lut_LC_21_17_1 .C_ON=1'b0;
    defparam \c0.i16_2_lut_4_lut_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_2_lut_4_lut_LC_21_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_2_lut_4_lut_LC_21_17_1  (
            .in0(N__63678),
            .in1(N__52184),
            .in2(N__48004),
            .in3(N__52158),
            .lcout(\c0.n35_adj_3317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_2_lut_3_lut_LC_21_17_2 .C_ON=1'b0;
    defparam \c0.i18_2_lut_3_lut_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i18_2_lut_3_lut_LC_21_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i18_2_lut_3_lut_LC_21_17_2  (
            .in0(N__52185),
            .in1(_gnd_net_),
            .in2(N__48001),
            .in3(N__47976),
            .lcout(\c0.n46 ),
            .ltout(\c0.n46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_3_lut_4_lut_LC_21_17_3 .C_ON=1'b0;
    defparam \c0.i32_3_lut_4_lut_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i32_3_lut_4_lut_LC_21_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_3_lut_4_lut_LC_21_17_3  (
            .in0(N__63679),
            .in1(N__47956),
            .in2(N__47944),
            .in3(N__52159),
            .lcout(\c0.n69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_2_lut_3_lut_LC_21_17_4 .C_ON=1'b0;
    defparam \c0.i25_2_lut_3_lut_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_2_lut_3_lut_LC_21_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i25_2_lut_3_lut_LC_21_17_4  (
            .in0(N__48131),
            .in1(N__48721),
            .in2(_gnd_net_),
            .in3(N__48931),
            .lcout(\c0.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_adj_451_LC_21_17_5 .C_ON=1'b0;
    defparam \c0.i23_4_lut_adj_451_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_adj_451_LC_21_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_adj_451_LC_21_17_5  (
            .in0(N__48722),
            .in1(N__48139),
            .in2(N__64018),
            .in3(N__48132),
            .lcout(\c0.n51_adj_3290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_3_lut_LC_21_17_6 .C_ON=1'b0;
    defparam \c0.i13_2_lut_3_lut_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_3_lut_LC_21_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i13_2_lut_3_lut_LC_21_17_6  (
            .in0(N__64056),
            .in1(N__57502),
            .in2(_gnd_net_),
            .in3(N__58998),
            .lcout(\c0.n6_adj_3137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_21_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_21_17_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_937_LC_21_17_7  (
            .in0(N__71793),
            .in1(N__55867),
            .in2(_gnd_net_),
            .in3(N__59478),
            .lcout(n19130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_2_lut_3_lut_LC_21_18_0 .C_ON=1'b0;
    defparam \c0.i33_2_lut_3_lut_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i33_2_lut_3_lut_LC_21_18_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i33_2_lut_3_lut_LC_21_18_0  (
            .in0(N__52879),
            .in1(_gnd_net_),
            .in2(N__58550),
            .in3(N__59046),
            .lcout(\c0.n84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_605_LC_21_18_1 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_605_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_605_LC_21_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_605_LC_21_18_1  (
            .in0(N__57969),
            .in1(N__58954),
            .in2(N__52399),
            .in3(N__52362),
            .lcout(\c0.n19824 ),
            .ltout(\c0.n19824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_501_LC_21_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_501_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_501_LC_21_18_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_501_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48085),
            .in3(N__69986),
            .lcout(),
            .ltout(\c0.n18_adj_3360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_503_LC_21_18_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_503_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_503_LC_21_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_503_LC_21_18_3  (
            .in0(N__51637),
            .in1(N__48081),
            .in2(N__48052),
            .in3(N__52019),
            .lcout(),
            .ltout(\c0.n32_adj_3362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_506_LC_21_18_4 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_506_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_506_LC_21_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_506_LC_21_18_4  (
            .in0(N__51972),
            .in1(N__52261),
            .in2(N__48049),
            .in3(N__48960),
            .lcout(\c0.n20112 ),
            .ltout(\c0.n20112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_517_LC_21_18_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_517_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_517_LC_21_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_517_LC_21_18_5  (
            .in0(N__65626),
            .in1(N__52134),
            .in2(N__48046),
            .in3(N__48932),
            .lcout(\c0.n51_adj_3376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_484_LC_21_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_484_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_484_LC_21_19_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_484_LC_21_19_0  (
            .in0(N__64623),
            .in1(N__48333),
            .in2(N__64708),
            .in3(N__55960),
            .lcout(\c0.n18398 ),
            .ltout(\c0.n18398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_622_LC_21_19_1 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_622_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_622_LC_21_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_622_LC_21_19_1  (
            .in0(N__64984),
            .in1(_gnd_net_),
            .in2(N__48304),
            .in3(N__64951),
            .lcout(\c0.n37_adj_3390 ),
            .ltout(\c0.n37_adj_3390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_LC_21_19_2 .C_ON=1'b0;
    defparam \c0.i9_3_lut_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_LC_21_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i9_3_lut_LC_21_19_2  (
            .in0(N__65722),
            .in1(_gnd_net_),
            .in2(N__48301),
            .in3(N__49143),
            .lcout(\c0.n25_adj_3431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_adj_507_LC_21_19_3 .C_ON=1'b0;
    defparam \c0.i27_4_lut_adj_507_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_adj_507_LC_21_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_adj_507_LC_21_19_3  (
            .in0(N__48193),
            .in1(N__48163),
            .in2(N__51457),
            .in3(N__48232),
            .lcout(),
            .ltout(\c0.n60_adj_3368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_adj_522_LC_21_19_4 .C_ON=1'b0;
    defparam \c0.i30_4_lut_adj_522_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_adj_522_LC_21_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i30_4_lut_adj_522_LC_21_19_4  (
            .in0(N__48298),
            .in1(N__48226),
            .in2(N__48292),
            .in3(N__48289),
            .lcout(\c0.n63_adj_3391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_LC_21_19_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_LC_21_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_LC_21_19_5  (
            .in0(N__48283),
            .in1(N__64624),
            .in2(_gnd_net_),
            .in3(N__48265),
            .lcout(\c0.n39_adj_3334 ),
            .ltout(\c0.n39_adj_3334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_568_LC_21_19_6 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_568_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_568_LC_21_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_568_LC_21_19_6  (
            .in0(N__48145),
            .in1(N__48225),
            .in2(N__48202),
            .in3(N__48199),
            .lcout(\c0.n17900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_565_LC_21_19_7 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_565_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_565_LC_21_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_565_LC_21_19_7  (
            .in0(N__48192),
            .in1(N__48181),
            .in2(N__51456),
            .in3(N__48162),
            .lcout(\c0.n30_adj_3429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_894_LC_21_20_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_894_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_894_LC_21_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_894_LC_21_20_0  (
            .in0(N__53751),
            .in1(N__58895),
            .in2(_gnd_net_),
            .in3(N__53494),
            .lcout(\c0.n35_adj_3274 ),
            .ltout(\c0.n35_adj_3274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_adj_739_LC_21_20_1 .C_ON=1'b0;
    defparam \c0.i26_4_lut_adj_739_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_adj_739_LC_21_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_adj_739_LC_21_20_1  (
            .in0(N__58247),
            .in1(N__58217),
            .in2(N__48547),
            .in3(N__58199),
            .lcout(\c0.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_21_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_21_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_21_20_2  (
            .in0(N__68227),
            .in1(N__68120),
            .in2(_gnd_net_),
            .in3(N__48527),
            .lcout(\c0.n11601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_825_LC_21_20_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_825_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_825_LC_21_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_825_LC_21_20_3  (
            .in0(N__57196),
            .in1(N__48511),
            .in2(N__55978),
            .in3(N__48490),
            .lcout(\c0.n12052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i40_4_lut_adj_438_LC_21_20_4 .C_ON=1'b0;
    defparam \c0.i40_4_lut_adj_438_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i40_4_lut_adj_438_LC_21_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i40_4_lut_adj_438_LC_21_20_4  (
            .in0(N__57987),
            .in1(N__58248),
            .in2(N__48451),
            .in3(N__48666),
            .lcout(\c0.n91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_628_LC_21_20_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_628_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_628_LC_21_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i5_2_lut_adj_628_LC_21_20_5  (
            .in0(N__58832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57747),
            .lcout(\c0.n38_adj_3270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i40_4_lut_adj_521_LC_21_20_6 .C_ON=1'b0;
    defparam \c0.i40_4_lut_adj_521_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i40_4_lut_adj_521_LC_21_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i40_4_lut_adj_521_LC_21_20_6  (
            .in0(N__57988),
            .in1(N__48450),
            .in2(N__68047),
            .in3(N__48667),
            .lcout(\c0.n91_adj_3389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_2_lut_4_lut_LC_21_21_0 .C_ON=1'b0;
    defparam \c0.i22_2_lut_4_lut_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i22_2_lut_4_lut_LC_21_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_2_lut_4_lut_LC_21_21_0  (
            .in0(N__48724),
            .in1(N__58649),
            .in2(N__69715),
            .in3(N__68022),
            .lcout(\c0.n49_adj_3316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_598_LC_21_21_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_598_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_598_LC_21_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_4_lut_adj_598_LC_21_21_1  (
            .in0(N__48436),
            .in1(N__48412),
            .in2(N__57732),
            .in3(N__48391),
            .lcout(\c0.n24_adj_3427 ),
            .ltout(\c0.n24_adj_3427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_3_lut_LC_21_21_2 .C_ON=1'b0;
    defparam \c0.i8_2_lut_3_lut_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_3_lut_LC_21_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i8_2_lut_3_lut_LC_21_21_2  (
            .in0(_gnd_net_),
            .in1(N__64899),
            .in2(N__48385),
            .in3(N__48382),
            .lcout(\c0.n32_adj_3057 ),
            .ltout(\c0.n32_adj_3057_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_2_lut_LC_21_21_3 .C_ON=1'b0;
    defparam \c0.i17_2_lut_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_2_lut_LC_21_21_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i17_2_lut_LC_21_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48727),
            .in3(N__48723),
            .lcout(\c0.n44_adj_3125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_896_LC_21_21_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_896_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_896_LC_21_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_896_LC_21_21_4  (
            .in0(N__68169),
            .in1(N__48697),
            .in2(N__48688),
            .in3(N__49401),
            .lcout(\c0.n55_adj_3273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_748_LC_21_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_748_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_748_LC_21_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_748_LC_21_21_5  (
            .in0(N__52338),
            .in1(N__68430),
            .in2(_gnd_net_),
            .in3(N__48658),
            .lcout(\c0.n20965 ),
            .ltout(\c0.n20965_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_767_LC_21_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_767_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_767_LC_21_21_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_767_LC_21_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48634),
            .in3(N__65781),
            .lcout(\c0.n19312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_478_LC_21_22_0 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_478_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_478_LC_21_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_478_LC_21_22_0  (
            .in0(N__48631),
            .in1(N__51786),
            .in2(N__63457),
            .in3(N__49087),
            .lcout(\c0.n20336 ),
            .ltout(\c0.n20336_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_456_LC_21_22_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_456_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_456_LC_21_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_4_lut_adj_456_LC_21_22_1  (
            .in0(N__48618),
            .in1(N__53587),
            .in2(N__48574),
            .in3(N__52446),
            .lcout(\c0.n30_adj_3295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_adj_523_LC_21_22_2 .C_ON=1'b0;
    defparam \c0.i32_4_lut_adj_523_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_adj_523_LC_21_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_4_lut_adj_523_LC_21_22_2  (
            .in0(N__48571),
            .in1(N__49111),
            .in2(N__63456),
            .in3(N__48559),
            .lcout(\c0.n21034 ),
            .ltout(\c0.n21034_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_493_LC_21_22_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_493_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_493_LC_21_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_493_LC_21_22_3  (
            .in0(_gnd_net_),
            .in1(N__52482),
            .in2(N__48550),
            .in3(N__52505),
            .lcout(\c0.n18377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_520_LC_21_22_4 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_520_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_520_LC_21_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_520_LC_21_22_4  (
            .in0(N__49147),
            .in1(N__53874),
            .in2(N__70165),
            .in3(N__51785),
            .lcout(\c0.n58_adj_3381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_3_lut_LC_21_22_5 .C_ON=1'b0;
    defparam \c0.i24_3_lut_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i24_3_lut_LC_21_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i24_3_lut_LC_21_22_5  (
            .in0(N__48876),
            .in1(N__58491),
            .in2(_gnd_net_),
            .in3(N__49105),
            .lcout(\c0.n50_adj_3331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_adj_440_LC_21_22_6 .C_ON=1'b0;
    defparam \c0.i13_2_lut_adj_440_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_adj_440_LC_21_22_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i13_2_lut_adj_440_LC_21_22_6  (
            .in0(_gnd_net_),
            .in1(N__48907),
            .in2(_gnd_net_),
            .in3(N__49080),
            .lcout(\c0.n33_adj_3097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_406_LC_21_23_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_406_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_406_LC_21_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_406_LC_21_23_0  (
            .in0(N__64949),
            .in1(N__58912),
            .in2(N__49006),
            .in3(N__48991),
            .lcout(),
            .ltout(\c0.n27_adj_3241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_409_LC_21_23_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_409_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_409_LC_21_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_409_LC_21_23_1  (
            .in0(N__48979),
            .in1(N__48964),
            .in2(N__48943),
            .in3(N__48940),
            .lcout(\c0.n19_adj_3135 ),
            .ltout(\c0.n19_adj_3135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_adj_347_LC_21_23_2 .C_ON=1'b0;
    defparam \c0.i8_2_lut_adj_347_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_adj_347_LC_21_23_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i8_2_lut_adj_347_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48901),
            .in3(N__48898),
            .lcout(),
            .ltout(\c0.n22_adj_3136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_348_LC_21_23_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_348_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_348_LC_21_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_348_LC_21_23_3  (
            .in0(N__63455),
            .in1(N__48880),
            .in2(N__48844),
            .in3(N__51787),
            .lcout(\c0.n11936 ),
            .ltout(\c0.n11936_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_700_LC_21_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_700_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_700_LC_21_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_700_LC_21_23_4  (
            .in0(N__49260),
            .in1(N__49227),
            .in2(N__48841),
            .in3(N__48837),
            .lcout(\c0.n20_adj_3293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_472_LC_21_23_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_472_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_472_LC_21_23_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_472_LC_21_23_5  (
            .in0(N__49536),
            .in1(N__48790),
            .in2(N__49182),
            .in3(N__52447),
            .lcout(\c0.n17_adj_3318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_774_LC_21_23_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_774_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_774_LC_21_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_774_LC_21_23_6  (
            .in0(N__49261),
            .in1(N__49228),
            .in2(N__59701),
            .in3(N__49535),
            .lcout(\c0.n12_adj_3141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_326_LC_21_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_326_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_326_LC_21_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_326_LC_21_24_1  (
            .in0(_gnd_net_),
            .in1(N__49506),
            .in2(_gnd_net_),
            .in3(N__49454),
            .lcout(),
            .ltout(\c0.n19465_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_331_LC_21_24_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_331_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_331_LC_21_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_331_LC_21_24_2  (
            .in0(N__68157),
            .in1(N__53280),
            .in2(N__49414),
            .in3(N__53837),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_379_LC_21_24_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_379_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_379_LC_21_24_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_379_LC_21_24_3  (
            .in0(N__53838),
            .in1(N__68158),
            .in2(N__53284),
            .in3(N__49402),
            .lcout(\c0.n19703 ),
            .ltout(\c0.n19703_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_443_LC_21_24_4 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_443_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_443_LC_21_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_443_LC_21_24_4  (
            .in0(N__49160),
            .in1(N__58715),
            .in2(N__49357),
            .in3(N__59588),
            .lcout(\c0.n44_adj_3278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_319_LC_21_24_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_319_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_319_LC_21_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_319_LC_21_24_5  (
            .in0(_gnd_net_),
            .in1(N__49328),
            .in2(_gnd_net_),
            .in3(N__49257),
            .lcout(\c0.n7_adj_3094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_adj_756_LC_21_24_7 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_adj_756_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_adj_756_LC_21_24_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i7_2_lut_3_lut_adj_756_LC_21_24_7  (
            .in0(N__69988),
            .in1(N__72859),
            .in2(_gnd_net_),
            .in3(N__49288),
            .lcout(\c0.n33_adj_3279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_381_LC_21_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_381_LC_21_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_381_LC_21_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_381_LC_21_25_2  (
            .in0(_gnd_net_),
            .in1(N__49258),
            .in2(_gnd_net_),
            .in3(N__49229),
            .lcout(\c0.n19400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_LC_21_25_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_LC_21_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_LC_21_25_3  (
            .in0(N__53768),
            .in1(N__70044),
            .in2(_gnd_net_),
            .in3(N__66395),
            .lcout(\c0.n36_adj_3275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_291_LC_21_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_291_LC_21_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_291_LC_21_25_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_291_LC_21_25_4  (
            .in0(N__49789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53255),
            .lcout(\c0.n17840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i185_LC_21_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i185_LC_21_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i185_LC_21_25_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i185_LC_21_25_5  (
            .in0(N__53769),
            .in1(N__65247),
            .in2(_gnd_net_),
            .in3(N__53721),
            .lcout(data_in_frame_23_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71217),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0__5173_LC_21_25_6 .C_ON=1'b0;
    defparam \c0.data_in_3__0__5173_LC_21_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0__5173_LC_21_25_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__0__5173_LC_21_25_6  (
            .in0(N__65246),
            .in1(N__53230),
            .in2(_gnd_net_),
            .in3(N__49730),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71217),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i192_LC_21_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i192_LC_21_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i192_LC_21_25_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i192_LC_21_25_7  (
            .in0(N__72293),
            .in1(N__53722),
            .in2(_gnd_net_),
            .in3(N__66396),
            .lcout(data_in_frame_23_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71217),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_769_LC_22_8_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_769_LC_22_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_769_LC_22_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_769_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__54842),
            .in2(_gnd_net_),
            .in3(N__54673),
            .lcout(\c0.n12_adj_3498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_5_i6_2_lut_LC_22_8_3 .C_ON=1'b0;
    defparam \c0.select_357_Select_5_i6_2_lut_LC_22_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_5_i6_2_lut_LC_22_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_5_i6_2_lut_LC_22_8_3  (
            .in0(_gnd_net_),
            .in1(N__49676),
            .in2(_gnd_net_),
            .in3(N__60729),
            .lcout(\c0.n6_adj_3149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_911_LC_22_8_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_911_LC_22_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_911_LC_22_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_911_LC_22_8_5  (
            .in0(N__54199),
            .in1(N__57005),
            .in2(N__49581),
            .in3(N__56399),
            .lcout(\c0.n13_adj_3344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_adj_907_LC_22_8_7 .C_ON=1'b0;
    defparam \c0.i7_2_lut_adj_907_LC_22_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_adj_907_LC_22_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i7_2_lut_adj_907_LC_22_8_7  (
            .in0(N__49577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57006),
            .lcout(\c0.n35_adj_3233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_837_LC_22_9_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_837_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_837_LC_22_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_837_LC_22_9_0  (
            .in0(N__62625),
            .in1(N__61198),
            .in2(N__49984),
            .in3(N__60908),
            .lcout(\c0.n17_adj_3113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_3_lut_adj_901_LC_22_9_1 .C_ON=1'b0;
    defparam \c0.i8_2_lut_3_lut_adj_901_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_3_lut_adj_901_LC_22_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i8_2_lut_3_lut_adj_901_LC_22_9_1  (
            .in0(N__54675),
            .in1(N__54308),
            .in2(_gnd_net_),
            .in3(N__54770),
            .lcout(\c0.n60 ),
            .ltout(\c0.n60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i41_4_lut_LC_22_9_2 .C_ON=1'b0;
    defparam \c0.i41_4_lut_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i41_4_lut_LC_22_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i41_4_lut_LC_22_9_2  (
            .in0(N__57004),
            .in1(N__49939),
            .in2(N__49933),
            .in3(N__54901),
            .lcout(\c0.n93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_22_9_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_22_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_22_9_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_frame_0__i16_LC_22_9_3  (
            .in0(N__72200),
            .in1(_gnd_net_),
            .in2(N__54684),
            .in3(N__59883),
            .lcout(data_in_frame_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71226),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_763_LC_22_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_763_LC_22_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_763_LC_22_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_763_LC_22_9_4  (
            .in0(_gnd_net_),
            .in1(N__49916),
            .in2(_gnd_net_),
            .in3(N__54851),
            .lcout(\c0.n5_adj_3028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_22_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_22_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i52_LC_22_9_5  (
            .in0(N__62009),
            .in1(N__61598),
            .in2(N__54022),
            .in3(N__69443),
            .lcout(\c0.data_in_frame_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71226),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_770_LC_22_9_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_770_LC_22_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_770_LC_22_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_770_LC_22_9_6  (
            .in0(N__54771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54676),
            .lcout(\c0.n7_adj_3520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_760_LC_22_9_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_760_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_760_LC_22_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_760_LC_22_9_7  (
            .in0(N__55584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55349),
            .lcout(\c0.n19443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_764_LC_22_10_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_764_LC_22_10_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_764_LC_22_10_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_764_LC_22_10_0  (
            .in0(N__61347),
            .in1(_gnd_net_),
            .in2(N__49809),
            .in3(N__55544),
            .lcout(\c0.n11687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_848_LC_22_10_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_848_LC_22_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_848_LC_22_10_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_848_LC_22_10_1  (
            .in0(N__62354),
            .in1(N__49802),
            .in2(N__55548),
            .in3(N__61346),
            .lcout(),
            .ltout(\c0.n8_adj_3066_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_292_LC_22_10_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_292_LC_22_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_292_LC_22_10_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_292_LC_22_10_2  (
            .in0(N__51478),
            .in1(N__55725),
            .in2(N__50185),
            .in3(N__60906),
            .lcout(\c0.n19170 ),
            .ltout(\c0.n19170_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_839_LC_22_10_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_839_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_839_LC_22_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_839_LC_22_10_3  (
            .in0(_gnd_net_),
            .in1(N__62399),
            .in2(N__50161),
            .in3(N__50150),
            .lcout(\c0.n21_adj_3053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_843_LC_22_10_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_843_LC_22_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_843_LC_22_10_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_843_LC_22_10_4  (
            .in0(N__54836),
            .in1(N__55015),
            .in2(N__55162),
            .in3(N__60905),
            .lcout(\c0.n15_adj_3545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_612_LC_22_10_5 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_612_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_612_LC_22_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_612_LC_22_10_5  (
            .in0(N__55016),
            .in1(N__61254),
            .in2(_gnd_net_),
            .in3(N__50313),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_22_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_22_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_22_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_22_10_6  (
            .in0(N__54126),
            .in1(N__59876),
            .in2(_gnd_net_),
            .in3(N__71419),
            .lcout(data_in_frame_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71218),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_22_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_22_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i12_LC_22_10_7  (
            .in0(N__59875),
            .in1(N__69425),
            .in2(_gnd_net_),
            .in3(N__61212),
            .lcout(data_in_frame_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71218),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_706_LC_22_11_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_706_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_706_LC_22_11_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_706_LC_22_11_0  (
            .in0(N__50022),
            .in1(N__50394),
            .in2(N__50432),
            .in3(N__50285),
            .lcout(\c0.n20340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i37_3_lut_LC_22_11_1 .C_ON=1'b0;
    defparam \c0.i37_3_lut_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i37_3_lut_LC_22_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i37_3_lut_LC_22_11_1  (
            .in0(N__55505),
            .in1(N__61205),
            .in2(_gnd_net_),
            .in3(N__50004),
            .lcout(\c0.n89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_22_11_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_22_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_22_11_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i28_LC_22_11_2  (
            .in0(N__61408),
            .in1(N__69438),
            .in2(N__50433),
            .in3(N__61744),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71206),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_22_11_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_22_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_22_11_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i27_LC_22_11_3  (
            .in0(N__50395),
            .in1(N__68674),
            .in2(N__61777),
            .in3(N__61407),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71206),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_615_LC_22_11_4 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_615_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_615_LC_22_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_615_LC_22_11_4  (
            .in0(N__50674),
            .in1(N__55128),
            .in2(_gnd_net_),
            .in3(N__50603),
            .lcout(\c0.n33_adj_3088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_22_11_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_22_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_22_11_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i8_LC_22_11_5  (
            .in0(N__72199),
            .in1(N__50361),
            .in2(N__61778),
            .in3(N__55885),
            .lcout(data_out_frame_29__3__N_647),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71206),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_22_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_22_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_22_11_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i7_LC_22_11_6  (
            .in0(N__55884),
            .in1(N__55129),
            .in2(N__68854),
            .in3(N__61745),
            .lcout(data_in_frame_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71206),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_845_LC_22_11_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_845_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_845_LC_22_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_845_LC_22_11_7  (
            .in0(N__50467),
            .in1(N__55724),
            .in2(N__50456),
            .in3(N__50425),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_419_LC_22_12_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_419_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_419_LC_22_12_0 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \c0.i1_2_lut_adj_419_LC_22_12_0  (
            .in0(N__59485),
            .in1(_gnd_net_),
            .in2(N__61424),
            .in3(_gnd_net_),
            .lcout(\c0.n19131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_576_LC_22_12_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_576_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_576_LC_22_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_576_LC_22_12_1  (
            .in0(N__50393),
            .in1(N__55109),
            .in2(_gnd_net_),
            .in3(N__50286),
            .lcout(\c0.n29_adj_3216 ),
            .ltout(\c0.n29_adj_3216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_22_12_2 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_22_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_22_12_2  (
            .in0(N__50226),
            .in1(N__50209),
            .in2(N__50194),
            .in3(N__50869),
            .lcout(\c0.n44_adj_3217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_382_LC_22_12_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_382_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_382_LC_22_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_382_LC_22_12_3  (
            .in0(N__50853),
            .in1(N__50933),
            .in2(N__57633),
            .in3(N__50977),
            .lcout(),
            .ltout(\c0.n36_adj_3212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_384_LC_22_12_4 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_384_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_384_LC_22_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_384_LC_22_12_4  (
            .in0(N__54966),
            .in1(N__55696),
            .in2(N__50872),
            .in3(N__54460),
            .lcout(\c0.n41_adj_3213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_722_LC_22_12_5 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_722_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_722_LC_22_12_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i4_2_lut_adj_722_LC_22_12_5  (
            .in0(N__50852),
            .in1(N__54965),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n11651 ),
            .ltout(\c0.n11651_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_LC_22_12_6 .C_ON=1'b0;
    defparam \c0.i10_3_lut_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_LC_22_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i10_3_lut_LC_22_12_6  (
            .in0(_gnd_net_),
            .in1(N__55697),
            .in2(N__50839),
            .in3(N__50796),
            .lcout(\c0.n27_adj_3082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_adj_380_LC_22_12_7 .C_ON=1'b0;
    defparam \c0.i8_2_lut_adj_380_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_adj_380_LC_22_12_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i8_2_lut_adj_380_LC_22_12_7  (
            .in0(N__51090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50822),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_394_LC_22_13_0 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_394_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_394_LC_22_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_394_LC_22_13_0  (
            .in0(N__51421),
            .in1(N__62889),
            .in2(N__50785),
            .in3(N__56848),
            .lcout(),
            .ltout(\c0.n52_adj_3223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_LC_22_13_1 .C_ON=1'b0;
    defparam \c0.i26_4_lut_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_LC_22_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_LC_22_13_1  (
            .in0(N__50749),
            .in1(N__50740),
            .in2(N__50716),
            .in3(N__56365),
            .lcout(\c0.n54_adj_3234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_22_13_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_22_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_22_13_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i63_LC_22_13_2  (
            .in0(N__61766),
            .in1(N__64413),
            .in2(N__56351),
            .in3(N__68825),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71184),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_4_lut_adj_732_LC_22_13_3 .C_ON=1'b0;
    defparam \c0.i32_4_lut_adj_732_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.i32_4_lut_adj_732_LC_22_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i32_4_lut_adj_732_LC_22_13_3  (
            .in0(N__54937),
            .in1(N__56272),
            .in2(N__50713),
            .in3(N__50698),
            .lcout(\c0.n46_adj_3443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i183_LC_22_13_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i183_LC_22_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i183_LC_22_13_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i183_LC_22_13_4  (
            .in0(N__53794),
            .in1(N__67531),
            .in2(_gnd_net_),
            .in3(N__68824),
            .lcout(data_in_frame_22_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71184),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_22_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_22_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_22_13_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i61_LC_22_13_5  (
            .in0(N__64412),
            .in1(N__61767),
            .in2(N__51104),
            .in3(N__72660),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71184),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_22_13_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_22_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_22_13_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i62_LC_22_13_7  (
            .in0(N__67948),
            .in1(N__61768),
            .in2(N__55708),
            .in3(N__64414),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71184),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i85_LC_22_14_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i85_LC_22_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i85_LC_22_14_0 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0__i85_LC_22_14_0  (
            .in0(N__51539),
            .in1(N__62810),
            .in2(N__66066),
            .in3(N__72738),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71173),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_3_lut_adj_878_LC_22_14_1 .C_ON=1'b0;
    defparam \c0.i12_2_lut_3_lut_adj_878_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_3_lut_adj_878_LC_22_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i12_2_lut_3_lut_adj_878_LC_22_14_1  (
            .in0(N__58431),
            .in1(N__51538),
            .in2(_gnd_net_),
            .in3(N__51061),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_222_LC_22_14_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_222_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_222_LC_22_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_222_LC_22_14_2  (
            .in0(_gnd_net_),
            .in1(N__65407),
            .in2(_gnd_net_),
            .in3(N__61285),
            .lcout(\c0.n4 ),
            .ltout(\c0.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_876_LC_22_14_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_876_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_876_LC_22_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_876_LC_22_14_3  (
            .in0(N__51037),
            .in1(N__51016),
            .in2(N__50992),
            .in3(N__50988),
            .lcout(\c0.n26_adj_3550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i81_LC_22_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i81_LC_22_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i81_LC_22_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i81_LC_22_14_4  (
            .in0(N__62830),
            .in1(N__66184),
            .in2(N__50937),
            .in3(N__65118),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71173),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i109_LC_22_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i109_LC_22_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i109_LC_22_14_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i109_LC_22_14_5  (
            .in0(N__72739),
            .in1(N__71970),
            .in2(N__63048),
            .in3(N__66007),
            .lcout(\c0.data_in_frame_13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71173),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i169_LC_22_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i169_LC_22_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i169_LC_22_14_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i169_LC_22_14_6  (
            .in0(N__71969),
            .in1(N__71800),
            .in2(N__50903),
            .in3(N__65117),
            .lcout(\c0.data_in_frame_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71173),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_393_LC_22_14_7 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_393_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_393_LC_22_14_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_393_LC_22_14_7  (
            .in0(N__51432),
            .in1(N__51711),
            .in2(N__63799),
            .in3(N__58599),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_880_LC_22_15_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_880_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_880_LC_22_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_880_LC_22_15_0  (
            .in0(N__51415),
            .in1(N__51349),
            .in2(N__51301),
            .in3(N__51292),
            .lcout(\c0.n27_adj_3551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i86_LC_22_15_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i86_LC_22_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i86_LC_22_15_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i86_LC_22_15_1  (
            .in0(N__56904),
            .in1(N__67947),
            .in2(N__66204),
            .in3(N__62844),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71162),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_280_LC_22_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_280_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_280_LC_22_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_280_LC_22_15_2  (
            .in0(N__63034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51706),
            .lcout(\c0.n11613 ),
            .ltout(\c0.n11613_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_669_LC_22_15_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_669_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_669_LC_22_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_669_LC_22_15_3  (
            .in0(N__51207),
            .in1(N__51178),
            .in2(N__51157),
            .in3(N__51153),
            .lcout(\c0.n17_adj_3482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3106_2_lut_LC_22_15_4 .C_ON=1'b0;
    defparam \c0.i3106_2_lut_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3106_2_lut_LC_22_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3106_2_lut_LC_22_15_4  (
            .in0(_gnd_net_),
            .in1(N__51122),
            .in2(_gnd_net_),
            .in3(N__56027),
            .lcout(\c0.n5753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i111_LC_22_15_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i111_LC_22_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i111_LC_22_15_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i111_LC_22_15_5  (
            .in0(N__66177),
            .in1(N__68923),
            .in2(N__51129),
            .in3(N__71948),
            .lcout(\c0.data_in_frame_13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71162),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i166_LC_22_15_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i166_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i166_LC_22_15_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i166_LC_22_15_6  (
            .in0(N__67945),
            .in1(N__67131),
            .in2(N__71806),
            .in3(N__72424),
            .lcout(\c0.data_in_frame_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71162),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i110_LC_22_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i110_LC_22_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i110_LC_22_15_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i110_LC_22_15_7  (
            .in0(N__51707),
            .in1(N__67946),
            .in2(N__66203),
            .in3(N__71947),
            .lcout(\c0.data_in_frame_13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71162),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_401_LC_22_16_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_401_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_401_LC_22_16_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_401_LC_22_16_0  (
            .in0(N__65406),
            .in1(N__51514),
            .in2(N__64821),
            .in3(N__51688),
            .lcout(),
            .ltout(\c0.n43_adj_3232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_22_16_1 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_22_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_LC_22_16_1  (
            .in0(N__51553),
            .in1(N__51649),
            .in2(N__51640),
            .in3(N__51601),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_3_lut_LC_22_16_2 .C_ON=1'b0;
    defparam \c0.i21_3_lut_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_3_lut_LC_22_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i21_3_lut_LC_22_16_2  (
            .in0(N__58404),
            .in1(N__51636),
            .in2(_gnd_net_),
            .in3(N__52015),
            .lcout(\c0.n49_adj_3237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_903_LC_22_16_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_903_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_903_LC_22_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_903_LC_22_16_3  (
            .in0(N__60843),
            .in1(N__62497),
            .in2(N__55959),
            .in3(N__60791),
            .lcout(\c0.n7_adj_3225 ),
            .ltout(\c0.n7_adj_3225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_666_LC_22_16_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_666_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_666_LC_22_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_666_LC_22_16_4  (
            .in0(N__56560),
            .in1(N__51588),
            .in2(N__51595),
            .in3(N__62307),
            .lcout(\c0.n11590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_395_LC_22_16_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_395_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_395_LC_22_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_395_LC_22_16_5  (
            .in0(N__62308),
            .in1(N__64703),
            .in2(N__51592),
            .in3(N__51559),
            .lcout(\c0.n44_adj_3226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_750_LC_22_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_750_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_750_LC_22_16_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_750_LC_22_16_6  (
            .in0(_gnd_net_),
            .in1(N__65680),
            .in2(_gnd_net_),
            .in3(N__65795),
            .lcout(\c0.n19202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_3_lut_adj_872_LC_22_17_0 .C_ON=1'b0;
    defparam \c0.i8_2_lut_3_lut_adj_872_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_3_lut_adj_872_LC_22_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i8_2_lut_3_lut_adj_872_LC_22_17_0  (
            .in0(N__51544),
            .in1(N__58462),
            .in2(_gnd_net_),
            .in3(N__51513),
            .lcout(\c0.n41_adj_3365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_3_lut_4_lut_LC_22_17_1 .C_ON=1'b0;
    defparam \c0.i19_3_lut_4_lut_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i19_3_lut_4_lut_LC_22_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_3_lut_4_lut_LC_22_17_1  (
            .in0(N__63630),
            .in1(N__51730),
            .in2(N__63688),
            .in3(N__52166),
            .lcout(),
            .ltout(\c0.n47_adj_3286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_450_LC_22_17_2 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_450_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_450_LC_22_17_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i24_4_lut_adj_450_LC_22_17_2  (
            .in0(N__67673),
            .in1(N__51892),
            .in2(N__51874),
            .in3(N__58068),
            .lcout(),
            .ltout(\c0.n52_adj_3288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_452_LC_22_17_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_452_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_452_LC_22_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_452_LC_22_17_3  (
            .in0(N__51871),
            .in1(N__65452),
            .in2(N__51865),
            .in3(N__57760),
            .lcout(\c0.n6_adj_3291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i95_LC_22_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i95_LC_22_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i95_LC_22_17_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i95_LC_22_17_4  (
            .in0(N__64542),
            .in1(N__51833),
            .in2(N__66205),
            .in3(N__69011),
            .lcout(\c0.data_in_frame_11_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71116),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_22_17_5 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_22_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_22_17_5  (
            .in0(N__63574),
            .in1(N__63495),
            .in2(_gnd_net_),
            .in3(N__51775),
            .lcout(\c0.n19909 ),
            .ltout(\c0.n19909_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i36_3_lut_4_lut_LC_22_17_6 .C_ON=1'b0;
    defparam \c0.i36_3_lut_4_lut_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i36_3_lut_4_lut_LC_22_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i36_3_lut_4_lut_LC_22_17_6  (
            .in0(N__63628),
            .in1(N__63683),
            .in2(N__51811),
            .in3(N__58067),
            .lcout(\c0.n87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_3_lut_adj_648_LC_22_17_7 .C_ON=1'b0;
    defparam \c0.i15_2_lut_3_lut_adj_648_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_3_lut_adj_648_LC_22_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i15_2_lut_3_lut_adj_648_LC_22_17_7  (
            .in0(N__63629),
            .in1(N__63496),
            .in2(_gnd_net_),
            .in3(N__51776),
            .lcout(\c0.n35_adj_3098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_adj_309_LC_22_18_0 .C_ON=1'b0;
    defparam \c0.i28_4_lut_adj_309_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_adj_309_LC_22_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i28_4_lut_adj_309_LC_22_18_0  (
            .in0(N__52543),
            .in1(N__59010),
            .in2(N__57820),
            .in3(N__53506),
            .lcout(\c0.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_2_lut_3_lut_LC_22_18_2 .C_ON=1'b0;
    defparam \c0.i12_2_lut_3_lut_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_2_lut_3_lut_LC_22_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i12_2_lut_3_lut_LC_22_18_2  (
            .in0(N__63776),
            .in1(N__65519),
            .in2(_gnd_net_),
            .in3(N__51729),
            .lcout(\c0.n45_adj_3423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_340_LC_22_18_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_340_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_340_LC_22_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_340_LC_22_18_3  (
            .in0(_gnd_net_),
            .in1(N__65796),
            .in2(_gnd_net_),
            .in3(N__53943),
            .lcout(\c0.n7_adj_3047 ),
            .ltout(\c0.n7_adj_3047_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_344_LC_22_18_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_344_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_344_LC_22_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_344_LC_22_18_4  (
            .in0(N__52231),
            .in1(N__52216),
            .in2(N__52195),
            .in3(N__59358),
            .lcout(\c0.n7_adj_3079 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_adj_603_LC_22_18_5 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_adj_603_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_adj_603_LC_22_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_2_lut_3_lut_adj_603_LC_22_18_5  (
            .in0(N__64057),
            .in1(N__57501),
            .in2(_gnd_net_),
            .in3(N__63485),
            .lcout(\c0.n28_adj_3059 ),
            .ltout(\c0.n28_adj_3059_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_3_lut_LC_22_18_6 .C_ON=1'b0;
    defparam \c0.i14_2_lut_3_lut_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_3_lut_LC_22_18_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i14_2_lut_3_lut_LC_22_18_6  (
            .in0(N__63627),
            .in1(_gnd_net_),
            .in2(N__52192),
            .in3(N__63560),
            .lcout(\c0.n33_adj_3315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_3_lut_4_lut_LC_22_18_7 .C_ON=1'b0;
    defparam \c0.i13_2_lut_3_lut_4_lut_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_3_lut_4_lut_LC_22_18_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_2_lut_3_lut_4_lut_LC_22_18_7  (
            .in0(N__63775),
            .in1(N__52189),
            .in2(N__65526),
            .in3(N__52167),
            .lcout(\c0.n32_adj_3465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_4_lut_LC_22_19_0 .C_ON=1'b0;
    defparam \c0.i10_3_lut_4_lut_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_4_lut_LC_22_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_3_lut_4_lut_LC_22_19_0  (
            .in0(N__52135),
            .in1(N__52108),
            .in2(N__55675),
            .in3(N__52060),
            .lcout(),
            .ltout(\c0.n29_adj_3461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_625_LC_22_19_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_625_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_625_LC_22_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_625_LC_22_19_1  (
            .in0(N__52249),
            .in1(N__52054),
            .in2(N__52024),
            .in3(N__52021),
            .lcout(),
            .ltout(\c0.n36_adj_3470_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_626_LC_22_19_2 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_626_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_626_LC_22_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_626_LC_22_19_2  (
            .in0(N__51973),
            .in1(N__51946),
            .in2(N__51919),
            .in3(N__51916),
            .lcout(\c0.n11_adj_3124 ),
            .ltout(\c0.n11_adj_3124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_629_LC_22_19_3 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_629_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_629_LC_22_19_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i4_2_lut_adj_629_LC_22_19_3  (
            .in0(N__53804),
            .in1(_gnd_net_),
            .in2(N__51895),
            .in3(_gnd_net_),
            .lcout(\c0.n37_adj_3268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_2_lut_LC_22_19_4 .C_ON=1'b0;
    defparam \c0.i27_2_lut_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i27_2_lut_LC_22_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i27_2_lut_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__52397),
            .in2(_gnd_net_),
            .in3(N__52405),
            .lcout(\c0.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_339_LC_22_19_5 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_339_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_339_LC_22_19_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_adj_339_LC_22_19_5  (
            .in0(_gnd_net_),
            .in1(N__58840),
            .in2(_gnd_net_),
            .in3(N__57952),
            .lcout(\c0.n42_adj_3086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_adj_471_LC_22_19_6 .C_ON=1'b0;
    defparam \c0.i26_4_lut_adj_471_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_adj_471_LC_22_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_adj_471_LC_22_19_6  (
            .in0(N__52398),
            .in1(N__52378),
            .in2(N__57940),
            .in3(N__52366),
            .lcout(\c0.n19764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_890_LC_22_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_890_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_890_LC_22_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_890_LC_22_20_0  (
            .in0(N__69965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72832),
            .lcout(\c0.n11971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_22_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_22_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_664_LC_22_20_1  (
            .in0(N__72833),
            .in1(N__69966),
            .in2(_gnd_net_),
            .in3(N__69636),
            .lcout(\c0.n18379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_683_LC_22_20_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_683_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_683_LC_22_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_683_LC_22_20_2  (
            .in0(N__52350),
            .in1(N__67404),
            .in2(N__68392),
            .in3(N__52282),
            .lcout(\c0.n22_adj_3363 ),
            .ltout(\c0.n22_adj_3363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_623_LC_22_20_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_623_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_623_LC_22_20_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i11_3_lut_adj_623_LC_22_20_3  (
            .in0(N__69496),
            .in1(_gnd_net_),
            .in2(N__52252),
            .in3(N__69964),
            .lcout(\c0.n30_adj_3468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_513_LC_22_20_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_513_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_513_LC_22_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_513_LC_22_20_4  (
            .in0(N__68300),
            .in1(N__68428),
            .in2(N__68391),
            .in3(N__69818),
            .lcout(\c0.n6009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i33_4_lut_LC_22_20_5 .C_ON=1'b0;
    defparam \c0.i33_4_lut_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i33_4_lut_LC_22_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i33_4_lut_LC_22_20_5  (
            .in0(N__57883),
            .in1(N__52240),
            .in2(N__57909),
            .in3(N__52416),
            .lcout(),
            .ltout(\c0.n70_adj_3087_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i36_4_lut_LC_22_20_6 .C_ON=1'b0;
    defparam \c0.i36_4_lut_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i36_4_lut_LC_22_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i36_4_lut_LC_22_20_6  (
            .in0(N__57838),
            .in1(N__58612),
            .in2(N__52693),
            .in3(N__57928),
            .lcout(\c0.n20339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_655_LC_22_20_7 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_655_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_655_LC_22_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_655_LC_22_20_7  (
            .in0(N__72834),
            .in1(N__69967),
            .in2(_gnd_net_),
            .in3(N__53459),
            .lcout(\c0.n27_adj_3311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_455_LC_22_21_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_455_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_455_LC_22_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_455_LC_22_21_0  (
            .in0(N__52645),
            .in1(N__52615),
            .in2(N__66694),
            .in3(N__52606),
            .lcout(),
            .ltout(\c0.n32_adj_3294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_459_LC_22_21_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_459_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_459_LC_22_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_459_LC_22_21_1  (
            .in0(N__53443),
            .in1(N__52588),
            .in2(N__52582),
            .in3(N__52525),
            .lcout(\c0.n21075 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_4_lut_LC_22_21_2 .C_ON=1'b0;
    defparam \c0.i11_3_lut_4_lut_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_4_lut_LC_22_21_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i11_3_lut_4_lut_LC_22_21_2  (
            .in0(N__52708),
            .in1(N__52559),
            .in2(N__52489),
            .in3(N__57857),
            .lcout(\c0.n29_adj_3299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i172_LC_22_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i172_LC_22_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i172_LC_22_21_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i172_LC_22_21_3  (
            .in0(N__71778),
            .in1(N__71977),
            .in2(N__69602),
            .in3(N__69287),
            .lcout(\c0.data_in_frame_21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71185),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_473_LC_22_21_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_473_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_473_LC_22_21_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_473_LC_22_21_4  (
            .in0(N__52507),
            .in1(N__52707),
            .in2(N__52490),
            .in3(N__57858),
            .lcout(\c0.n19_adj_3320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_4_lut_adj_783_LC_22_21_5 .C_ON=1'b0;
    defparam \c0.i20_3_lut_4_lut_adj_783_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_4_lut_adj_783_LC_22_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_3_lut_4_lut_adj_783_LC_22_21_5  (
            .in0(N__52706),
            .in1(N__52506),
            .in2(N__52492),
            .in3(N__52445),
            .lcout(\c0.n57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_584_LC_22_21_6 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_584_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_584_LC_22_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_584_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__52875),
            .in2(_gnd_net_),
            .in3(N__59032),
            .lcout(\c0.n39_adj_3384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_695_LC_22_22_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_695_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_695_LC_22_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_695_LC_22_22_0  (
            .in0(N__53342),
            .in1(N__53391),
            .in2(N__68125),
            .in3(N__53298),
            .lcout(\c0.n11714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_457_LC_22_22_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_457_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_457_LC_22_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_457_LC_22_22_1  (
            .in0(N__52735),
            .in1(N__68124),
            .in2(N__53395),
            .in3(N__53343),
            .lcout(\c0.n22_adj_3296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_321_LC_22_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_321_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_321_LC_22_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_321_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(N__68236),
            .in2(_gnd_net_),
            .in3(N__53297),
            .lcout(\c0.n19159 ),
            .ltout(\c0.n19159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_749_LC_22_22_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_749_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_749_LC_22_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_749_LC_22_22_3  (
            .in0(N__53808),
            .in1(N__72438),
            .in2(N__52831),
            .in3(N__52828),
            .lcout(\c0.n12206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_adj_504_LC_22_22_4 .C_ON=1'b0;
    defparam \c0.i30_4_lut_adj_504_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_adj_504_LC_22_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i30_4_lut_adj_504_LC_22_22_4  (
            .in0(N__52804),
            .in1(N__53353),
            .in2(N__52798),
            .in3(N__53585),
            .lcout(\c0.n79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_373_LC_22_22_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_373_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_373_LC_22_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_373_LC_22_22_5  (
            .in0(N__58041),
            .in1(N__58794),
            .in2(_gnd_net_),
            .in3(N__53421),
            .lcout(\c0.n19151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_364_LC_22_22_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_364_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_364_LC_22_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_364_LC_22_22_6  (
            .in0(N__52762),
            .in1(N__59011),
            .in2(N__57256),
            .in3(N__52734),
            .lcout(\c0.n11776 ),
            .ltout(\c0.n11776_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_561_LC_22_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_561_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_561_LC_22_22_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_561_LC_22_22_7  (
            .in0(N__68235),
            .in1(N__72437),
            .in2(N__52711),
            .in3(N__59504),
            .lcout(\c0.n6_adj_3319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_317_LC_22_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_317_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_317_LC_22_23_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_317_LC_22_23_0  (
            .in0(N__53626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53601),
            .lcout(\c0.n19268 ),
            .ltout(\c0.n19268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_649_LC_22_23_1 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_649_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_649_LC_22_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_649_LC_22_23_1  (
            .in0(N__53511),
            .in1(N__66647),
            .in2(N__53563),
            .in3(N__53539),
            .lcout(\c0.n20_adj_3301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_22_23_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_22_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_22_23_2  (
            .in0(N__53538),
            .in1(N__53510),
            .in2(N__66649),
            .in3(N__53469),
            .lcout(\c0.n42_adj_3055 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_323_LC_22_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_323_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_323_LC_22_23_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_323_LC_22_23_3  (
            .in0(N__67697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53425),
            .lcout(\c0.n4_adj_3100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_375_LC_22_23_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_375_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_375_LC_22_23_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_375_LC_22_23_4  (
            .in0(N__53272),
            .in1(N__53375),
            .in2(N__58114),
            .in3(N__64632),
            .lcout(\c0.n19436 ),
            .ltout(\c0.n19436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_adj_697_LC_22_23_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_adj_697_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_adj_697_LC_22_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_adj_697_LC_22_23_5  (
            .in0(N__53344),
            .in1(N__68119),
            .in2(N__53302),
            .in3(N__53299),
            .lcout(\c0.n6_adj_3112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_336_LC_22_23_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_336_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_336_LC_22_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_336_LC_22_23_6  (
            .in0(N__53271),
            .in1(N__69787),
            .in2(N__58849),
            .in3(N__67696),
            .lcout(\c0.n20933 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6__5175_LC_22_23_7 .C_ON=1'b0;
    defparam \c0.data_in_2__6__5175_LC_22_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6__5175_LC_22_23_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__6__5175_LC_22_23_7  (
            .in0(N__53135),
            .in1(N__52960),
            .in2(_gnd_net_),
            .in3(N__52903),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71207),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_LC_22_24_0 .C_ON=1'b0;
    defparam \c0.i7_3_lut_LC_22_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_LC_22_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_3_lut_LC_22_24_0  (
            .in0(N__59274),
            .in1(N__59230),
            .in2(_gnd_net_),
            .in3(N__59828),
            .lcout(\c0.n25_adj_3048 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_377_LC_22_24_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_377_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_377_LC_22_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_377_LC_22_24_1  (
            .in0(N__72392),
            .in1(N__53973),
            .in2(N__69606),
            .in3(N__53947),
            .lcout(),
            .ltout(\c0.n12_adj_3210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_378_LC_22_24_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_378_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_378_LC_22_24_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_378_LC_22_24_2  (
            .in0(N__53911),
            .in1(N__66453),
            .in2(N__53884),
            .in3(N__53881),
            .lcout(\c0.n17834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_109_2_lut_LC_22_24_3 .C_ON=1'b0;
    defparam \c0.i1_rep_109_2_lut_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_109_2_lut_LC_22_24_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_rep_109_2_lut_LC_22_24_3  (
            .in0(N__59231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59275),
            .lcout(\c0.n21767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_338_LC_22_24_4 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_338_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_338_LC_22_24_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i4_2_lut_adj_338_LC_22_24_4  (
            .in0(N__53809),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53770),
            .lcout(\c0.n41_adj_3085 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i189_LC_22_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i189_LC_22_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i189_LC_22_24_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i189_LC_22_24_5  (
            .in0(N__72733),
            .in1(N__53709),
            .in2(_gnd_net_),
            .in3(N__53744),
            .lcout(data_in_frame_23_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71219),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i190_LC_22_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i190_LC_22_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i190_LC_22_24_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i190_LC_22_24_6  (
            .in0(N__53710),
            .in1(N__67980),
            .in2(_gnd_net_),
            .in3(N__66454),
            .lcout(data_in_frame_23_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71219),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_67_i9_2_lut_3_lut_LC_23_7_0 .C_ON=1'b0;
    defparam \c0.equal_67_i9_2_lut_3_lut_LC_23_7_0 .SEQ_MODE=4'b0000;
    defparam \c0.equal_67_i9_2_lut_3_lut_LC_23_7_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.equal_67_i9_2_lut_3_lut_LC_23_7_0  (
            .in0(N__60268),
            .in1(N__59996),
            .in2(_gnd_net_),
            .in3(N__60117),
            .lcout(\c0.n9_adj_3211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_4_lut_LC_23_8_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_4_lut_LC_23_8_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_4_lut_LC_23_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_4_lut_LC_23_8_0  (
            .in0(N__54211),
            .in1(N__54187),
            .in2(N__53662),
            .in3(N__54579),
            .lcout(\c0.n7_adj_3347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_812_LC_23_8_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_812_LC_23_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_812_LC_23_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i13_4_lut_adj_812_LC_23_8_2  (
            .in0(N__54680),
            .in1(N__55377),
            .in2(N__54628),
            .in3(N__60922),
            .lcout(\c0.n34_adj_3326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_adj_912_LC_23_8_3 .C_ON=1'b0;
    defparam \c0.i7_3_lut_adj_912_LC_23_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_adj_912_LC_23_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i7_3_lut_adj_912_LC_23_8_3  (
            .in0(N__54186),
            .in1(_gnd_net_),
            .in2(N__54580),
            .in3(N__54210),
            .lcout(\c0.n11982 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_719_LC_23_8_4 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_719_LC_23_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_719_LC_23_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_719_LC_23_8_4  (
            .in0(N__54568),
            .in1(N__54530),
            .in2(N__54502),
            .in3(N__54480),
            .lcout(\c0.n58_adj_3497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_771_LC_23_8_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_771_LC_23_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_771_LC_23_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_771_LC_23_8_5  (
            .in0(_gnd_net_),
            .in1(N__54315),
            .in2(_gnd_net_),
            .in3(N__54271),
            .lcout(\c0.n8_adj_3345 ),
            .ltout(\c0.n8_adj_3345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_779_LC_23_8_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_779_LC_23_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_779_LC_23_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_779_LC_23_8_6  (
            .in0(N__54198),
            .in1(N__54185),
            .in2(N__54172),
            .in3(N__56398),
            .lcout(\c0.n11626 ),
            .ltout(\c0.n11626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_372_LC_23_8_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_372_LC_23_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_372_LC_23_8_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_372_LC_23_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54169),
            .in3(N__54166),
            .lcout(\c0.n12209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_519_LC_23_9_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_519_LC_23_9_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_519_LC_23_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_519_LC_23_9_0  (
            .in0(N__54634),
            .in1(N__54115),
            .in2(N__54858),
            .in3(N__55277),
            .lcout(\c0.n19970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_728_LC_23_9_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_728_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_728_LC_23_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_728_LC_23_9_1  (
            .in0(N__54031),
            .in1(N__54834),
            .in2(N__54020),
            .in3(N__54672),
            .lcout(\c0.n11478 ),
            .ltout(\c0.n11478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_4_lut_LC_23_9_2 .C_ON=1'b0;
    defparam \c0.i29_4_lut_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.i29_4_lut_LC_23_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i29_4_lut_LC_23_9_2  (
            .in0(N__56630),
            .in1(N__54781),
            .in2(N__54904),
            .in3(N__54731),
            .lcout(\c0.n81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_23_9_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_23_9_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_23_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i15_LC_23_9_3  (
            .in0(N__68866),
            .in1(N__59884),
            .in2(_gnd_net_),
            .in3(N__54835),
            .lcout(data_in_frame_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71231),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_835_LC_23_9_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_835_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_835_LC_23_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_835_LC_23_9_4  (
            .in0(_gnd_net_),
            .in1(N__60907),
            .in2(_gnd_net_),
            .in3(N__62624),
            .lcout(\c0.n11526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_23_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_23_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_23_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i54_LC_23_9_5  (
            .in0(N__62030),
            .in1(N__61615),
            .in2(N__54775),
            .in3(N__67912),
            .lcout(\c0.data_in_frame_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71231),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_606_LC_23_9_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_606_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_606_LC_23_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_606_LC_23_9_6  (
            .in0(N__56938),
            .in1(N__57043),
            .in2(N__54757),
            .in3(N__54732),
            .lcout(\c0.n27_adj_3457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_805_LC_23_9_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_805_LC_23_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_805_LC_23_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_adj_805_LC_23_9_7  (
            .in0(_gnd_net_),
            .in1(N__61193),
            .in2(_gnd_net_),
            .in3(N__54671),
            .lcout(\c0.n12_adj_3378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_23_10_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_23_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_23_10_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i48_LC_23_10_0  (
            .in0(N__61757),
            .in1(N__60352),
            .in2(N__62681),
            .in3(N__72149),
            .lcout(\c0.data_in_frame_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71227),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_23_10_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_23_10_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_23_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i13_LC_23_10_1  (
            .in0(N__59866),
            .in1(N__72613),
            .in2(_gnd_net_),
            .in3(N__60916),
            .lcout(data_in_frame_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71227),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_23_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_23_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i14_LC_23_10_2  (
            .in0(N__67911),
            .in1(N__59867),
            .in2(_gnd_net_),
            .in3(N__55345),
            .lcout(data_in_frame_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71227),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_564_LC_23_10_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_564_LC_23_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_564_LC_23_10_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i11_3_lut_adj_564_LC_23_10_3  (
            .in0(N__55420),
            .in1(N__55411),
            .in2(_gnd_net_),
            .in3(N__60842),
            .lcout(\c0.n28_adj_3428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_800_LC_23_10_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_800_LC_23_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_800_LC_23_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_800_LC_23_10_4  (
            .in0(N__60388),
            .in1(N__60899),
            .in2(_gnd_net_),
            .in3(N__55344),
            .lcout(\c0.n7_adj_3509 ),
            .ltout(\c0.n7_adj_3509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_803_LC_23_10_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_803_LC_23_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_803_LC_23_10_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_803_LC_23_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55294),
            .in3(N__55010),
            .lcout(\c0.n10_adj_3012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_23_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_23_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_23_10_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.data_in_frame_0__i9_LC_23_10_6  (
            .in0(_gnd_net_),
            .in1(N__65259),
            .in2(N__55031),
            .in3(N__59868),
            .lcout(data_in_frame_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71227),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_4_lut_adj_862_LC_23_10_7 .C_ON=1'b0;
    defparam \c0.i23_3_lut_4_lut_adj_862_LC_23_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_4_lut_adj_862_LC_23_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_3_lut_4_lut_adj_862_LC_23_10_7  (
            .in0(N__62409),
            .in1(N__55264),
            .in2(N__62464),
            .in3(N__55240),
            .lcout(\c0.n56_adj_3505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_709_LC_23_11_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_709_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_709_LC_23_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_709_LC_23_11_0  (
            .in0(N__55108),
            .in1(N__55014),
            .in2(_gnd_net_),
            .in3(N__60389),
            .lcout(\c0.n20341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_4_lut_adj_731_LC_23_11_1 .C_ON=1'b0;
    defparam \c0.i31_4_lut_adj_731_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.i31_4_lut_adj_731_LC_23_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i31_4_lut_adj_731_LC_23_11_1  (
            .in0(N__54910),
            .in1(N__54952),
            .in2(N__61141),
            .in3(N__54943),
            .lcout(\c0.n64_adj_3506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_838_LC_23_11_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_838_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_838_LC_23_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_838_LC_23_11_2  (
            .in0(_gnd_net_),
            .in1(N__61326),
            .in2(_gnd_net_),
            .in3(N__60390),
            .lcout(\c0.n4_adj_3036 ),
            .ltout(\c0.n4_adj_3036_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_723_LC_23_11_3 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_723_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_723_LC_23_11_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_adj_723_LC_23_11_3  (
            .in0(N__62353),
            .in1(N__54925),
            .in2(N__54913),
            .in3(N__62619),
            .lcout(\c0.n57_adj_3499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_899_LC_23_11_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_899_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_899_LC_23_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_899_LC_23_11_4  (
            .in0(N__62618),
            .in1(N__61327),
            .in2(_gnd_net_),
            .in3(N__60391),
            .lcout(\c0.n6_adj_3019 ),
            .ltout(\c0.n6_adj_3019_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_244_LC_23_11_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_244_LC_23_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_244_LC_23_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_244_LC_23_11_5  (
            .in0(N__62320),
            .in1(N__55704),
            .in2(N__55678),
            .in3(N__60909),
            .lcout(\c0.n20386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i79_LC_23_11_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i79_LC_23_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i79_LC_23_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i79_LC_23_11_6  (
            .in0(N__66145),
            .in1(N__63418),
            .in2(N__55614),
            .in3(N__68826),
            .lcout(\c0.data_in_frame_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71220),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i64_LC_23_12_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i64_LC_23_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i64_LC_23_12_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i64_LC_23_12_0  (
            .in0(N__64409),
            .in1(N__61756),
            .in2(N__62410),
            .in3(N__72132),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_23_12_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_23_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_23_12_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i32_LC_23_12_1  (
            .in0(N__61752),
            .in1(N__61455),
            .in2(N__72201),
            .in3(N__55583),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_23_12_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_23_12_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_23_12_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i30_LC_23_12_2  (
            .in0(N__61454),
            .in1(N__61754),
            .in2(N__62626),
            .in3(N__67952),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_23_12_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_23_12_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_23_12_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i46_LC_23_12_3  (
            .in0(N__61753),
            .in1(N__67951),
            .in2(N__60358),
            .in3(N__55540),
            .lcout(\c0.data_in_frame_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_23_12_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_23_12_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_23_12_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i44_LC_23_12_4  (
            .in0(N__69442),
            .in1(N__61755),
            .in2(N__55515),
            .in3(N__60354),
            .lcout(\c0.data_in_frame_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_23_12_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_23_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_23_12_5 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_23_12_5  (
            .in0(N__72128),
            .in1(N__56266),
            .in2(N__56226),
            .in3(N__55468),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_3_lut_4_lut_LC_23_12_6 .C_ON=1'b0;
    defparam \c0.i18_3_lut_4_lut_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i18_3_lut_4_lut_LC_23_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_3_lut_4_lut_LC_23_12_6  (
            .in0(N__60487),
            .in1(N__60448),
            .in2(N__62496),
            .in3(N__56295),
            .lcout(\c0.n51_adj_3426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_12_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_23_12_7 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_23_12_7  (
            .in0(N__56259),
            .in1(N__68853),
            .in2(N__56225),
            .in3(N__56085),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71208),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_823_LC_23_13_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_823_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_823_LC_23_13_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_823_LC_23_13_0  (
            .in0(N__64438),
            .in1(N__56028),
            .in2(N__57500),
            .in3(N__61873),
            .lcout(\c0.n13_adj_3541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i102_LC_23_13_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i102_LC_23_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i102_LC_23_13_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i102_LC_23_13_1  (
            .in0(N__67949),
            .in1(N__67220),
            .in2(N__66189),
            .in3(N__57632),
            .lcout(\c0.data_in_frame_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i107_LC_23_13_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i107_LC_23_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i107_LC_23_13_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i107_LC_23_13_2  (
            .in0(N__68725),
            .in1(N__71972),
            .in2(N__55951),
            .in3(N__66162),
            .lcout(\c0.data_in_frame_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i78_LC_23_13_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i78_LC_23_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i78_LC_23_13_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i78_LC_23_13_3  (
            .in0(N__67950),
            .in1(N__66193),
            .in2(N__55920),
            .in3(N__63380),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i65_LC_23_13_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i65_LC_23_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i65_LC_23_13_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i65_LC_23_13_4  (
            .in0(N__65230),
            .in1(N__62447),
            .in2(N__64249),
            .in3(N__55812),
            .lcout(\c0.data_in_frame_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i97_LC_23_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i97_LC_23_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i97_LC_23_13_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i97_LC_23_13_5  (
            .in0(N__66157),
            .in1(N__67221),
            .in2(N__57195),
            .in3(N__65234),
            .lcout(\c0.data_in_frame_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i73_LC_23_13_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i73_LC_23_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i73_LC_23_13_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i73_LC_23_13_6  (
            .in0(N__63379),
            .in1(N__66158),
            .in2(N__65258),
            .in3(N__63104),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71196),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_LC_23_13_7 .C_ON=1'b0;
    defparam \c0.i6_3_lut_LC_23_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_LC_23_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_3_lut_LC_23_13_7  (
            .in0(N__62250),
            .in1(N__56410),
            .in2(_gnd_net_),
            .in3(N__56847),
            .lcout(\c0.n17_adj_3544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_359_LC_23_14_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_359_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_359_LC_23_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_359_LC_23_14_0  (
            .in0(N__56939),
            .in1(N__57103),
            .in2(_gnd_net_),
            .in3(N__57044),
            .lcout(),
            .ltout(\c0.n11858_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_371_LC_23_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_371_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_371_LC_23_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_371_LC_23_14_1  (
            .in0(_gnd_net_),
            .in1(N__56727),
            .in2(N__56671),
            .in3(N__61871),
            .lcout(\c0.n19446 ),
            .ltout(\c0.n19446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_376_LC_23_14_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_376_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_376_LC_23_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_376_LC_23_14_2  (
            .in0(_gnd_net_),
            .in1(N__62904),
            .in2(N__56656),
            .in3(N__56653),
            .lcout(\c0.n33_adj_3209 ),
            .ltout(\c0.n33_adj_3209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_adj_827_LC_23_14_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_827_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_827_LC_23_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i3_3_lut_adj_827_LC_23_14_3  (
            .in0(_gnd_net_),
            .in1(N__56578),
            .in2(N__56569),
            .in3(N__56440),
            .lcout(\c0.n5598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_809_LC_23_14_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_809_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_809_LC_23_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_809_LC_23_14_4  (
            .in0(N__61872),
            .in1(N__56529),
            .in2(N__65433),
            .in3(N__56488),
            .lcout(\c0.n29_adj_3533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_3_lut_LC_23_14_5 .C_ON=1'b0;
    defparam \c0.i17_3_lut_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i17_3_lut_LC_23_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i17_3_lut_LC_23_14_5  (
            .in0(N__56458),
            .in1(N__56441),
            .in2(_gnd_net_),
            .in3(N__56409),
            .lcout(\c0.n45_adj_3224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_23_14_6 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_23_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i5_2_lut_LC_23_14_6  (
            .in0(_gnd_net_),
            .in1(N__56341),
            .in2(_gnd_net_),
            .in3(N__62679),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_391_LC_23_15_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_391_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_391_LC_23_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_391_LC_23_15_0  (
            .in0(N__57401),
            .in1(N__57271),
            .in2(N__57251),
            .in3(N__57187),
            .lcout(\c0.n19430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_917_LC_23_15_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_917_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_917_LC_23_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i6_2_lut_adj_917_LC_23_15_1  (
            .in0(_gnd_net_),
            .in1(N__62720),
            .in2(_gnd_net_),
            .in3(N__57157),
            .lcout(\c0.n20_adj_3536 ),
            .ltout(\c0.n20_adj_3536_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_918_LC_23_15_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_918_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_918_LC_23_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_918_LC_23_15_2  (
            .in0(_gnd_net_),
            .in1(N__56917),
            .in2(N__57121),
            .in3(N__58598),
            .lcout(),
            .ltout(\c0.n12_adj_3558_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_919_LC_23_15_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_919_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_919_LC_23_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_919_LC_23_15_3  (
            .in0(N__66354),
            .in1(N__60745),
            .in2(N__57118),
            .in3(N__58461),
            .lcout(\c0.n18420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_906_LC_23_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_906_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_906_LC_23_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_906_LC_23_15_4  (
            .in0(N__57115),
            .in1(N__56940),
            .in2(N__57076),
            .in3(N__57046),
            .lcout(\c0.n19359 ),
            .ltout(\c0.n19359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_392_LC_23_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_392_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_392_LC_23_15_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_392_LC_23_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56974),
            .in3(N__56902),
            .lcout(\c0.n19502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_914_LC_23_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_914_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_914_LC_23_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_914_LC_23_15_6  (
            .in0(_gnd_net_),
            .in1(N__56970),
            .in2(_gnd_net_),
            .in3(N__56941),
            .lcout(\c0.n19199 ),
            .ltout(\c0.n19199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_820_LC_23_15_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_820_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_820_LC_23_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_820_LC_23_15_7  (
            .in0(N__59530),
            .in1(N__56903),
            .in2(N__56881),
            .in3(N__66294),
            .lcout(\c0.n19_adj_3540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i142_LC_23_16_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i142_LC_23_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i142_LC_23_16_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i142_LC_23_16_0  (
            .in0(N__63416),
            .in1(N__67981),
            .in2(N__65326),
            .in3(N__71802),
            .lcout(\c0.data_in_frame_17_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i122_LC_23_16_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i122_LC_23_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i122_LC_23_16_1 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i122_LC_23_16_1  (
            .in0(N__71488),
            .in1(N__64254),
            .in2(N__64389),
            .in3(N__64979),
            .lcout(\c0.data_in_frame_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i208_LC_23_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i208_LC_23_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i208_LC_23_16_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i208_LC_23_16_2  (
            .in0(N__63417),
            .in1(N__66898),
            .in2(N__59783),
            .in3(N__72206),
            .lcout(\c0.data_in_frame_25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i114_LC_23_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i114_LC_23_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i114_LC_23_16_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i114_LC_23_16_3  (
            .in0(N__71487),
            .in1(N__64252),
            .in2(N__57499),
            .in3(N__62058),
            .lcout(\c0.data_in_frame_14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i128_LC_23_16_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i128_LC_23_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i128_LC_23_16_4 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i128_LC_23_16_4  (
            .in0(N__64251),
            .in1(N__64362),
            .in2(N__57434),
            .in3(N__72205),
            .lcout(\c0.data_in_frame_15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i115_LC_23_16_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i115_LC_23_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i115_LC_23_16_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i115_LC_23_16_5  (
            .in0(N__68722),
            .in1(N__64253),
            .in2(N__57408),
            .in3(N__62059),
            .lcout(\c0.data_in_frame_14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_23_16_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_23_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_23_16_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_in_frame_0__i59_LC_23_16_6  (
            .in0(N__57361),
            .in1(N__68723),
            .in2(N__61599),
            .in3(N__64366),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71163),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_360_LC_23_16_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_360_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_360_LC_23_16_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i8_4_lut_adj_360_LC_23_16_7  (
            .in0(N__62527),
            .in1(N__62680),
            .in2(N__62551),
            .in3(N__57331),
            .lcout(\c0.n25_adj_3157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_4_lut_adj_865_LC_23_17_0 .C_ON=1'b0;
    defparam \c0.i11_3_lut_4_lut_adj_865_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_4_lut_adj_865_LC_23_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_3_lut_4_lut_adj_865_LC_23_17_0  (
            .in0(N__69688),
            .in1(N__70083),
            .in2(N__58899),
            .in3(N__59009),
            .lcout(\c0.n32_adj_3060 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_290_LC_23_17_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_290_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_290_LC_23_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_290_LC_23_17_1  (
            .in0(N__59047),
            .in1(N__58667),
            .in2(N__70498),
            .in3(N__58629),
            .lcout(),
            .ltout(\c0.n38_adj_3058_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_23_17_2 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_23_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_23_17_2  (
            .in0(N__57837),
            .in1(N__57819),
            .in2(N__57802),
            .in3(N__57799),
            .lcout(\c0.n8_adj_3061 ),
            .ltout(\c0.n8_adj_3061_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_3_lut_LC_23_17_3 .C_ON=1'b0;
    defparam \c0.i19_3_lut_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i19_3_lut_LC_23_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i19_3_lut_LC_23_17_3  (
            .in0(_gnd_net_),
            .in1(N__70460),
            .in2(N__57793),
            .in3(N__59178),
            .lcout(\c0.n52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_449_LC_23_17_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_449_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_449_LC_23_17_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_449_LC_23_17_4  (
            .in0(N__70021),
            .in1(N__70242),
            .in2(N__70465),
            .in3(N__57769),
            .lcout(),
            .ltout(\c0.n43_adj_3285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_3_lut_4_lut_LC_23_17_5 .C_ON=1'b0;
    defparam \c0.i25_3_lut_4_lut_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i25_3_lut_4_lut_LC_23_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_3_lut_4_lut_LC_23_17_5  (
            .in0(N__58668),
            .in1(N__68023),
            .in2(N__57763),
            .in3(N__67303),
            .lcout(\c0.n53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_23_18_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_23_18_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i6_2_lut_LC_23_18_0  (
            .in0(N__67264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57754),
            .lcout(\c0.n43_adj_3089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_883_LC_23_18_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_883_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_883_LC_23_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_883_LC_23_18_1  (
            .in0(N__57736),
            .in1(N__67386),
            .in2(N__64831),
            .in3(N__57645),
            .lcout(),
            .ltout(\c0.n12_adj_3554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_884_LC_23_18_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_884_LC_23_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_884_LC_23_18_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_884_LC_23_18_2  (
            .in0(N__67438),
            .in1(N__67354),
            .in2(N__57589),
            .in3(N__57586),
            .lcout(\c0.n20542 ),
            .ltout(\c0.n20542_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_891_LC_23_18_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_891_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_891_LC_23_18_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_891_LC_23_18_3  (
            .in0(N__67613),
            .in1(N__58798),
            .in2(N__57535),
            .in3(N__67263),
            .lcout(\c0.n25_adj_3510 ),
            .ltout(\c0.n25_adj_3510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_737_LC_23_18_4 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_737_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_737_LC_23_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_adj_737_LC_23_18_4  (
            .in0(N__63647),
            .in1(N__57525),
            .in2(N__57514),
            .in3(N__66582),
            .lcout(\c0.n58_adj_3511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i37_3_lut_4_lut_LC_23_18_5 .C_ON=1'b0;
    defparam \c0.i37_3_lut_4_lut_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i37_3_lut_4_lut_LC_23_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i37_3_lut_4_lut_LC_23_18_5  (
            .in0(N__58072),
            .in1(N__67675),
            .in2(N__63652),
            .in3(N__58042),
            .lcout(\c0.n88_adj_3422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_adj_893_LC_23_18_6 .C_ON=1'b0;
    defparam \c0.i5_2_lut_adj_893_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_adj_893_LC_23_18_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i5_2_lut_adj_893_LC_23_18_6  (
            .in0(N__59779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57994),
            .lcout(\c0.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i29_3_lut_LC_23_19_0 .C_ON=1'b0;
    defparam \c0.i29_3_lut_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i29_3_lut_LC_23_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i29_3_lut_LC_23_19_0  (
            .in0(N__58336),
            .in1(N__58306),
            .in2(_gnd_net_),
            .in3(N__57973),
            .lcout(\c0.n60_adj_3127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_469_LC_23_19_1 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_469_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_469_LC_23_19_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i21_4_lut_adj_469_LC_23_19_1  (
            .in0(N__59004),
            .in1(N__58287),
            .in2(N__67270),
            .in3(N__57951),
            .lcout(\c0.n48_adj_3313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_824_LC_23_19_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_824_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_824_LC_23_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_824_LC_23_19_2  (
            .in0(N__68113),
            .in1(_gnd_net_),
            .in2(N__68228),
            .in3(N__58099),
            .lcout(),
            .ltout(\c0.n35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_LC_23_19_3 .C_ON=1'b0;
    defparam \c0.i30_4_lut_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_LC_23_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i30_4_lut_LC_23_19_3  (
            .in0(N__69919),
            .in1(N__69714),
            .in2(N__57931),
            .in3(N__57922),
            .lcout(\c0.n67_adj_3092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_341_LC_23_19_4 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_341_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_341_LC_23_19_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i24_4_lut_adj_341_LC_23_19_4  (
            .in0(N__57921),
            .in1(N__59005),
            .in2(N__57910),
            .in3(N__57882),
            .lcout(),
            .ltout(\c0.n55_adj_3128_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30_4_lut_adj_343_LC_23_19_5 .C_ON=1'b0;
    defparam \c0.i30_4_lut_adj_343_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30_4_lut_adj_343_LC_23_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i30_4_lut_adj_343_LC_23_19_5  (
            .in0(N__58288),
            .in1(N__57871),
            .in2(N__57865),
            .in3(N__67993),
            .lcout(\c0.n19749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_698_LC_23_19_6 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_698_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_698_LC_23_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i14_4_lut_adj_698_LC_23_19_6  (
            .in0(N__58335),
            .in1(N__59003),
            .in2(N__58327),
            .in3(N__58305),
            .lcout(\c0.n10_adj_3425 ),
            .ltout(\c0.n10_adj_3425_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_23_19_7 .C_ON=1'b0;
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_3_lut_4_lut_LC_23_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_2_lut_3_lut_4_lut_LC_23_19_7  (
            .in0(N__69918),
            .in1(N__68217),
            .in2(N__58291),
            .in3(N__68112),
            .lcout(\c0.n42_adj_3130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i41_4_lut_adj_437_LC_23_20_0 .C_ON=1'b0;
    defparam \c0.i41_4_lut_adj_437_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i41_4_lut_adj_437_LC_23_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i41_4_lut_adj_437_LC_23_20_0  (
            .in0(N__58264),
            .in1(N__67242),
            .in2(N__58228),
            .in3(N__58200),
            .lcout(\c0.n92_adj_3272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_adj_707_LC_23_20_1 .C_ON=1'b0;
    defparam \c0.i6_2_lut_adj_707_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_adj_707_LC_23_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i6_2_lut_adj_707_LC_23_20_1  (
            .in0(_gnd_net_),
            .in1(N__67266),
            .in2(_gnd_net_),
            .in3(N__58098),
            .lcout(\c0.n39_adj_3269 ),
            .ltout(\c0.n39_adj_3269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i41_4_lut_adj_518_LC_23_20_2 .C_ON=1'b0;
    defparam \c0.i41_4_lut_adj_518_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i41_4_lut_adj_518_LC_23_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i41_4_lut_adj_518_LC_23_20_2  (
            .in0(N__58258),
            .in1(N__58227),
            .in2(N__58204),
            .in3(N__58201),
            .lcout(),
            .ltout(\c0.n92_adj_3377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i49_4_lut_adj_557_LC_23_20_3 .C_ON=1'b0;
    defparam \c0.i49_4_lut_adj_557_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i49_4_lut_adj_557_LC_23_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i49_4_lut_adj_557_LC_23_20_3  (
            .in0(N__58186),
            .in1(N__58675),
            .in2(N__58171),
            .in3(N__58168),
            .lcout(\c0.n100_adj_3420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_374_LC_23_20_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_374_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_374_LC_23_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_374_LC_23_20_4  (
            .in0(N__64707),
            .in1(N__58368),
            .in2(N__58150),
            .in3(N__66243),
            .lcout(\c0.n12_adj_3208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_2_lut_3_lut_LC_23_20_5 .C_ON=1'b0;
    defparam \c0.i31_2_lut_3_lut_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i31_2_lut_3_lut_LC_23_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i31_2_lut_3_lut_LC_23_20_5  (
            .in0(N__67241),
            .in1(N__67265),
            .in2(_gnd_net_),
            .in3(N__58097),
            .lcout(\c0.n82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i42_4_lut_LC_23_20_6 .C_ON=1'b0;
    defparam \c0.i42_4_lut_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i42_4_lut_LC_23_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i42_4_lut_LC_23_20_6  (
            .in0(N__69853),
            .in1(N__67243),
            .in2(N__59179),
            .in3(N__58507),
            .lcout(\c0.n93_adj_3385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i31_2_lut_3_lut_adj_841_LC_23_20_7 .C_ON=1'b0;
    defparam \c0.i31_2_lut_3_lut_adj_841_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i31_2_lut_3_lut_adj_841_LC_23_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i31_2_lut_3_lut_adj_841_LC_23_20_7  (
            .in0(N__68018),
            .in1(N__58669),
            .in2(_gnd_net_),
            .in3(N__58633),
            .lcout(\c0.n68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_815_LC_23_21_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_815_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_815_LC_23_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_815_LC_23_21_0  (
            .in0(N__58606),
            .in1(N__58582),
            .in2(N__58573),
            .in3(N__60844),
            .lcout(\c0.n26_adj_3537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_21_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_23_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_2_lut_3_lut_4_lut_LC_23_21_1  (
            .in0(N__69682),
            .in1(N__69825),
            .in2(N__69657),
            .in3(N__69746),
            .lcout(\c0.n38_adj_3062 ),
            .ltout(\c0.n38_adj_3062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i42_2_lut_4_lut_LC_23_21_2 .C_ON=1'b0;
    defparam \c0.i42_2_lut_4_lut_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i42_2_lut_4_lut_LC_23_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i42_2_lut_4_lut_LC_23_21_2  (
            .in0(N__58551),
            .in1(N__69848),
            .in2(N__58510),
            .in3(N__58506),
            .lcout(\c0.n93_adj_3329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_816_LC_23_21_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_816_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_816_LC_23_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_816_LC_23_21_3  (
            .in0(N__66256),
            .in1(N__58468),
            .in2(N__58408),
            .in3(N__58381),
            .lcout(\c0.n20917 ),
            .ltout(\c0.n20917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_570_LC_23_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_570_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_570_LC_23_21_4 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_adj_570_LC_23_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__58375),
            .in3(N__72346),
            .lcout(),
            .ltout(\c0.n6_adj_3433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_572_LC_23_21_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_572_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_572_LC_23_21_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_572_LC_23_21_5  (
            .in0(N__58372),
            .in1(N__69745),
            .in2(N__58342),
            .in3(N__58942),
            .lcout(\c0.n18375 ),
            .ltout(\c0.n18375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_adj_636_LC_23_21_6 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_adj_636_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_adj_636_LC_23_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i7_2_lut_3_lut_adj_636_LC_23_21_6  (
            .in0(_gnd_net_),
            .in1(N__69652),
            .in2(N__58339),
            .in3(N__59039),
            .lcout(\c0.n32_adj_3310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i32_2_lut_LC_23_21_7 .C_ON=1'b0;
    defparam \c0.i32_2_lut_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i32_2_lut_LC_23_21_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i32_2_lut_LC_23_21_7  (
            .in0(N__69849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59165),
            .lcout(\c0.n83_adj_3442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_742_LC_23_22_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_742_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_4_lut_adj_742_LC_23_22_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_2_lut_3_lut_4_lut_adj_742_LC_23_22_0  (
            .in0(N__63741),
            .in1(N__58940),
            .in2(N__59137),
            .in3(N__59086),
            .lcout(\c0.n19_adj_3056 ),
            .ltout(\c0.n19_adj_3056_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_4_lut_adj_614_LC_23_22_1 .C_ON=1'b0;
    defparam \c0.i10_3_lut_4_lut_adj_614_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_4_lut_adj_614_LC_23_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_3_lut_4_lut_adj_614_LC_23_22_1  (
            .in0(N__69744),
            .in1(N__69817),
            .in2(N__59014),
            .in3(N__59002),
            .lcout(\c0.n29_adj_3454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_553_LC_23_22_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_553_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_553_LC_23_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_553_LC_23_22_2  (
            .in0(_gnd_net_),
            .in1(N__64983),
            .in2(_gnd_net_),
            .in3(N__58941),
            .lcout(\c0.n6_adj_3239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_325_LC_23_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_325_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_325_LC_23_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_325_LC_23_22_3  (
            .in0(_gnd_net_),
            .in1(N__58900),
            .in2(_gnd_net_),
            .in3(N__69683),
            .lcout(\c0.n19354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i184_LC_23_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i184_LC_23_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i184_LC_23_22_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i184_LC_23_22_4  (
            .in0(N__67527),
            .in1(N__72217),
            .in2(_gnd_net_),
            .in3(N__58822),
            .lcout(data_in_frame_22_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71209),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i180_LC_23_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i180_LC_23_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i180_LC_23_22_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0__i180_LC_23_22_5  (
            .in0(N__58790),
            .in1(N__67528),
            .in2(_gnd_net_),
            .in3(N__69381),
            .lcout(data_in_frame_22_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71209),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_284_LC_23_22_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_284_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_284_LC_23_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_284_LC_23_22_6  (
            .in0(N__58768),
            .in1(N__66661),
            .in2(N__58724),
            .in3(N__59191),
            .lcout(\c0.n20642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i132_LC_23_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i132_LC_23_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i132_LC_23_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i132_LC_23_22_7  (
            .in0(N__65605),
            .in1(N__69380),
            .in2(_gnd_net_),
            .in3(N__63742),
            .lcout(data_in_frame_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71209),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_759_LC_23_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_759_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_759_LC_23_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_759_LC_23_23_0  (
            .in0(N__66545),
            .in1(N__69565),
            .in2(N__59324),
            .in3(N__59511),
            .lcout(\c0.n17942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_23_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_23_23_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_921_LC_23_23_1  (
            .in0(N__71754),
            .in1(N__61456),
            .in2(_gnd_net_),
            .in3(N__59479),
            .lcout(n19128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i163_LC_23_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i163_LC_23_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i163_LC_23_23_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i163_LC_23_23_2  (
            .in0(N__67198),
            .in1(N__71755),
            .in2(N__67704),
            .in3(N__68712),
            .lcout(\c0.data_in_frame_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71221),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_283_LC_23_23_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_283_LC_23_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_283_LC_23_23_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_283_LC_23_23_3  (
            .in0(N__72385),
            .in1(N__59380),
            .in2(N__66514),
            .in3(N__59359),
            .lcout(\c0.n20709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i209_LC_23_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i209_LC_23_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i209_LC_23_23_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i209_LC_23_23_4  (
            .in0(N__65241),
            .in1(N__66979),
            .in2(N__59325),
            .in3(N__62848),
            .lcout(\c0.data_in_frame_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71221),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i210_LC_23_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i210_LC_23_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i210_LC_23_23_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i210_LC_23_23_5  (
            .in0(N__62847),
            .in1(N__71504),
            .in2(N__66987),
            .in3(N__66546),
            .lcout(\c0.data_in_frame_26_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71221),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i218_LC_23_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i218_LC_23_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i218_LC_23_23_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i218_LC_23_23_6  (
            .in0(N__71503),
            .in1(N__66980),
            .in2(N__59300),
            .in3(N__64583),
            .lcout(\c0.data_in_frame_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71221),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i219_LC_23_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i219_LC_23_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i219_LC_23_23_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i219_LC_23_23_7  (
            .in0(N__64582),
            .in1(N__68711),
            .in2(N__66988),
            .in3(N__59237),
            .lcout(\c0.data_in_frame_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71221),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_adj_528_LC_23_24_0 .C_ON=1'b0;
    defparam \c0.i26_4_lut_adj_528_LC_23_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_adj_528_LC_23_24_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i26_4_lut_adj_528_LC_23_24_0  (
            .in0(N__59549),
            .in1(N__59212),
            .in2(N__59784),
            .in3(N__59190),
            .lcout(),
            .ltout(\c0.n77_adj_3396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i39_4_lut_LC_23_24_1 .C_ON=1'b0;
    defparam \c0.i39_4_lut_LC_23_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i39_4_lut_LC_23_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i39_4_lut_LC_23_24_1  (
            .in0(N__68043),
            .in1(N__59832),
            .in2(N__59812),
            .in3(N__66589),
            .lcout(\c0.n90_adj_3400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_383_LC_23_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_383_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_383_LC_23_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_383_LC_23_24_2  (
            .in0(_gnd_net_),
            .in1(N__59548),
            .in2(_gnd_net_),
            .in3(N__59775),
            .lcout(),
            .ltout(\c0.n19214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_385_LC_23_24_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_385_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_385_LC_23_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_385_LC_23_24_3  (
            .in0(N__59743),
            .in1(N__59699),
            .in2(N__59623),
            .in3(N__59620),
            .lcout(\c0.n12_adj_3214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i207_LC_23_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i207_LC_23_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i207_LC_23_24_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i207_LC_23_24_4  (
            .in0(N__69040),
            .in1(N__66957),
            .in2(N__59556),
            .in3(N__63378),
            .lcout(\c0.data_in_frame_25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71228),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i120_LC_23_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i120_LC_23_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i120_LC_23_24_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i120_LC_23_24_5  (
            .in0(N__62034),
            .in1(N__64199),
            .in2(N__64942),
            .in3(N__72242),
            .lcout(\c0.data_in_frame_14_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71228),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3137_2_lut_LC_23_25_1 .C_ON=1'b0;
    defparam \c0.i3137_2_lut_LC_23_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3137_2_lut_LC_23_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3137_2_lut_LC_23_25_1  (
            .in0(_gnd_net_),
            .in1(N__64920),
            .in2(_gnd_net_),
            .in3(N__64888),
            .lcout(\c0.n5784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i124_LC_24_9_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i124_LC_24_9_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i124_LC_24_9_0 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i124_LC_24_9_0  (
            .in0(N__64183),
            .in1(N__64387),
            .in2(N__64683),
            .in3(N__69445),
            .lcout(\c0.data_in_frame_15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71233),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i121_LC_24_9_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i121_LC_24_9_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i121_LC_24_9_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i121_LC_24_9_1  (
            .in0(N__64386),
            .in1(N__64184),
            .in2(N__63534),
            .in3(N__65190),
            .lcout(\c0.data_in_frame_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71233),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_24_9_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_24_9_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_24_9_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i57_LC_24_9_2  (
            .in0(N__65189),
            .in1(N__61595),
            .in2(N__65397),
            .in3(N__64388),
            .lcout(\c0.data_in_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71233),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_238_LC_24_9_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_238_LC_24_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_238_LC_24_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_238_LC_24_9_3  (
            .in0(N__60829),
            .in1(N__62495),
            .in2(_gnd_net_),
            .in3(N__60792),
            .lcout(\c0.n5595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_357_Select_1_i6_2_lut_LC_24_9_4 .C_ON=1'b0;
    defparam \c0.select_357_Select_1_i6_2_lut_LC_24_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_357_Select_1_i6_2_lut_LC_24_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_357_Select_1_i6_2_lut_LC_24_9_4  (
            .in0(_gnd_net_),
            .in1(N__60128),
            .in2(_gnd_net_),
            .in3(N__60733),
            .lcout(\c0.n6_adj_3140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_24_9_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_24_9_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_24_9_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i49_LC_24_9_5  (
            .in0(N__61593),
            .in1(N__60478),
            .in2(N__62049),
            .in3(N__65191),
            .lcout(\c0.data_in_frame_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71233),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_24_9_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_24_9_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_24_9_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i51_LC_24_9_7  (
            .in0(N__61594),
            .in1(N__62041),
            .in2(N__60449),
            .in3(N__68746),
            .lcout(\c0.data_in_frame_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71233),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_24_10_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_24_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i11_LC_24_10_0  (
            .in0(N__68745),
            .in1(N__59869),
            .in2(_gnd_net_),
            .in3(N__60398),
            .lcout(data_in_frame_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71232),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2593_2_lut_LC_24_10_1 .C_ON=1'b0;
    defparam \c0.i2593_2_lut_LC_24_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2593_2_lut_LC_24_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2593_2_lut_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(N__62512),
            .in2(_gnd_net_),
            .in3(N__61826),
            .lcout(\c0.n5240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_24_10_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_24_10_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i47_LC_24_10_2  (
            .in0(N__61550),
            .in1(N__60353),
            .in2(N__62359),
            .in3(N__68844),
            .lcout(\c0.data_in_frame_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71232),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_866_LC_24_10_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_866_LC_24_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_866_LC_24_10_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_866_LC_24_10_3  (
            .in0(N__60273),
            .in1(N__61549),
            .in2(N__60133),
            .in3(N__60001),
            .lcout(n19100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_793_LC_24_10_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_793_LC_24_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_793_LC_24_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_793_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(N__62206),
            .in2(_gnd_net_),
            .in3(N__62181),
            .lcout(\c0.n7 ),
            .ltout(\c0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_24_10_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_24_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_24_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(N__62076),
            .in2(N__62062),
            .in3(N__60987),
            .lcout(\c0.n12_adj_2998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_24_10_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_24_10_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_24_10_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i55_LC_24_10_6  (
            .in0(N__61551),
            .in1(N__68843),
            .in2(N__62522),
            .in3(N__62040),
            .lcout(\c0.data_in_frame_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71232),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_24_10_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_24_10_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_24_10_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i56_LC_24_10_7  (
            .in0(N__62039),
            .in1(N__61552),
            .in2(N__61861),
            .in3(N__72207),
            .lcout(\c0.data_in_frame_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71232),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_24_11_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_24_11_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i29_LC_24_11_0  (
            .in0(N__72698),
            .in1(N__61560),
            .in2(N__61345),
            .in3(N__61453),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71229),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_221_LC_24_11_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_221_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_221_LC_24_11_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_221_LC_24_11_2  (
            .in0(N__61306),
            .in1(N__61300),
            .in2(N__61011),
            .in3(N__61126),
            .lcout(\c0.n11953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_724_LC_24_11_4 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_724_LC_24_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_724_LC_24_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_adj_724_LC_24_11_4  (
            .in0(N__61261),
            .in1(N__61227),
            .in2(N__63166),
            .in3(N__60901),
            .lcout(\c0.n55_adj_3500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_599_LC_24_11_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_599_LC_24_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_599_LC_24_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_599_LC_24_11_5  (
            .in0(N__61127),
            .in1(N__61018),
            .in2(N__61012),
            .in3(N__60976),
            .lcout(\c0.data_out_frame_0__7__N_1540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_729_LC_24_11_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_729_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_729_LC_24_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_729_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(N__62343),
            .in2(_gnd_net_),
            .in3(N__60900),
            .lcout(\c0.n6_adj_3037 ),
            .ltout(\c0.n6_adj_3037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_266_LC_24_11_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_266_LC_24_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_266_LC_24_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_266_LC_24_11_7  (
            .in0(N__62658),
            .in1(N__62635),
            .in2(N__62629),
            .in3(N__62620),
            .lcout(\c0.n19560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_235_LC_24_12_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_235_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_235_LC_24_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_235_LC_24_12_1  (
            .in0(N__62935),
            .in1(N__63099),
            .in2(N__62544),
            .in3(N__62523),
            .lcout(\c0.n19258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_863_LC_24_12_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_863_LC_24_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_863_LC_24_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_863_LC_24_12_6  (
            .in0(N__62440),
            .in1(N__62382),
            .in2(_gnd_net_),
            .in3(N__62355),
            .lcout(\c0.n8_adj_3020 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i108_LC_24_13_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i108_LC_24_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i108_LC_24_13_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i108_LC_24_13_0  (
            .in0(N__71971),
            .in1(N__66146),
            .in2(N__62309),
            .in3(N__69410),
            .lcout(\c0.data_in_frame_13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i94_LC_24_13_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i94_LC_24_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i94_LC_24_13_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i94_LC_24_13_1  (
            .in0(N__67932),
            .in1(N__63201),
            .in2(N__66188),
            .in3(N__64550),
            .lcout(\c0.data_in_frame_11_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i75_LC_24_13_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i75_LC_24_13_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i75_LC_24_13_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i75_LC_24_13_2  (
            .in0(N__68726),
            .in1(N__63415),
            .in2(N__62254),
            .in3(N__66153),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i92_LC_24_13_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i92_LC_24_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i92_LC_24_13_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i92_LC_24_13_3  (
            .in0(N__69414),
            .in1(N__64549),
            .in2(N__66187),
            .in3(N__63066),
            .lcout(\c0.data_in_frame_11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i154_LC_24_13_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i154_LC_24_13_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i154_LC_24_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i154_LC_24_13_4  (
            .in0(N__71526),
            .in1(N__69169),
            .in2(_gnd_net_),
            .in3(N__65661),
            .lcout(data_in_frame_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i76_LC_24_13_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i76_LC_24_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i76_LC_24_13_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i76_LC_24_13_5  (
            .in0(N__63414),
            .in1(N__63224),
            .in2(N__69437),
            .in3(N__66144),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71210),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_316_LC_24_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_316_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_316_LC_24_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_316_LC_24_13_6  (
            .in0(_gnd_net_),
            .in1(N__63218),
            .in2(_gnd_net_),
            .in3(N__63197),
            .lcout(\c0.n5_adj_3043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_909_LC_24_13_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_909_LC_24_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_909_LC_24_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_909_LC_24_13_7  (
            .in0(N__63162),
            .in1(N__63100),
            .in2(_gnd_net_),
            .in3(N__63065),
            .lcout(\c0.n19381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_708_LC_24_14_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_708_LC_24_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_708_LC_24_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_708_LC_24_14_0  (
            .in0(N__62927),
            .in1(N__64039),
            .in2(N__62724),
            .in3(N__63044),
            .lcout(\c0.n11_adj_3492 ),
            .ltout(\c0.n11_adj_3492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_798_LC_24_14_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_798_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_798_LC_24_14_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_798_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62995),
            .in3(N__62988),
            .lcout(\c0.n20_adj_3527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i90_LC_24_14_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i90_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i90_LC_24_14_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i90_LC_24_14_2  (
            .in0(N__71527),
            .in1(N__64548),
            .in2(N__62934),
            .in3(N__66067),
            .lcout(\c0.data_in_frame_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71197),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_711_LC_24_14_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_711_LC_24_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_711_LC_24_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_711_LC_24_14_3  (
            .in0(N__65398),
            .in1(N__62716),
            .in2(N__62878),
            .in3(N__62926),
            .lcout(\c0.n19229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i91_LC_24_14_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i91_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i91_LC_24_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i91_LC_24_14_4  (
            .in0(N__66139),
            .in1(N__64546),
            .in2(N__62885),
            .in3(N__68727),
            .lcout(\c0.data_in_frame_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71197),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i88_LC_24_14_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i88_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i88_LC_24_14_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i88_LC_24_14_5  (
            .in0(N__62811),
            .in1(N__66140),
            .in2(N__62725),
            .in3(N__72145),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71197),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i96_LC_24_14_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i96_LC_24_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i96_LC_24_14_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i96_LC_24_14_6  (
            .in0(N__72144),
            .in1(N__64547),
            .in2(N__66186),
            .in3(N__64442),
            .lcout(\c0.data_in_frame_11_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71197),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i126_LC_24_14_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i126_LC_24_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i126_LC_24_14_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i126_LC_24_14_7  (
            .in0(N__67921),
            .in1(N__64397),
            .in2(N__64049),
            .in3(N__64250),
            .lcout(\c0.data_in_frame_15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71197),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_adj_934_LC_24_15_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_adj_934_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_adj_934_LC_24_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_adj_934_LC_24_15_1  (
            .in0(N__65495),
            .in1(N__63795),
            .in2(_gnd_net_),
            .in3(N__63766),
            .lcout(),
            .ltout(\c0.n9_adj_3552_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_881_LC_24_15_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_881_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_881_LC_24_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_881_LC_24_15_2  (
            .in0(N__72425),
            .in1(N__63805),
            .in2(N__64021),
            .in3(N__64013),
            .lcout(\c0.n25_adj_3553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i149_LC_24_15_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i149_LC_24_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i149_LC_24_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i149_LC_24_15_3  (
            .in0(N__63871),
            .in1(N__72700),
            .in2(_gnd_net_),
            .in3(N__63955),
            .lcout(data_in_frame_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71186),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_224_LC_24_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_224_LC_24_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_224_LC_24_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_224_LC_24_15_4  (
            .in0(_gnd_net_),
            .in1(N__63870),
            .in2(_gnd_net_),
            .in3(N__63861),
            .lcout(\c0.n7_adj_3000 ),
            .ltout(\c0.n7_adj_3000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_932_LC_24_15_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_932_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_932_LC_24_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_932_LC_24_15_5  (
            .in0(N__65494),
            .in1(N__63794),
            .in2(N__63781),
            .in3(N__63765),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_2_lut_3_lut_4_lut_LC_24_15_6 .C_ON=1'b0;
    defparam \c0.i19_2_lut_3_lut_4_lut_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19_2_lut_3_lut_4_lut_LC_24_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_2_lut_3_lut_4_lut_LC_24_15_6  (
            .in0(N__63687),
            .in1(N__63646),
            .in2(N__63573),
            .in3(N__63494),
            .lcout(\c0.n45_adj_3138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_834_LC_24_15_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_834_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_834_LC_24_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_834_LC_24_15_7  (
            .in0(_gnd_net_),
            .in1(N__65429),
            .in2(_gnd_net_),
            .in3(N__65399),
            .lcout(\c0.n7_adj_3355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_24_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_24_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_24_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_630_LC_24_16_0  (
            .in0(N__65299),
            .in1(N__65321),
            .in2(_gnd_net_),
            .in3(N__64770),
            .lcout(\c0.n4_adj_3435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_631_LC_24_16_1 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_631_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_631_LC_24_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_631_LC_24_16_1  (
            .in0(N__65320),
            .in1(N__65618),
            .in2(_gnd_net_),
            .in3(N__65298),
            .lcout(\c0.n14_adj_3449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i158_LC_24_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i158_LC_24_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i158_LC_24_16_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i158_LC_24_16_2  (
            .in0(N__69167),
            .in1(N__67971),
            .in2(_gnd_net_),
            .in3(N__65715),
            .lcout(data_in_frame_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71174),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i161_LC_24_16_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i161_LC_24_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i161_LC_24_16_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i161_LC_24_16_3  (
            .in0(N__71740),
            .in1(N__65226),
            .in2(N__69777),
            .in3(N__67218),
            .lcout(\c0.data_in_frame_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71174),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_782_LC_24_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_782_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_782_LC_24_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_782_LC_24_16_5  (
            .in0(N__64972),
            .in1(N__64950),
            .in2(_gnd_net_),
            .in3(N__64900),
            .lcout(\c0.n19554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_754_LC_24_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_754_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_754_LC_24_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_754_LC_24_16_6  (
            .in0(N__65619),
            .in1(N__64771),
            .in2(_gnd_net_),
            .in3(N__68308),
            .lcout(\c0.n18_adj_3235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_676_LC_24_16_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_676_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_676_LC_24_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i5_3_lut_adj_676_LC_24_16_7  (
            .in0(N__64699),
            .in1(N__64645),
            .in2(_gnd_net_),
            .in3(N__64608),
            .lcout(\c0.n20576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i164_LC_24_17_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i164_LC_24_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i164_LC_24_17_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i164_LC_24_17_0  (
            .in0(N__67224),
            .in1(N__68084),
            .in2(N__69363),
            .in3(N__71739),
            .lcout(\c0.data_in_frame_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71147),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_789_LC_24_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_789_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_789_LC_24_17_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_789_LC_24_17_1  (
            .in0(_gnd_net_),
            .in1(N__68070),
            .in2(_gnd_net_),
            .in3(N__68195),
            .lcout(\c0.n19251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_814_LC_24_17_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_814_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_814_LC_24_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_814_LC_24_17_2  (
            .in0(N__66361),
            .in1(N__66337),
            .in2(N__66310),
            .in3(N__66298),
            .lcout(\c0.n22_adj_3535 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i165_LC_24_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i165_LC_24_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i165_LC_24_17_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i165_LC_24_17_3  (
            .in0(N__72699),
            .in1(N__67226),
            .in2(N__71781),
            .in3(N__68196),
            .lcout(\c0.data_in_frame_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71147),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i162_LC_24_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i162_LC_24_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i162_LC_24_17_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i162_LC_24_17_4  (
            .in0(N__67223),
            .in1(N__71738),
            .in2(N__66239),
            .in3(N__71524),
            .lcout(\c0.data_in_frame_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71147),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i100_LC_24_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i100_LC_24_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i100_LC_24_17_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i100_LC_24_17_5  (
            .in0(N__66185),
            .in1(N__67225),
            .in2(N__65869),
            .in3(N__69316),
            .lcout(\c0.data_in_frame_12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71147),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_617_LC_24_17_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_617_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_617_LC_24_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_617_LC_24_17_6  (
            .in0(N__65780),
            .in1(N__65711),
            .in2(N__65674),
            .in3(N__69492),
            .lcout(\c0.n6166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i131_LC_24_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i131_LC_24_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i131_LC_24_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i131_LC_24_17_7  (
            .in0(N__65580),
            .in1(N__68750),
            .in2(_gnd_net_),
            .in3(N__65493),
            .lcout(data_in_frame_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71147),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i230_LC_24_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i230_LC_24_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i230_LC_24_18_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i230_LC_24_18_0  (
            .in0(N__65448),
            .in1(N__66956),
            .in2(N__67944),
            .in3(N__67227),
            .lcout(\c0.data_in_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71175),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i228_LC_24_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i228_LC_24_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i228_LC_24_18_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i228_LC_24_18_1  (
            .in0(N__66953),
            .in1(N__69277),
            .in2(N__67231),
            .in3(N__66571),
            .lcout(\c0.data_in_frame_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71175),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i236_LC_24_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i236_LC_24_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i236_LC_24_18_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i236_LC_24_18_2  (
            .in0(N__69278),
            .in1(N__66955),
            .in2(N__67020),
            .in3(N__71958),
            .lcout(\c0.data_in_frame_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71175),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i238_LC_24_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i238_LC_24_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i238_LC_24_18_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i238_LC_24_18_3  (
            .in0(N__66954),
            .in1(N__67889),
            .in2(N__71973),
            .in3(N__66690),
            .lcout(\c0.data_in_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71175),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_712_LC_24_18_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_712_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_712_LC_24_18_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_712_LC_24_18_4  (
            .in0(N__68245),
            .in1(N__69834),
            .in2(N__72851),
            .in3(N__66673),
            .lcout(\c0.n20503 ),
            .ltout(\c0.n20503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_718_LC_24_18_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_718_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_718_LC_24_18_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_718_LC_24_18_5  (
            .in0(N__66648),
            .in1(N__66427),
            .in2(N__66604),
            .in3(N__66601),
            .lcout(\c0.n27_adj_3399 ),
            .ltout(\c0.n27_adj_3399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_adj_549_LC_24_18_6 .C_ON=1'b0;
    defparam \c0.i27_4_lut_adj_549_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_adj_549_LC_24_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_adj_549_LC_24_18_6  (
            .in0(N__69937),
            .in1(N__66570),
            .in2(N__66559),
            .in3(N__66556),
            .lcout(\c0.n78_adj_3414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_715_LC_24_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_715_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_715_LC_24_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_715_LC_24_18_7  (
            .in0(N__66510),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66464),
            .lcout(\c0.n19487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_892_LC_24_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_892_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_892_LC_24_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_892_LC_24_19_0  (
            .in0(N__70063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66416),
            .lcout(\c0.n19484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_842_LC_24_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_842_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_842_LC_24_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_842_LC_24_19_1  (
            .in0(N__69079),
            .in1(N__67614),
            .in2(N__69564),
            .in3(N__69648),
            .lcout(),
            .ltout(\c0.n7_adj_3072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_299_LC_24_19_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_299_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_299_LC_24_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_299_LC_24_19_2  (
            .in0(N__67582),
            .in1(N__70494),
            .in2(N__67576),
            .in3(N__67360),
            .lcout(\c0.n18413 ),
            .ltout(\c0.n18413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_289_LC_24_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_289_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_289_LC_24_19_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_289_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67573),
            .in3(N__67570),
            .lcout(\c0.n18525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i182_LC_24_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i182_LC_24_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i182_LC_24_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i182_LC_24_19_4  (
            .in0(N__67529),
            .in1(N__67940),
            .in2(_gnd_net_),
            .in3(N__67427),
            .lcout(data_in_frame_22_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71187),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_297_LC_24_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_297_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_297_LC_24_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_297_LC_24_19_5  (
            .in0(N__70016),
            .in1(N__67408),
            .in2(_gnd_net_),
            .in3(N__67387),
            .lcout(\c0.n8_adj_3070 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_796_LC_24_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_796_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_796_LC_24_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_796_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(N__69557),
            .in2(_gnd_net_),
            .in3(N__69078),
            .lcout(\c0.n19315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_882_LC_24_19_7 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_882_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_882_LC_24_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_882_LC_24_19_7  (
            .in0(N__67348),
            .in1(N__67330),
            .in2(N__67315),
            .in3(N__67302),
            .lcout(\c0.n17832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i159_LC_24_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i159_LC_24_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i159_LC_24_20_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_in_frame_0__i159_LC_24_20_0  (
            .in0(_gnd_net_),
            .in1(N__69151),
            .in2(N__72342),
            .in3(N__69006),
            .lcout(data_in_frame_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71198),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_2_lut_3_lut_adj_574_LC_24_20_1 .C_ON=1'b0;
    defparam \c0.i7_2_lut_3_lut_adj_574_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_2_lut_3_lut_adj_574_LC_24_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_2_lut_3_lut_adj_574_LC_24_20_1  (
            .in0(N__68104),
            .in1(N__68213),
            .in2(_gnd_net_),
            .in3(N__67629),
            .lcout(\c0.n40_adj_3271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i157_LC_24_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i157_LC_24_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i157_LC_24_20_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i157_LC_24_20_2  (
            .in0(N__72754),
            .in1(N__69150),
            .in2(_gnd_net_),
            .in3(N__72827),
            .lcout(data_in_frame_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71198),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i175_LC_24_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i175_LC_24_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i175_LC_24_20_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i175_LC_24_20_3  (
            .in0(N__71779),
            .in1(N__71960),
            .in2(N__72473),
            .in3(N__69007),
            .lcout(\c0.data_in_frame_21_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71198),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i171_LC_24_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i171_LC_24_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i171_LC_24_20_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i171_LC_24_20_4  (
            .in0(N__71959),
            .in1(N__71780),
            .in2(N__69896),
            .in3(N__68682),
            .lcout(\c0.data_in_frame_21_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71198),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_573_LC_24_20_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_573_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_573_LC_24_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_573_LC_24_20_5  (
            .in0(N__68429),
            .in1(N__68384),
            .in2(N__69555),
            .in3(N__68307),
            .lcout(\c0.n14_adj_3436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_871_LC_24_20_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_871_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_871_LC_24_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_871_LC_24_20_6  (
            .in0(N__69658),
            .in1(N__68234),
            .in2(N__68173),
            .in3(N__68105),
            .lcout(\c0.n54_adj_3388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_2_lut_LC_24_20_7 .C_ON=1'b0;
    defparam \c0.i16_2_lut_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i16_2_lut_LC_24_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i16_2_lut_LC_24_20_7  (
            .in0(_gnd_net_),
            .in1(N__69707),
            .in2(_gnd_net_),
            .in3(N__68017),
            .lcout(\c0.n43_adj_3131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i174_LC_24_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i174_LC_24_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i174_LC_24_21_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i174_LC_24_21_0  (
            .in0(N__67964),
            .in1(N__71801),
            .in2(N__69556),
            .in3(N__71964),
            .lcout(\c0.data_in_frame_21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71211),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_684_LC_24_21_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_684_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_684_LC_24_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_684_LC_24_21_1  (
            .in0(N__72304),
            .in1(N__70069),
            .in2(N__67705),
            .in3(N__67674),
            .lcout(\c0.n22_adj_3322 ),
            .ltout(\c0.n22_adj_3322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_4_lut_LC_24_21_2 .C_ON=1'b0;
    defparam \c0.i5_2_lut_4_lut_LC_24_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_4_lut_LC_24_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_2_lut_4_lut_LC_24_21_2  (
            .in0(N__69510),
            .in1(N__69879),
            .in2(N__69922),
            .in3(N__71266),
            .lcout(\c0.n36_adj_3090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_2_lut_4_lut_LC_24_21_3 .C_ON=1'b0;
    defparam \c0.i8_2_lut_4_lut_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_2_lut_4_lut_LC_24_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_2_lut_4_lut_LC_24_21_3  (
            .in0(N__71265),
            .in1(N__69772),
            .in2(N__69889),
            .in3(N__69509),
            .lcout(\c0.n29_adj_3383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_589_LC_24_21_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_589_LC_24_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_589_LC_24_21_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i2_2_lut_adj_589_LC_24_21_4  (
            .in0(N__69748),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69827),
            .lcout(\c0.n18415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_adj_699_LC_24_21_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_adj_699_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_adj_699_LC_24_21_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i6_2_lut_3_lut_adj_699_LC_24_21_5  (
            .in0(N__69826),
            .in1(N__69773),
            .in2(_gnd_net_),
            .in3(N__69747),
            .lcout(\c0.n6_adj_3091 ),
            .ltout(\c0.n6_adj_3091_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_634_LC_24_21_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_634_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_634_LC_24_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_634_LC_24_21_6  (
            .in0(N__70481),
            .in1(N__69684),
            .in2(N__69661),
            .in3(N__69656),
            .lcout(\c0.n18498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_548_LC_24_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_548_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_548_LC_24_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_548_LC_24_21_7  (
            .in0(_gnd_net_),
            .in1(N__69595),
            .in2(_gnd_net_),
            .in3(N__69543),
            .lcout(\c0.n19321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_618_LC_24_22_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_618_LC_24_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_618_LC_24_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_618_LC_24_22_0  (
            .in0(N__72335),
            .in1(N__69055),
            .in2(N__72844),
            .in3(N__69458),
            .lcout(\c0.n12037 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i160_LC_24_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i160_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i160_LC_24_22_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_frame_0__i160_LC_24_22_1  (
            .in0(N__69138),
            .in1(_gnd_net_),
            .in2(N__69465),
            .in3(N__72254),
            .lcout(data_in_frame_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71222),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i156_LC_24_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i156_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i156_LC_24_22_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_frame_0__i156_LC_24_22_2  (
            .in0(N__69422),
            .in1(N__69139),
            .in2(_gnd_net_),
            .in3(N__69056),
            .lcout(data_in_frame_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71222),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_295_LC_24_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_295_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_295_LC_24_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_295_LC_24_22_3  (
            .in0(_gnd_net_),
            .in1(N__71998),
            .in2(_gnd_net_),
            .in3(N__72336),
            .lcout(\c0.n19162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_296_LC_24_22_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_296_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_296_LC_24_22_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_296_LC_24_22_4  (
            .in0(N__70464),
            .in1(N__69933),
            .in2(N__70224),
            .in3(N__70188),
            .lcout(\c0.n20332 ),
            .ltout(\c0.n20332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_301_LC_24_22_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_301_LC_24_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_301_LC_24_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_301_LC_24_22_5  (
            .in0(N__70389),
            .in1(N__70339),
            .in2(N__70291),
            .in3(N__70288),
            .lcout(\c0.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_541_LC_24_22_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_541_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_541_LC_24_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_541_LC_24_22_6  (
            .in0(N__70257),
            .in1(N__70243),
            .in2(N__70225),
            .in3(N__70189),
            .lcout(\c0.n10_adj_3410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_adj_578_LC_24_22_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_adj_578_LC_24_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_adj_578_LC_24_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i4_2_lut_3_lut_adj_578_LC_24_22_7  (
            .in0(N__70161),
            .in1(N__70124),
            .in2(_gnd_net_),
            .in3(N__70084),
            .lcout(\c0.n12_adj_3439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_846_LC_24_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_846_LC_24_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_846_LC_24_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_846_LC_24_23_0  (
            .in0(N__70056),
            .in1(N__71993),
            .in2(_gnd_net_),
            .in3(N__72467),
            .lcout(),
            .ltout(\c0.n4_adj_3067_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_293_LC_24_23_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_293_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_293_LC_24_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_293_LC_24_23_1  (
            .in0(N__72781),
            .in1(N__70017),
            .in2(N__69991),
            .in3(N__69987),
            .lcout(\c0.n19369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_592_LC_24_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_592_LC_24_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_592_LC_24_23_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_592_LC_24_23_2  (
            .in0(N__72338),
            .in1(N__72831),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n11669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i173_LC_24_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i173_LC_24_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i173_LC_24_23_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i173_LC_24_23_3  (
            .in0(N__71962),
            .in1(N__71745),
            .in2(N__72393),
            .in3(N__72740),
            .lcout(\c0.data_in_frame_21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71230),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_660_LC_24_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_660_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_660_LC_24_23_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_660_LC_24_23_4  (
            .in0(_gnd_net_),
            .in1(N__71992),
            .in2(_gnd_net_),
            .in3(N__72466),
            .lcout(),
            .ltout(\c0.n11939_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_679_LC_24_23_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_679_LC_24_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_679_LC_24_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_679_LC_24_23_5  (
            .in0(N__72439),
            .in1(N__72369),
            .in2(N__72349),
            .in3(N__72337),
            .lcout(\c0.n13_adj_3485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i176_LC_24_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i176_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i176_LC_24_23_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i176_LC_24_23_6  (
            .in0(N__72256),
            .in1(N__71963),
            .in2(N__71782),
            .in3(N__71994),
            .lcout(\c0.data_in_frame_21_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71230),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i170_LC_24_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i170_LC_24_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i170_LC_24_23_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i170_LC_24_23_7  (
            .in0(N__71961),
            .in1(N__71744),
            .in2(N__71273),
            .in3(N__71547),
            .lcout(\c0.data_in_frame_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__71230),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
