// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 16:24:44

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__35917;
    wire N__35916;
    wire N__35915;
    wire N__35908;
    wire N__35907;
    wire N__35906;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35881;
    wire N__35880;
    wire N__35879;
    wire N__35872;
    wire N__35871;
    wire N__35870;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35832;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35817;
    wire N__35816;
    wire N__35815;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35758;
    wire N__35745;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35736;
    wire N__35735;
    wire N__35732;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35704;
    wire N__35699;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35689;
    wire N__35684;
    wire N__35683;
    wire N__35682;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35661;
    wire N__35658;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35638;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35617;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35580;
    wire N__35577;
    wire N__35574;
    wire N__35573;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35556;
    wire N__35555;
    wire N__35554;
    wire N__35553;
    wire N__35552;
    wire N__35551;
    wire N__35550;
    wire N__35547;
    wire N__35546;
    wire N__35545;
    wire N__35540;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35536;
    wire N__35535;
    wire N__35534;
    wire N__35531;
    wire N__35526;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35513;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35498;
    wire N__35493;
    wire N__35486;
    wire N__35475;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35453;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35436;
    wire N__35435;
    wire N__35434;
    wire N__35433;
    wire N__35432;
    wire N__35431;
    wire N__35430;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35423;
    wire N__35422;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35418;
    wire N__35417;
    wire N__35416;
    wire N__35415;
    wire N__35414;
    wire N__35413;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35402;
    wire N__35401;
    wire N__35400;
    wire N__35399;
    wire N__35398;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35389;
    wire N__35388;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35369;
    wire N__35368;
    wire N__35367;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35363;
    wire N__35362;
    wire N__35361;
    wire N__35360;
    wire N__35359;
    wire N__35358;
    wire N__35357;
    wire N__35356;
    wire N__35355;
    wire N__35354;
    wire N__35353;
    wire N__35352;
    wire N__35351;
    wire N__35350;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35346;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35341;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35335;
    wire N__35334;
    wire N__35333;
    wire N__35332;
    wire N__35331;
    wire N__35330;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35323;
    wire N__35322;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35318;
    wire N__35317;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35292;
    wire N__35291;
    wire N__35290;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34826;
    wire N__34825;
    wire N__34822;
    wire N__34817;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34789;
    wire N__34780;
    wire N__34771;
    wire N__34768;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34697;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34624;
    wire N__34619;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34600;
    wire N__34595;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34551;
    wire N__34548;
    wire N__34547;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34524;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34480;
    wire N__34479;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34463;
    wire N__34454;
    wire N__34443;
    wire N__34440;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34419;
    wire N__34414;
    wire N__34411;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34397;
    wire N__34394;
    wire N__34389;
    wire N__34384;
    wire N__34381;
    wire N__34376;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34352;
    wire N__34351;
    wire N__34350;
    wire N__34349;
    wire N__34348;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34340;
    wire N__34339;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34329;
    wire N__34322;
    wire N__34319;
    wire N__34308;
    wire N__34295;
    wire N__34284;
    wire N__34283;
    wire N__34282;
    wire N__34281;
    wire N__34280;
    wire N__34279;
    wire N__34278;
    wire N__34277;
    wire N__34276;
    wire N__34275;
    wire N__34274;
    wire N__34273;
    wire N__34272;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34254;
    wire N__34239;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34218;
    wire N__34213;
    wire N__34208;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34200;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34178;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34157;
    wire N__34156;
    wire N__34155;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34140;
    wire N__34137;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34101;
    wire N__34098;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34052;
    wire N__34047;
    wire N__34044;
    wire N__34043;
    wire N__34038;
    wire N__34035;
    wire N__34034;
    wire N__34033;
    wire N__34032;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34017;
    wire N__34008;
    wire N__34005;
    wire N__34004;
    wire N__34003;
    wire N__34000;
    wire N__33995;
    wire N__33990;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33981;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33973;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33958;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33920;
    wire N__33919;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33913;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33907;
    wire N__33900;
    wire N__33897;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33878;
    wire N__33875;
    wire N__33864;
    wire N__33861;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33842;
    wire N__33839;
    wire N__33838;
    wire N__33837;
    wire N__33836;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33824;
    wire N__33823;
    wire N__33822;
    wire N__33821;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33806;
    wire N__33801;
    wire N__33796;
    wire N__33793;
    wire N__33780;
    wire N__33779;
    wire N__33778;
    wire N__33777;
    wire N__33776;
    wire N__33771;
    wire N__33770;
    wire N__33767;
    wire N__33762;
    wire N__33759;
    wire N__33758;
    wire N__33755;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33735;
    wire N__33732;
    wire N__33731;
    wire N__33728;
    wire N__33727;
    wire N__33726;
    wire N__33725;
    wire N__33724;
    wire N__33723;
    wire N__33720;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33706;
    wire N__33701;
    wire N__33700;
    wire N__33697;
    wire N__33688;
    wire N__33685;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33666;
    wire N__33661;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33611;
    wire N__33608;
    wire N__33603;
    wire N__33600;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33585;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33543;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33531;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33506;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33483;
    wire N__33482;
    wire N__33477;
    wire N__33474;
    wire N__33473;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33461;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33432;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33408;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33396;
    wire N__33395;
    wire N__33392;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33376;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33358;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33338;
    wire N__33333;
    wire N__33330;
    wire N__33329;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33303;
    wire N__33302;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33280;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33228;
    wire N__33225;
    wire N__33220;
    wire N__33217;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33201;
    wire N__33200;
    wire N__33199;
    wire N__33194;
    wire N__33193;
    wire N__33192;
    wire N__33191;
    wire N__33190;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33178;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33174;
    wire N__33173;
    wire N__33164;
    wire N__33161;
    wire N__33152;
    wire N__33151;
    wire N__33150;
    wire N__33149;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33130;
    wire N__33125;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33096;
    wire N__33095;
    wire N__33092;
    wire N__33091;
    wire N__33090;
    wire N__33085;
    wire N__33082;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33064;
    wire N__33057;
    wire N__33054;
    wire N__33047;
    wire N__33042;
    wire N__33035;
    wire N__33034;
    wire N__33033;
    wire N__33032;
    wire N__33031;
    wire N__33030;
    wire N__33029;
    wire N__33028;
    wire N__33025;
    wire N__33024;
    wire N__33023;
    wire N__33020;
    wire N__33019;
    wire N__33018;
    wire N__33015;
    wire N__33014;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32966;
    wire N__32963;
    wire N__32958;
    wire N__32957;
    wire N__32956;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32945;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32922;
    wire N__32919;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32885;
    wire N__32884;
    wire N__32883;
    wire N__32878;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32867;
    wire N__32860;
    wire N__32857;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32843;
    wire N__32840;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32815;
    wire N__32812;
    wire N__32807;
    wire N__32806;
    wire N__32799;
    wire N__32796;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32775;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32742;
    wire N__32733;
    wire N__32728;
    wire N__32709;
    wire N__32706;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32678;
    wire N__32675;
    wire N__32668;
    wire N__32663;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32556;
    wire N__32555;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32538;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32509;
    wire N__32508;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32474;
    wire N__32471;
    wire N__32466;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32378;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32349;
    wire N__32348;
    wire N__32345;
    wire N__32344;
    wire N__32339;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32319;
    wire N__32310;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32273;
    wire N__32272;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32233;
    wire N__32230;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32198;
    wire N__32193;
    wire N__32190;
    wire N__32185;
    wire N__32182;
    wire N__32179;
    wire N__32172;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32164;
    wire N__32161;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32128;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32105;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32063;
    wire N__32058;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32044;
    wire N__32043;
    wire N__32042;
    wire N__32041;
    wire N__32040;
    wire N__32039;
    wire N__32038;
    wire N__32037;
    wire N__32036;
    wire N__32035;
    wire N__32034;
    wire N__32033;
    wire N__32032;
    wire N__32031;
    wire N__32030;
    wire N__32027;
    wire N__32022;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32012;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31972;
    wire N__31971;
    wire N__31968;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31956;
    wire N__31953;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31897;
    wire N__31894;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31853;
    wire N__31850;
    wire N__31837;
    wire N__31834;
    wire N__31829;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31807;
    wire N__31804;
    wire N__31797;
    wire N__31788;
    wire N__31785;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31763;
    wire N__31754;
    wire N__31749;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31731;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31686;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31678;
    wire N__31675;
    wire N__31674;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31647;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31631;
    wire N__31630;
    wire N__31629;
    wire N__31628;
    wire N__31627;
    wire N__31620;
    wire N__31619;
    wire N__31618;
    wire N__31617;
    wire N__31616;
    wire N__31615;
    wire N__31614;
    wire N__31607;
    wire N__31606;
    wire N__31605;
    wire N__31604;
    wire N__31601;
    wire N__31594;
    wire N__31587;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31580;
    wire N__31573;
    wire N__31572;
    wire N__31571;
    wire N__31570;
    wire N__31569;
    wire N__31564;
    wire N__31561;
    wire N__31556;
    wire N__31553;
    wire N__31552;
    wire N__31551;
    wire N__31548;
    wire N__31543;
    wire N__31536;
    wire N__31533;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31521;
    wire N__31516;
    wire N__31513;
    wire N__31506;
    wire N__31503;
    wire N__31498;
    wire N__31493;
    wire N__31488;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31461;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31446;
    wire N__31443;
    wire N__31436;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31415;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31399;
    wire N__31396;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31379;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31360;
    wire N__31355;
    wire N__31352;
    wire N__31347;
    wire N__31344;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31303;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31259;
    wire N__31256;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31245;
    wire N__31244;
    wire N__31243;
    wire N__31242;
    wire N__31239;
    wire N__31234;
    wire N__31233;
    wire N__31232;
    wire N__31231;
    wire N__31230;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31204;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31193;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31179;
    wire N__31178;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31141;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31123;
    wire N__31116;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31076;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31058;
    wire N__31055;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31022;
    wire N__31021;
    wire N__31020;
    wire N__31017;
    wire N__31016;
    wire N__31013;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30992;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30965;
    wire N__30964;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30952;
    wire N__30947;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30920;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30912;
    wire N__30911;
    wire N__30910;
    wire N__30909;
    wire N__30904;
    wire N__30895;
    wire N__30892;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30875;
    wire N__30874;
    wire N__30873;
    wire N__30870;
    wire N__30869;
    wire N__30868;
    wire N__30867;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30849;
    wire N__30846;
    wire N__30837;
    wire N__30836;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30789;
    wire N__30788;
    wire N__30787;
    wire N__30786;
    wire N__30785;
    wire N__30784;
    wire N__30783;
    wire N__30778;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30760;
    wire N__30757;
    wire N__30752;
    wire N__30747;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30724;
    wire N__30723;
    wire N__30722;
    wire N__30721;
    wire N__30720;
    wire N__30719;
    wire N__30716;
    wire N__30715;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30679;
    wire N__30676;
    wire N__30663;
    wire N__30660;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30647;
    wire N__30646;
    wire N__30643;
    wire N__30642;
    wire N__30641;
    wire N__30636;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30592;
    wire N__30589;
    wire N__30584;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30567;
    wire N__30564;
    wire N__30563;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30544;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30511;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30491;
    wire N__30490;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30474;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30452;
    wire N__30451;
    wire N__30450;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30435;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30413;
    wire N__30412;
    wire N__30411;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30396;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30359;
    wire N__30356;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30323;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30273;
    wire N__30270;
    wire N__30269;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30035;
    wire N__30034;
    wire N__30033;
    wire N__30032;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30023;
    wire N__30022;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30008;
    wire N__30007;
    wire N__30006;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29980;
    wire N__29979;
    wire N__29978;
    wire N__29977;
    wire N__29976;
    wire N__29975;
    wire N__29974;
    wire N__29973;
    wire N__29972;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29956;
    wire N__29955;
    wire N__29954;
    wire N__29953;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29930;
    wire N__29929;
    wire N__29928;
    wire N__29927;
    wire N__29926;
    wire N__29925;
    wire N__29924;
    wire N__29923;
    wire N__29908;
    wire N__29905;
    wire N__29894;
    wire N__29887;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29870;
    wire N__29867;
    wire N__29866;
    wire N__29863;
    wire N__29862;
    wire N__29861;
    wire N__29860;
    wire N__29859;
    wire N__29846;
    wire N__29845;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29840;
    wire N__29839;
    wire N__29838;
    wire N__29837;
    wire N__29830;
    wire N__29825;
    wire N__29816;
    wire N__29805;
    wire N__29804;
    wire N__29803;
    wire N__29802;
    wire N__29801;
    wire N__29800;
    wire N__29797;
    wire N__29796;
    wire N__29795;
    wire N__29794;
    wire N__29793;
    wire N__29782;
    wire N__29781;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29777;
    wire N__29776;
    wire N__29775;
    wire N__29774;
    wire N__29771;
    wire N__29770;
    wire N__29769;
    wire N__29768;
    wire N__29767;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29759;
    wire N__29756;
    wire N__29743;
    wire N__29740;
    wire N__29735;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29714;
    wire N__29713;
    wire N__29712;
    wire N__29705;
    wire N__29702;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29697;
    wire N__29694;
    wire N__29685;
    wire N__29676;
    wire N__29671;
    wire N__29660;
    wire N__29657;
    wire N__29656;
    wire N__29655;
    wire N__29654;
    wire N__29653;
    wire N__29652;
    wire N__29651;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29647;
    wire N__29646;
    wire N__29645;
    wire N__29644;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29634;
    wire N__29633;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29627;
    wire N__29626;
    wire N__29625;
    wire N__29624;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29616;
    wire N__29615;
    wire N__29614;
    wire N__29611;
    wire N__29604;
    wire N__29599;
    wire N__29594;
    wire N__29587;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29567;
    wire N__29560;
    wire N__29551;
    wire N__29536;
    wire N__29531;
    wire N__29528;
    wire N__29521;
    wire N__29508;
    wire N__29503;
    wire N__29498;
    wire N__29497;
    wire N__29494;
    wire N__29493;
    wire N__29492;
    wire N__29489;
    wire N__29488;
    wire N__29487;
    wire N__29486;
    wire N__29485;
    wire N__29482;
    wire N__29477;
    wire N__29472;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29452;
    wire N__29447;
    wire N__29444;
    wire N__29437;
    wire N__29428;
    wire N__29425;
    wire N__29414;
    wire N__29409;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29380;
    wire N__29375;
    wire N__29372;
    wire N__29359;
    wire N__29358;
    wire N__29353;
    wire N__29332;
    wire N__29325;
    wire N__29322;
    wire N__29311;
    wire N__29288;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29258;
    wire N__29255;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29238;
    wire N__29235;
    wire N__29230;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29195;
    wire N__29184;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29166;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29096;
    wire N__29093;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29073;
    wire N__29072;
    wire N__29071;
    wire N__29070;
    wire N__29069;
    wire N__29068;
    wire N__29067;
    wire N__29066;
    wire N__29065;
    wire N__29064;
    wire N__29063;
    wire N__29062;
    wire N__29059;
    wire N__29058;
    wire N__29057;
    wire N__29056;
    wire N__29055;
    wire N__29054;
    wire N__29053;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29046;
    wire N__29043;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29020;
    wire N__29019;
    wire N__29016;
    wire N__29015;
    wire N__29014;
    wire N__29013;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28996;
    wire N__28993;
    wire N__28992;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28986;
    wire N__28985;
    wire N__28984;
    wire N__28981;
    wire N__28976;
    wire N__28973;
    wire N__28972;
    wire N__28969;
    wire N__28968;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28958;
    wire N__28957;
    wire N__28954;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28937;
    wire N__28934;
    wire N__28925;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28869;
    wire N__28868;
    wire N__28867;
    wire N__28864;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28856;
    wire N__28855;
    wire N__28854;
    wire N__28853;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28823;
    wire N__28814;
    wire N__28809;
    wire N__28802;
    wire N__28799;
    wire N__28794;
    wire N__28791;
    wire N__28784;
    wire N__28773;
    wire N__28772;
    wire N__28769;
    wire N__28764;
    wire N__28761;
    wire N__28756;
    wire N__28753;
    wire N__28752;
    wire N__28751;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28747;
    wire N__28746;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28742;
    wire N__28739;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28723;
    wire N__28714;
    wire N__28711;
    wire N__28700;
    wire N__28697;
    wire N__28690;
    wire N__28685;
    wire N__28674;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28658;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28647;
    wire N__28644;
    wire N__28643;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28613;
    wire N__28606;
    wire N__28603;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28550;
    wire N__28547;
    wire N__28542;
    wire N__28531;
    wire N__28526;
    wire N__28521;
    wire N__28518;
    wire N__28503;
    wire N__28486;
    wire N__28471;
    wire N__28466;
    wire N__28455;
    wire N__28440;
    wire N__28425;
    wire N__28398;
    wire N__28397;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28353;
    wire N__28344;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28320;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28305;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28248;
    wire N__28245;
    wire N__28244;
    wire N__28241;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28230;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28215;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28157;
    wire N__28156;
    wire N__28153;
    wire N__28152;
    wire N__28151;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28133;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28098;
    wire N__28097;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28043;
    wire N__28042;
    wire N__28041;
    wire N__28038;
    wire N__28033;
    wire N__28030;
    wire N__28023;
    wire N__28020;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27993;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27975;
    wire N__27972;
    wire N__27967;
    wire N__27964;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27932;
    wire N__27931;
    wire N__27930;
    wire N__27927;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27906;
    wire N__27897;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27843;
    wire N__27840;
    wire N__27835;
    wire N__27832;
    wire N__27827;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27791;
    wire N__27788;
    wire N__27787;
    wire N__27786;
    wire N__27785;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27749;
    wire N__27746;
    wire N__27739;
    wire N__27736;
    wire N__27729;
    wire N__27728;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27704;
    wire N__27703;
    wire N__27698;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27679;
    wire N__27672;
    wire N__27671;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27659;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27647;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27635;
    wire N__27630;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27557;
    wire N__27552;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27544;
    wire N__27539;
    wire N__27536;
    wire N__27535;
    wire N__27530;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27519;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27504;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27429;
    wire N__27426;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27405;
    wire N__27400;
    wire N__27397;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27329;
    wire N__27328;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27308;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27290;
    wire N__27285;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27162;
    wire N__27161;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27102;
    wire N__27099;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27081;
    wire N__27078;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27067;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27055;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27034;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27016;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26996;
    wire N__26995;
    wire N__26992;
    wire N__26987;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26943;
    wire N__26942;
    wire N__26939;
    wire N__26938;
    wire N__26935;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26921;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26898;
    wire N__26893;
    wire N__26880;
    wire N__26877;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26816;
    wire N__26815;
    wire N__26814;
    wire N__26813;
    wire N__26810;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26794;
    wire N__26787;
    wire N__26784;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26772;
    wire N__26769;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26739;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26721;
    wire N__26718;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26691;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26685;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26659;
    wire N__26656;
    wire N__26655;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26640;
    wire N__26637;
    wire N__26628;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26620;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26612;
    wire N__26607;
    wire N__26606;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26592;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26541;
    wire N__26536;
    wire N__26533;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26518;
    wire N__26515;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26486;
    wire N__26485;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26473;
    wire N__26466;
    wire N__26463;
    wire N__26462;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26441;
    wire N__26438;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26409;
    wire N__26408;
    wire N__26405;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26381;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26353;
    wire N__26346;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26292;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26212;
    wire N__26207;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26190;
    wire N__26187;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26172;
    wire N__26169;
    wire N__26164;
    wire N__26161;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26132;
    wire N__26127;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26097;
    wire N__26096;
    wire N__26095;
    wire N__26092;
    wire N__26087;
    wire N__26082;
    wire N__26081;
    wire N__26080;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26046;
    wire N__26043;
    wire N__26038;
    wire N__26031;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25977;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25950;
    wire N__25949;
    wire N__25948;
    wire N__25947;
    wire N__25938;
    wire N__25935;
    wire N__25934;
    wire N__25929;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25896;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25882;
    wire N__25875;
    wire N__25874;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25863;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25844;
    wire N__25843;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25831;
    wire N__25824;
    wire N__25823;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25805;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25745;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25729;
    wire N__25722;
    wire N__25719;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25711;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25613;
    wire N__25612;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25604;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25586;
    wire N__25581;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25489;
    wire N__25482;
    wire N__25481;
    wire N__25480;
    wire N__25477;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25454;
    wire N__25445;
    wire N__25442;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25339;
    wire N__25338;
    wire N__25335;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25318;
    wire N__25315;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25303;
    wire N__25300;
    wire N__25295;
    wire N__25290;
    wire N__25287;
    wire N__25278;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25251;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25224;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25170;
    wire N__25167;
    wire N__25166;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25140;
    wire N__25139;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25095;
    wire N__25092;
    wire N__25083;
    wire N__25080;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25023;
    wire N__25020;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24986;
    wire N__24985;
    wire N__24984;
    wire N__24981;
    wire N__24980;
    wire N__24975;
    wire N__24970;
    wire N__24967;
    wire N__24960;
    wire N__24959;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24948;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24918;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24887;
    wire N__24882;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24861;
    wire N__24860;
    wire N__24857;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24820;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24800;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24785;
    wire N__24782;
    wire N__24781;
    wire N__24780;
    wire N__24777;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24756;
    wire N__24755;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24743;
    wire N__24738;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24656;
    wire N__24655;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24618;
    wire N__24615;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24568;
    wire N__24561;
    wire N__24560;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24513;
    wire N__24504;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24466;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24442;
    wire N__24441;
    wire N__24438;
    wire N__24437;
    wire N__24434;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24407;
    wire N__24402;
    wire N__24399;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24391;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24379;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24332;
    wire N__24331;
    wire N__24328;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24313;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24299;
    wire N__24298;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24281;
    wire N__24278;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24242;
    wire N__24241;
    wire N__24240;
    wire N__24237;
    wire N__24230;
    wire N__24225;
    wire N__24224;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24213;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24189;
    wire N__24188;
    wire N__24185;
    wire N__24184;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24158;
    wire N__24155;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24136;
    wire N__24129;
    wire N__24128;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24090;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24082;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24048;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23980;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23944;
    wire N__23943;
    wire N__23938;
    wire N__23933;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23851;
    wire N__23850;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23796;
    wire N__23787;
    wire N__23786;
    wire N__23783;
    wire N__23782;
    wire N__23781;
    wire N__23776;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23748;
    wire N__23745;
    wire N__23740;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23720;
    wire N__23715;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23667;
    wire N__23664;
    wire N__23663;
    wire N__23662;
    wire N__23661;
    wire N__23660;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23640;
    wire N__23635;
    wire N__23630;
    wire N__23623;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23576;
    wire N__23575;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23562;
    wire N__23561;
    wire N__23560;
    wire N__23559;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23552;
    wire N__23551;
    wire N__23550;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23540;
    wire N__23537;
    wire N__23528;
    wire N__23527;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23521;
    wire N__23520;
    wire N__23517;
    wire N__23516;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23494;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23481;
    wire N__23480;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23471;
    wire N__23470;
    wire N__23469;
    wire N__23468;
    wire N__23465;
    wire N__23460;
    wire N__23457;
    wire N__23452;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23438;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23424;
    wire N__23421;
    wire N__23420;
    wire N__23419;
    wire N__23418;
    wire N__23415;
    wire N__23410;
    wire N__23403;
    wire N__23402;
    wire N__23401;
    wire N__23400;
    wire N__23397;
    wire N__23386;
    wire N__23383;
    wire N__23372;
    wire N__23361;
    wire N__23350;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23332;
    wire N__23327;
    wire N__23326;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23308;
    wire N__23301;
    wire N__23294;
    wire N__23291;
    wire N__23286;
    wire N__23275;
    wire N__23268;
    wire N__23267;
    wire N__23266;
    wire N__23263;
    wire N__23262;
    wire N__23259;
    wire N__23248;
    wire N__23241;
    wire N__23234;
    wire N__23229;
    wire N__23224;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23189;
    wire N__23184;
    wire N__23181;
    wire N__23180;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23154;
    wire N__23153;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23114;
    wire N__23109;
    wire N__23106;
    wire N__23105;
    wire N__23100;
    wire N__23097;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23067;
    wire N__23066;
    wire N__23061;
    wire N__23058;
    wire N__23057;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23016;
    wire N__23013;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22995;
    wire N__22992;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22984;
    wire N__22983;
    wire N__22978;
    wire N__22977;
    wire N__22976;
    wire N__22973;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22957;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22848;
    wire N__22845;
    wire N__22844;
    wire N__22839;
    wire N__22836;
    wire N__22835;
    wire N__22830;
    wire N__22827;
    wire N__22826;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22805;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22779;
    wire N__22778;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22760;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22715;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22693;
    wire N__22686;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22675;
    wire N__22674;
    wire N__22673;
    wire N__22672;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22575;
    wire N__22574;
    wire N__22571;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22559;
    wire N__22554;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22536;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22524;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22502;
    wire N__22499;
    wire N__22494;
    wire N__22489;
    wire N__22484;
    wire N__22479;
    wire N__22476;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22468;
    wire N__22467;
    wire N__22464;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22443;
    wire N__22438;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22411;
    wire N__22408;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22383;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22332;
    wire N__22329;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22305;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22284;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22227;
    wire N__22224;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22209;
    wire N__22208;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22196;
    wire N__22191;
    wire N__22186;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22157;
    wire N__22152;
    wire N__22151;
    wire N__22148;
    wire N__22147;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22135;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22058;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22039;
    wire N__22036;
    wire N__22031;
    wire N__22028;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21973;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21903;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21844;
    wire N__21837;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21794;
    wire N__21793;
    wire N__21788;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21766;
    wire N__21763;
    wire N__21758;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21731;
    wire N__21730;
    wire N__21727;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21698;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21647;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21627;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21603;
    wire N__21598;
    wire N__21591;
    wire N__21590;
    wire N__21585;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21538;
    wire N__21537;
    wire N__21532;
    wire N__21529;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21486;
    wire N__21483;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21375;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21337;
    wire N__21330;
    wire N__21327;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21234;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21192;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21168;
    wire N__21165;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21150;
    wire N__21145;
    wire N__21144;
    wire N__21141;
    wire N__21136;
    wire N__21133;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21075;
    wire N__21072;
    wire N__21067;
    wire N__21064;
    wire N__21063;
    wire N__21060;
    wire N__21055;
    wire N__21052;
    wire N__21045;
    wire N__21044;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21023;
    wire N__21020;
    wire N__21019;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__20997;
    wire N__20994;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20982;
    wire N__20979;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20892;
    wire N__20889;
    wire N__20880;
    wire N__20879;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20776;
    wire N__20775;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20760;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20719;
    wire N__20718;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20700;
    wire N__20697;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20672;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20630;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20593;
    wire N__20590;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20515;
    wire N__20510;
    wire N__20505;
    wire N__20502;
    wire N__20501;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20475;
    wire N__20474;
    wire N__20473;
    wire N__20468;
    wire N__20465;
    wire N__20460;
    wire N__20457;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20441;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20397;
    wire N__20396;
    wire N__20391;
    wire N__20388;
    wire N__20387;
    wire N__20382;
    wire N__20379;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20367;
    wire N__20366;
    wire N__20365;
    wire N__20362;
    wire N__20357;
    wire N__20352;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20337;
    wire N__20336;
    wire N__20335;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20271;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20259;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20247;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20208;
    wire N__20207;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20178;
    wire N__20175;
    wire N__20174;
    wire N__20169;
    wire N__20166;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20154;
    wire N__20153;
    wire N__20148;
    wire N__20145;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20115;
    wire N__20114;
    wire N__20109;
    wire N__20106;
    wire N__20105;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20093;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20070;
    wire N__20067;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19983;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19962;
    wire N__19961;
    wire N__19956;
    wire N__19953;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19941;
    wire N__19940;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19910;
    wire N__19907;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19887;
    wire N__19886;
    wire N__19883;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19875;
    wire N__19872;
    wire N__19867;
    wire N__19864;
    wire N__19857;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19818;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19800;
    wire N__19795;
    wire N__19790;
    wire N__19787;
    wire N__19782;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19771;
    wire N__19770;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19747;
    wire N__19744;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19715;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19686;
    wire N__19685;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19677;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19650;
    wire N__19645;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19611;
    wire N__19610;
    wire N__19607;
    wire N__19602;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19539;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19489;
    wire N__19486;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19462;
    wire N__19459;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19424;
    wire N__19421;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19354;
    wire N__19353;
    wire N__19352;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19304;
    wire N__19303;
    wire N__19300;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19273;
    wire N__19272;
    wire N__19265;
    wire N__19262;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19185;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19168;
    wire N__19165;
    wire N__19158;
    wire N__19155;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19148;
    wire N__19147;
    wire N__19146;
    wire N__19143;
    wire N__19138;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19129;
    wire N__19128;
    wire N__19127;
    wire N__19126;
    wire N__19125;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19119;
    wire N__19118;
    wire N__19117;
    wire N__19114;
    wire N__19113;
    wire N__19112;
    wire N__19109;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19089;
    wire N__19088;
    wire N__19087;
    wire N__19086;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19067;
    wire N__19066;
    wire N__19065;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19056;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19041;
    wire N__19040;
    wire N__19039;
    wire N__19036;
    wire N__19027;
    wire N__19020;
    wire N__19017;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__18992;
    wire N__18987;
    wire N__18982;
    wire N__18971;
    wire N__18964;
    wire N__18959;
    wire N__18956;
    wire N__18949;
    wire N__18934;
    wire N__18923;
    wire N__18912;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18896;
    wire N__18889;
    wire N__18858;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18850;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18762;
    wire N__18759;
    wire N__18758;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18729;
    wire N__18720;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18712;
    wire N__18711;
    wire N__18708;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18681;
    wire N__18678;
    wire N__18677;
    wire N__18676;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18642;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18636;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18617;
    wire N__18606;
    wire N__18603;
    wire N__18602;
    wire N__18601;
    wire N__18598;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18582;
    wire N__18579;
    wire N__18578;
    wire N__18577;
    wire N__18574;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18552;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18519;
    wire N__18516;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18508;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18483;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18471;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18393;
    wire N__18392;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18380;
    wire N__18379;
    wire N__18376;
    wire N__18375;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18354;
    wire N__18353;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18341;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18312;
    wire N__18311;
    wire N__18310;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18290;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18270;
    wire N__18269;
    wire N__18268;
    wire N__18261;
    wire N__18258;
    wire N__18257;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18243;
    wire N__18240;
    wire N__18239;
    wire N__18234;
    wire N__18231;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18219;
    wire N__18218;
    wire N__18213;
    wire N__18210;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18198;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18186;
    wire N__18185;
    wire N__18180;
    wire N__18177;
    wire N__18176;
    wire N__18171;
    wire N__18168;
    wire N__18167;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18144;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18129;
    wire N__18126;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18058;
    wire N__18057;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18029;
    wire N__18024;
    wire N__18021;
    wire N__18020;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17955;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17944;
    wire N__17943;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17928;
    wire N__17925;
    wire N__17922;
    wire N__17913;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17898;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17757;
    wire N__17756;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17741;
    wire N__17736;
    wire N__17733;
    wire N__17732;
    wire N__17729;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17714;
    wire N__17709;
    wire N__17706;
    wire N__17705;
    wire N__17704;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17692;
    wire N__17687;
    wire N__17682;
    wire N__17679;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17604;
    wire N__17603;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17595;
    wire N__17594;
    wire N__17593;
    wire N__17590;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17563;
    wire N__17550;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17542;
    wire N__17541;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17514;
    wire N__17511;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17479;
    wire N__17472;
    wire N__17469;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17450;
    wire N__17447;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17436;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17413;
    wire N__17406;
    wire N__17403;
    wire N__17402;
    wire N__17399;
    wire N__17398;
    wire N__17395;
    wire N__17394;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17358;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17274;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17126;
    wire N__17125;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17113;
    wire N__17110;
    wire N__17103;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17094;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17073;
    wire N__17070;
    wire N__17069;
    wire N__17068;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17046;
    wire N__17043;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16995;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16971;
    wire N__16968;
    wire N__16963;
    wire N__16960;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16942;
    wire N__16937;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16884;
    wire N__16883;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16848;
    wire N__16847;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16818;
    wire N__16817;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16806;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16738;
    wire N__16735;
    wire N__16728;
    wire N__16725;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16698;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16686;
    wire N__16683;
    wire N__16680;
    wire N__16677;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16646;
    wire N__16643;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16616;
    wire N__16615;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16603;
    wire N__16596;
    wire N__16595;
    wire N__16594;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16566;
    wire N__16563;
    wire N__16562;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16544;
    wire N__16543;
    wire N__16542;
    wire N__16539;
    wire N__16534;
    wire N__16531;
    wire N__16524;
    wire N__16521;
    wire N__16520;
    wire N__16519;
    wire N__16518;
    wire N__16515;
    wire N__16508;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16473;
    wire N__16464;
    wire N__16461;
    wire N__16460;
    wire N__16459;
    wire N__16458;
    wire N__16451;
    wire N__16448;
    wire N__16443;
    wire N__16440;
    wire N__16439;
    wire N__16436;
    wire N__16435;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16413;
    wire N__16412;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16390;
    wire N__16383;
    wire N__16380;
    wire N__16379;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16347;
    wire N__16344;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16317;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16305;
    wire N__16304;
    wire N__16299;
    wire N__16296;
    wire N__16295;
    wire N__16290;
    wire N__16287;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16275;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16263;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16224;
    wire N__16221;
    wire N__16220;
    wire N__16219;
    wire N__16216;
    wire N__16211;
    wire N__16208;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16196;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16179;
    wire N__16178;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16171;
    wire N__16166;
    wire N__16163;
    wire N__16158;
    wire N__16155;
    wire N__16146;
    wire N__16145;
    wire N__16144;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16128;
    wire N__16127;
    wire N__16122;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16110;
    wire N__16109;
    wire N__16108;
    wire N__16107;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16082;
    wire N__16075;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16050;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16005;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15993;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15981;
    wire N__15980;
    wire N__15975;
    wire N__15972;
    wire N__15971;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15943;
    wire N__15942;
    wire N__15941;
    wire N__15940;
    wire N__15939;
    wire N__15938;
    wire N__15937;
    wire N__15934;
    wire N__15925;
    wire N__15922;
    wire N__15915;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15878;
    wire N__15873;
    wire N__15872;
    wire N__15871;
    wire N__15870;
    wire N__15869;
    wire N__15866;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15846;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15838;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15823;
    wire N__15818;
    wire N__15815;
    wire N__15810;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15769;
    wire N__15764;
    wire N__15761;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15668;
    wire N__15667;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15655;
    wire N__15652;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15625;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15613;
    wire N__15606;
    wire N__15605;
    wire N__15604;
    wire N__15599;
    wire N__15596;
    wire N__15595;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15575;
    wire N__15570;
    wire N__15569;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15550;
    wire N__15547;
    wire N__15542;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15444;
    wire N__15441;
    wire N__15440;
    wire N__15437;
    wire N__15436;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15421;
    wire N__15416;
    wire N__15415;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15403;
    wire N__15400;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15375;
    wire N__15372;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15293;
    wire N__15292;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15244;
    wire N__15239;
    wire N__15236;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15215;
    wire N__15212;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15101;
    wire N__15100;
    wire N__15097;
    wire N__15092;
    wire N__15087;
    wire N__15086;
    wire N__15085;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15064;
    wire N__15063;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15026;
    wire N__15023;
    wire N__15022;
    wire N__15019;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__14997;
    wire N__14994;
    wire N__14993;
    wire N__14990;
    wire N__14989;
    wire N__14986;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14965;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14942;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14913;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14898;
    wire N__14897;
    wire N__14894;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14861;
    wire N__14858;
    wire N__14857;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14835;
    wire N__14832;
    wire N__14831;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14796;
    wire N__14793;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14781;
    wire N__14778;
    wire N__14777;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14709;
    wire N__14706;
    wire N__14705;
    wire N__14704;
    wire N__14701;
    wire N__14696;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14681;
    wire N__14680;
    wire N__14679;
    wire N__14676;
    wire N__14669;
    wire N__14664;
    wire N__14661;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14653;
    wire N__14652;
    wire N__14649;
    wire N__14642;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14613;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14601;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14589;
    wire N__14588;
    wire N__14585;
    wire N__14584;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14566;
    wire N__14563;
    wire N__14556;
    wire N__14555;
    wire N__14552;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14504;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14481;
    wire N__14480;
    wire N__14475;
    wire N__14472;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14460;
    wire N__14459;
    wire N__14454;
    wire N__14451;
    wire N__14450;
    wire N__14445;
    wire N__14442;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14430;
    wire N__14429;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14417;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14388;
    wire N__14385;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14349;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14333;
    wire N__14332;
    wire N__14327;
    wire N__14324;
    wire N__14319;
    wire N__14318;
    wire N__14317;
    wire N__14316;
    wire N__14315;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14304;
    wire N__14301;
    wire N__14300;
    wire N__14299;
    wire N__14292;
    wire N__14289;
    wire N__14284;
    wire N__14277;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14261;
    wire N__14252;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14233;
    wire N__14230;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14177;
    wire N__14176;
    wire N__14173;
    wire N__14168;
    wire N__14163;
    wire N__14160;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14145;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14003;
    wire N__14000;
    wire N__13999;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13980;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13972;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13960;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13938;
    wire N__13935;
    wire N__13934;
    wire N__13933;
    wire N__13932;
    wire N__13931;
    wire N__13928;
    wire N__13921;
    wire N__13918;
    wire N__13913;
    wire N__13908;
    wire N__13905;
    wire N__13904;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13881;
    wire N__13878;
    wire N__13877;
    wire N__13876;
    wire N__13873;
    wire N__13868;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13838;
    wire N__13837;
    wire N__13836;
    wire N__13833;
    wire N__13828;
    wire N__13825;
    wire N__13818;
    wire N__13817;
    wire N__13814;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13797;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13777;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13753;
    wire N__13752;
    wire N__13749;
    wire N__13742;
    wire N__13737;
    wire N__13734;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13648;
    wire N__13643;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13624;
    wire N__13619;
    wire N__13616;
    wire N__13611;
    wire N__13610;
    wire N__13607;
    wire N__13606;
    wire N__13605;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13591;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13565;
    wire N__13562;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13554;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13540;
    wire N__13533;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13521;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13509;
    wire N__13508;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13496;
    wire N__13493;
    wire N__13492;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13477;
    wire N__13470;
    wire N__13467;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13398;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13374;
    wire N__13373;
    wire N__13368;
    wire N__13365;
    wire N__13364;
    wire N__13359;
    wire N__13356;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13290;
    wire N__13287;
    wire N__13286;
    wire N__13285;
    wire N__13284;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13270;
    wire N__13263;
    wire N__13262;
    wire N__13261;
    wire N__13260;
    wire N__13253;
    wire N__13250;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13195;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13155;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13143;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13128;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13116;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13073;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12951;
    wire N__12948;
    wire N__12941;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12850;
    wire N__12847;
    wire N__12840;
    wire N__12839;
    wire N__12834;
    wire N__12831;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12819;
    wire N__12818;
    wire N__12813;
    wire N__12810;
    wire N__12809;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12773;
    wire N__12768;
    wire N__12765;
    wire N__12764;
    wire N__12759;
    wire N__12756;
    wire N__12755;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12563;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12536;
    wire N__12535;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12520;
    wire N__12515;
    wire N__12510;
    wire N__12509;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12486;
    wire N__12485;
    wire N__12480;
    wire N__12477;
    wire N__12476;
    wire N__12471;
    wire N__12468;
    wire N__12467;
    wire N__12462;
    wire N__12459;
    wire N__12458;
    wire N__12453;
    wire N__12450;
    wire N__12449;
    wire N__12444;
    wire N__12441;
    wire N__12440;
    wire N__12435;
    wire N__12432;
    wire N__12431;
    wire N__12426;
    wire N__12423;
    wire N__12422;
    wire N__12417;
    wire N__12414;
    wire N__12413;
    wire N__12408;
    wire N__12405;
    wire N__12404;
    wire N__12399;
    wire N__12396;
    wire N__12395;
    wire N__12390;
    wire N__12387;
    wire N__12386;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire data_in_10_1;
    wire data_in_11_1;
    wire data_in_14_1;
    wire data_in_13_1;
    wire data_in_12_1;
    wire data_in_7_4;
    wire data_in_8_4;
    wire data_in_9_4;
    wire data_in_10_4;
    wire data_in_11_4;
    wire data_in_12_4;
    wire data_in_5_1;
    wire data_in_6_1;
    wire data_in_7_1;
    wire data_in_9_1;
    wire data_in_8_1;
    wire \c0.n4431_cascade_ ;
    wire n1902;
    wire data_in_6_4;
    wire \c0.n24_cascade_ ;
    wire \c0.n4_adj_1594_cascade_ ;
    wire \c0.n9674_cascade_ ;
    wire \c0.n9677_cascade_ ;
    wire \c0.n4431 ;
    wire \c0.n8849_cascade_ ;
    wire \c0.n20_adj_1622_cascade_ ;
    wire \c0.data_in_frame_19_5 ;
    wire \c0.n10_adj_1637_cascade_ ;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n9686_cascade_ ;
    wire \c0.n9689_cascade_ ;
    wire \c0.n10_adj_1646 ;
    wire \c0.n8779 ;
    wire \c0.n54_cascade_ ;
    wire \c0.n49 ;
    wire \c0.n9001 ;
    wire \c0.n9001_cascade_ ;
    wire \c0.n9464_cascade_ ;
    wire \c0.n9470_cascade_ ;
    wire \c0.n9216 ;
    wire \c0.n9213_cascade_ ;
    wire \c0.n9210 ;
    wire \c0.n9458_cascade_ ;
    wire \c0.n9461_cascade_ ;
    wire \c0.n9530_cascade_ ;
    wire \c0.n9524_cascade_ ;
    wire \c0.n9183 ;
    wire \c0.n9186_cascade_ ;
    wire \c0.n9518_cascade_ ;
    wire \c0.n22_adj_1680 ;
    wire \c0.n9521_cascade_ ;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire bfn_1_31_0_;
    wire \c0.tx2.n8105 ;
    wire \c0.tx2.n8106 ;
    wire \c0.tx2.n8107 ;
    wire \c0.tx2.n8108 ;
    wire \c0.tx2.n8109 ;
    wire \c0.tx2.n8110 ;
    wire \c0.tx2.n8111 ;
    wire \c0.tx2.n8112 ;
    wire bfn_1_32_0_;
    wire data_in_7_7;
    wire data_in_10_7;
    wire data_in_11_7;
    wire data_in_12_7;
    wire data_in_13_4;
    wire data_in_14_4;
    wire data_in_10_0;
    wire data_in_11_0;
    wire \c0.n9548_cascade_ ;
    wire \c0.n9177 ;
    wire \c0.data_in_field_10 ;
    wire \c0.n8801_cascade_ ;
    wire \c0.data_in_field_11 ;
    wire \c0.n4276 ;
    wire \c0.n4276_cascade_ ;
    wire \c0.n12_adj_1633_cascade_ ;
    wire \c0.n4327 ;
    wire \c0.n4434_cascade_ ;
    wire \c0.n8766 ;
    wire \c0.n9482_cascade_ ;
    wire \c0.n9207 ;
    wire n1894;
    wire \c0.n9542_cascade_ ;
    wire \c0.n9180 ;
    wire \c0.n4114_cascade_ ;
    wire \c0.n17_cascade_ ;
    wire \c0.n4324_cascade_ ;
    wire \c0.n8951 ;
    wire \c0.n8951_cascade_ ;
    wire \c0.n48 ;
    wire \c0.n4406 ;
    wire \c0.n4406_cascade_ ;
    wire \c0.n43_adj_1610 ;
    wire \c0.data_in_frame_20_5 ;
    wire \c0.n4215_cascade_ ;
    wire \c0.n18_adj_1593_cascade_ ;
    wire \c0.n20_adj_1596 ;
    wire \c0.n4568_cascade_ ;
    wire \c0.n46 ;
    wire data_in_6_7;
    wire \c0.n8816 ;
    wire \c0.n4282_cascade_ ;
    wire \c0.n4577 ;
    wire \c0.n4282 ;
    wire \c0.n4476_cascade_ ;
    wire \c0.n19_adj_1623 ;
    wire data_in_5_7;
    wire tx2_enable;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire \c0.tx2.n5_cascade_ ;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire \c0.tx2.n4081 ;
    wire \c0.tx2.n4081_cascade_ ;
    wire \c0.tx2.n7 ;
    wire \c0.tx2.n8196_cascade_ ;
    wire \c0.tx2.n5146 ;
    wire n9075_cascade_;
    wire \c0.tx2.r_Clock_Count_8 ;
    wire \c0.tx2.n7399 ;
    wire \c0.tx2.n7236 ;
    wire \c0.tx2.n7236_cascade_ ;
    wire n3220_cascade_;
    wire data_in_9_7;
    wire data_in_8_7;
    wire n1900;
    wire data_in_7_3;
    wire data_in_8_3;
    wire data_in_9_0;
    wire data_in_8_0;
    wire data_in_7_0;
    wire data_in_1_5;
    wire data_in_12_0;
    wire \c0.n14_adj_1670 ;
    wire \c0.n14_adj_1669 ;
    wire \c0.n26_adj_1673 ;
    wire \c0.n25_adj_1675 ;
    wire \c0.n9033_cascade_ ;
    wire \c0.n9578 ;
    wire \c0.n8794 ;
    wire data_in_3_1;
    wire data_in_0_2;
    wire \c0.n4381 ;
    wire \c0.n4381_cascade_ ;
    wire \c0.data_in_field_20 ;
    wire data_in_4_1;
    wire \c0.data_in_field_35 ;
    wire \c0.n4154_cascade_ ;
    wire \c0.data_in_field_19 ;
    wire \c0.n14 ;
    wire \c0.n10_adj_1631_cascade_ ;
    wire data_in_1_1;
    wire data_in_4_7;
    wire \c0.n47 ;
    wire \c0.data_in_field_4 ;
    wire data_in_0_7;
    wire \c0.n8776 ;
    wire \c0.n4131_cascade_ ;
    wire \c0.n8927_cascade_ ;
    wire n1896;
    wire data_in_2_7;
    wire data_in_0_6;
    wire \c0.n10_adj_1647_cascade_ ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.n9704_cascade_ ;
    wire \c0.data_in_frame_20_1 ;
    wire \c0.n9707_cascade_ ;
    wire \c0.n22_adj_1682 ;
    wire \c0.n9722_cascade_ ;
    wire \c0.data_in_field_7 ;
    wire \c0.data_in_field_23 ;
    wire \c0.n4514 ;
    wire \c0.n9007 ;
    wire \c0.n18_adj_1589_cascade_ ;
    wire \c0.n20_adj_1590_cascade_ ;
    wire \c0.n29 ;
    wire \c0.n4114 ;
    wire \c0.n4448 ;
    wire \c0.n4445 ;
    wire \c0.n8896 ;
    wire n6164;
    wire data_in_field_105;
    wire \c0.n8890_cascade_ ;
    wire \c0.n14_adj_1638 ;
    wire \c0.n4285 ;
    wire data_in_field_83;
    wire \c0.n9126 ;
    wire \c0.n9123_cascade_ ;
    wire \c0.n9240 ;
    wire \c0.n9644_cascade_ ;
    wire \c0.n9647_cascade_ ;
    wire \c0.n9656 ;
    wire \c0.n9752_cascade_ ;
    wire \c0.data_in_field_39 ;
    wire \c0.n9120 ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.n9692_cascade_ ;
    wire \c0.tx2.n9695_cascade_ ;
    wire \c0.tx2.o_Tx_Serial_N_1511_cascade_ ;
    wire n2207_cascade_;
    wire r_Bit_Index_2_adj_1741;
    wire r_SM_Main_0_adj_1740;
    wire r_SM_Main_2_N_1480_1_adj_1744;
    wire data_in_13_7;
    wire data_in_16_6;
    wire data_in_9_6;
    wire data_in_10_6;
    wire data_in_11_6;
    wire data_in_13_6;
    wire data_in_12_6;
    wire data_in_15_6;
    wire data_in_14_6;
    wire data_in_20_4;
    wire data_in_3_0;
    wire data_in_0_5;
    wire \c0.n28_adj_1668_cascade_ ;
    wire \c0.n30_adj_1674 ;
    wire \c0.n22_adj_1667 ;
    wire data_in_0_0;
    wire data_in_13_0;
    wire data_in_4_0;
    wire \c0.n13_adj_1671 ;
    wire \c0.n13_adj_1672 ;
    wire data_in_1_2;
    wire data_in_6_3;
    wire data_in_1_3;
    wire data_in_2_3;
    wire \c0.n4495 ;
    wire \c0.data_in_field_2 ;
    wire \c0.data_in_field_33 ;
    wire \c0.n6_adj_1632_cascade_ ;
    wire \c0.n8804 ;
    wire data_in_1_6;
    wire data_in_3_7;
    wire \c0.n4127 ;
    wire data_in_0_3;
    wire \c0.data_in_field_3 ;
    wire \c0.n20_adj_1597 ;
    wire \c0.n22_adj_1595 ;
    wire data_in_2_6;
    wire n9069_cascade_;
    wire data_in_3_3;
    wire \c0.n8849 ;
    wire n4_adj_1750_cascade_;
    wire n1892;
    wire n1891;
    wire \c0.n8831 ;
    wire \c0.data_in_field_9 ;
    wire \c0.n8831_cascade_ ;
    wire data_in_1_0;
    wire n1888;
    wire data_in_5_3;
    wire data_in_4_3;
    wire \c0.n4131 ;
    wire \c0.n4224 ;
    wire \c0.n10_adj_1640_cascade_ ;
    wire \c0.n4434 ;
    wire \c0.n8933_cascade_ ;
    wire \c0.n8822 ;
    wire \c0.n8314_cascade_ ;
    wire data_in_field_145;
    wire \c0.n4556 ;
    wire \c0.n8861 ;
    wire \c0.n6 ;
    wire \c0.n4452_cascade_ ;
    wire \c0.n8906 ;
    wire \c0.n4452 ;
    wire \c0.n4253_cascade_ ;
    wire data_in_field_71;
    wire data_in_field_147;
    wire data_in_field_127;
    wire \c0.n9650 ;
    wire \c0.n16_adj_1598 ;
    wire \c0.n9016 ;
    wire \c0.n6_adj_1645_cascade_ ;
    wire \c0.n4154 ;
    wire \c0.n8788_cascade_ ;
    wire \c0.n14_adj_1648 ;
    wire \c0.n8936 ;
    wire \c0.n24_adj_1600_cascade_ ;
    wire \c0.n18_adj_1603 ;
    wire \c0.n4107 ;
    wire \c0.tx2_transmit_N_1334_cascade_ ;
    wire \c0.n8980 ;
    wire \c0.n22_adj_1601_cascade_ ;
    wire \c0.n26 ;
    wire \c0.n16 ;
    wire data_in_field_115;
    wire \c0.n4574_cascade_ ;
    wire data_in_field_81;
    wire data_in_field_47;
    wire \c0.n4333 ;
    wire \c0.n4333_cascade_ ;
    wire n3_adj_1749;
    wire tx2_o;
    wire \c0.n24_adj_1615 ;
    wire \c0.n34 ;
    wire r_SM_Main_1_adj_1739;
    wire n8747;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire \c0.tx2.n9716_cascade_ ;
    wire \c0.tx2.n9719 ;
    wire n4691_cascade_;
    wire r_Bit_Index_0_adj_1743;
    wire n9075;
    wire n5346;
    wire r_Bit_Index_1_adj_1742;
    wire data_in_15_1;
    wire data_in_5_4;
    wire data_in_17_1;
    wire data_in_16_1;
    wire data_in_14_7;
    wire data_in_15_7;
    wire data_in_16_7;
    wire data_in_15_4;
    wire data_in_17_4;
    wire data_in_16_4;
    wire data_in_17_7;
    wire data_in_19_4;
    wire data_in_18_4;
    wire data_in_2_5;
    wire data_in_5_6;
    wire data_in_4_6;
    wire data_in_6_6;
    wire data_in_8_6;
    wire data_in_7_6;
    wire data_in_3_5;
    wire data_in_3_6;
    wire \c0.n8843_cascade_ ;
    wire \c0.data_in_field_31 ;
    wire \c0.n4151_cascade_ ;
    wire \c0.data_in_field_30 ;
    wire \c0.data_in_field_22 ;
    wire \c0.data_in_field_14 ;
    wire \c0.n9638_cascade_ ;
    wire \c0.data_in_field_6 ;
    wire data_in_2_0;
    wire \c0.data_in_field_26 ;
    wire \c0.data_in_field_18 ;
    wire \c0.n9512 ;
    wire data_in_2_1;
    wire \c0.n4492 ;
    wire \c0.n24 ;
    wire \c0.n8902 ;
    wire \c0.n4492_cascade_ ;
    wire \c0.n8948_cascade_ ;
    wire \c0.n8858 ;
    wire \c0.n19_adj_1602 ;
    wire data_in_0_1;
    wire \c0.data_in_field_1 ;
    wire data_in_1_7;
    wire \c0.data_in_field_15 ;
    wire n1895_cascade_;
    wire n1889;
    wire n1897;
    wire data_in_4_4;
    wire \c0.n9506_cascade_ ;
    wire \c0.data_in_field_34 ;
    wire \c0.n4_adj_1592_cascade_ ;
    wire \c0.n4324 ;
    wire \c0.n21_adj_1599 ;
    wire \c0.n4200 ;
    wire \c0.n28 ;
    wire \c0.n23_adj_1608 ;
    wire \c0.n8864 ;
    wire \c0.n8843 ;
    wire \c0.n8930 ;
    wire \c0.n20 ;
    wire \c0.n21_cascade_ ;
    wire \c0.n19 ;
    wire \c0.n18 ;
    wire \c0.n8421_cascade_ ;
    wire \c0.tx2_transmit_N_1334 ;
    wire \c0.n24_adj_1605 ;
    wire data_in_field_75;
    wire data_in_field_67;
    wire \c0.n6_adj_1654 ;
    wire \c0.n4253 ;
    wire \c0.n4151 ;
    wire \c0.data_in_field_17 ;
    wire \c0.n45 ;
    wire \c0.n4183 ;
    wire data_in_field_63;
    wire data_in_field_59;
    wire data_in_field_51;
    wire \c0.n4302 ;
    wire data_in_field_79;
    wire data_in_field_139;
    wire \c0.n8825 ;
    wire data_in_field_111;
    wire \c0.n4525_cascade_ ;
    wire data_in_field_107;
    wire data_in_field_137;
    wire \c0.n8874_cascade_ ;
    wire data_in_field_55;
    wire \c0.n6_adj_1636 ;
    wire \c0.n8989 ;
    wire \c0.n6_adj_1604_cascade_ ;
    wire \c0.n8983 ;
    wire \c0.n8948 ;
    wire \c0.n8945 ;
    wire \c0.n8983_cascade_ ;
    wire \c0.n9004 ;
    wire data_in_field_89;
    wire \c0.n4203 ;
    wire \c0.n8890 ;
    wire \c0.n8874 ;
    wire \c0.n24_adj_1607 ;
    wire \c0.n23 ;
    wire \c0.n25_cascade_ ;
    wire \c0.n26_adj_1606 ;
    wire \c0.data_in_frame_20_3 ;
    wire \c0.n8974 ;
    wire \c0.n22_adj_1617 ;
    wire \c0.n8933 ;
    wire \c0.data_in_frame_20_7 ;
    wire \c0.n3056_cascade_ ;
    wire \c0.n22_adj_1676 ;
    wire \c0.n38_adj_1616 ;
    wire \c0.n36 ;
    wire \c0.n37 ;
    wire \c0.data_in_frame_19_7 ;
    wire data_in_field_135;
    wire \c0.n9662_cascade_ ;
    wire \c0.n9665 ;
    wire data_in_13_3;
    wire data_in_14_3;
    wire data_in_16_3;
    wire data_in_15_3;
    wire data_in_17_3;
    wire data_in_18_3;
    wire data_in_19_3;
    wire data_in_20_3;
    wire data_in_19_5;
    wire data_in_17_6;
    wire data_in_10_3;
    wire data_in_9_3;
    wire data_in_20_5;
    wire data_in_5_5;
    wire data_in_4_5;
    wire data_in_6_5;
    wire data_in_7_5;
    wire data_in_8_5;
    wire data_in_9_5;
    wire data_in_14_0;
    wire data_in_15_0;
    wire data_in_2_2;
    wire data_in_16_0;
    wire data_in_20_0;
    wire n1898;
    wire \c0.n9746_cascade_ ;
    wire \c0.data_in_field_32 ;
    wire data_in_field_42;
    wire data_in_field_40;
    wire \c0.n4208 ;
    wire data_in_3_4;
    wire data_in_3_2;
    wire data_in_2_4;
    wire data_in_17_0;
    wire \c0.n8960 ;
    wire data_in_0_4;
    wire n1890;
    wire data_in_1_4;
    wire n9069;
    wire data_in_field_45;
    wire \c0.n9602 ;
    wire \c0.data_in_field_12 ;
    wire \c0.n9019 ;
    wire \c0.data_in_field_28 ;
    wire n9091;
    wire n9092_cascade_;
    wire LED_c;
    wire n8761;
    wire data_in_field_48;
    wire \c0.n4897_cascade_ ;
    wire bfn_6_27_0_;
    wire n8155;
    wire n8156;
    wire n8157;
    wire n8158;
    wire rand_data_5;
    wire n8159;
    wire n8160;
    wire n8161;
    wire n8162;
    wire bfn_6_28_0_;
    wire n8163;
    wire n8164;
    wire n8165;
    wire n8166;
    wire n8167;
    wire rand_data_14;
    wire n8168;
    wire n8169;
    wire n8170;
    wire bfn_6_29_0_;
    wire n8171;
    wire n8172;
    wire rand_data_19;
    wire n8173;
    wire n8174;
    wire n8175;
    wire n8176;
    wire n8177;
    wire n8178;
    wire bfn_6_30_0_;
    wire rand_data_25;
    wire n8179;
    wire n8180;
    wire rand_data_27;
    wire n8181;
    wire n8182;
    wire n8183;
    wire n8184;
    wire n8185;
    wire rand_data_31;
    wire data_in_field_104;
    wire \c0.n9734_cascade_ ;
    wire data_in_field_141;
    wire rand_data_21;
    wire rand_data_17;
    wire data_in_field_113;
    wire data_in_field_149;
    wire \c0.n1893_adj_1635 ;
    wire rand_data_23;
    wire data_in_field_85;
    wire \c0.n9596_cascade_ ;
    wire data_in_field_117;
    wire \c0.n9590_cascade_ ;
    wire \c0.n9153 ;
    wire \c0.n9156_cascade_ ;
    wire \c0.n9584_cascade_ ;
    wire \c0.n9150 ;
    wire \c0.n22_adj_1678 ;
    wire \c0.n9587_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire data_in_10_5;
    wire data_in_11_5;
    wire data_in_13_5;
    wire data_in_12_5;
    wire data_in_14_5;
    wire data_in_15_5;
    wire data_in_16_5;
    wire data_in_18_5;
    wire data_in_17_5;
    wire data_in_18_6;
    wire data_in_18_1;
    wire data_in_19_1;
    wire data_in_20_1;
    wire rx_data_2;
    wire data_in_12_3;
    wire data_in_11_3;
    wire n4;
    wire rx_data_3;
    wire data_in_19_6;
    wire rx_data_0;
    wire data_in_18_7;
    wire data_in_20_6;
    wire n4_adj_1725;
    wire n4_adj_1725_cascade_;
    wire rx_data_1;
    wire n4044_cascade_;
    wire rx_data_6;
    wire rx_data_4;
    wire rx_data_7;
    wire data_in_20_7;
    wire data_in_19_7;
    wire n4044;
    wire rx_data_5;
    wire n4049;
    wire \c0.n9476 ;
    wire rand_data_24;
    wire n1903;
    wire data_in_field_129;
    wire \c0.n8791 ;
    wire data_in_6_0;
    wire data_in_5_0;
    wire \c0.n19_adj_1665_cascade_ ;
    wire tx2_active;
    wire \c0.r_SM_Main_2_N_1483_0 ;
    wire \c0.n19_adj_1665 ;
    wire \c0.n7194_cascade_ ;
    wire \c0.n8449 ;
    wire n4839;
    wire n4839_cascade_;
    wire n31;
    wire data_in_field_65;
    wire \c0.tx2_transmit_N_1444 ;
    wire bfn_7_25_0_;
    wire \c0.n8113 ;
    wire \c0.n8114 ;
    wire \c0.n8115 ;
    wire \c0.n8116 ;
    wire \c0.byte_transmit_counter2_5 ;
    wire \c0.n8117 ;
    wire \c0.byte_transmit_counter2_6 ;
    wire \c0.n8118 ;
    wire \c0.n8119 ;
    wire \c0.byte_transmit_counter2_7 ;
    wire \c0.n4897 ;
    wire \c0.n5154 ;
    wire rand_data_8;
    wire rand_data_22;
    wire rand_data_3;
    wire \c0.n8992 ;
    wire \c0.n21_adj_1624 ;
    wire rand_data_7;
    wire rand_data_1;
    wire rand_data_15;
    wire data_in_field_143;
    wire rand_data_28;
    wire rand_data_13;
    wire \c0.data_in_field_29 ;
    wire \c0.data_in_field_21 ;
    wire \c0.n9608_cascade_ ;
    wire \c0.data_in_field_5 ;
    wire \c0.n9147 ;
    wire rand_data_29;
    wire data_in_field_109;
    wire rand_data_4;
    wire \c0.n8942 ;
    wire data_in_field_57;
    wire data_in_field_93;
    wire \c0.n4390 ;
    wire data_in_field_87;
    wire data_in_field_91;
    wire \c0.n8909 ;
    wire \c0.n4197 ;
    wire data_in_field_60;
    wire \c0.n4197_cascade_ ;
    wire \c0.n4399 ;
    wire data_in_field_61;
    wire \c0.n4399_cascade_ ;
    wire \c0.n4288 ;
    wire \c0.n10 ;
    wire rand_data_9;
    wire data_in_field_121;
    wire data_in_field_44;
    wire \c0.n9572 ;
    wire data_in_field_77;
    wire data_in_field_49;
    wire \c0.n8887_cascade_ ;
    wire data_in_field_120;
    wire rand_data_30;
    wire \c0.n8785 ;
    wire \c0.n8887 ;
    wire \c0.n4240_cascade_ ;
    wire \c0.data_in_field_13 ;
    wire \c0.n44_adj_1609 ;
    wire \c0.n4553 ;
    wire data_in_field_53;
    wire \c0.n8964 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \c0.n18_adj_1666 ;
    wire data_in_field_36;
    wire \c0.n1645 ;
    wire data_in_field_62;
    wire data_in_field_46;
    wire \c0.n9632_cascade_ ;
    wire \c0.data_in_field_38 ;
    wire data_in_field_126;
    wire \c0.n9620_cascade_ ;
    wire data_in_field_94;
    wire \c0.n9626_cascade_ ;
    wire \c0.n9141 ;
    wire \c0.n9138_cascade_ ;
    wire \c0.n9132 ;
    wire \c0.n9135 ;
    wire \c0.n9614_cascade_ ;
    wire \c0.n9617_cascade_ ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire data_in_11_2;
    wire data_in_12_2;
    wire data_in_13_2;
    wire data_in_14_2;
    wire data_in_15_2;
    wire data_in_16_2;
    wire data_in_18_2;
    wire data_in_17_2;
    wire data_in_20_2;
    wire data_in_19_2;
    wire n7171;
    wire \c0.n9668 ;
    wire \c0.n8878 ;
    wire \c0.n8813 ;
    wire data_in_field_43;
    wire \c0.n28_adj_1619 ;
    wire \c0.n29_adj_1620_cascade_ ;
    wire \c0.data_in_frame_19_6 ;
    wire n1901;
    wire FRAME_MATCHER_state_2;
    wire \c0.n7194 ;
    wire n9262;
    wire data_in_6_2;
    wire FRAME_MATCHER_state_0;
    wire n1893;
    wire data_in_7_2;
    wire data_in_8_2;
    wire data_in_10_2;
    wire data_in_9_2;
    wire \c0.n8921 ;
    wire \c0.n4562_cascade_ ;
    wire \c0.n4479 ;
    wire \c0.n4235_cascade_ ;
    wire \c0.n4562 ;
    wire data_in_field_99;
    wire data_in_field_131;
    wire \c0.n8846 ;
    wire rand_data_2;
    wire \c0.n30 ;
    wire rand_data_26;
    wire data_in_field_58;
    wire data_in_field_118;
    wire \c0.n4534 ;
    wire \c0.n27_adj_1621 ;
    wire rand_data_10;
    wire \c0.n4473 ;
    wire \c0.n4473_cascade_ ;
    wire \c0.n9010 ;
    wire \c0.n4244_cascade_ ;
    wire rand_data_6;
    wire data_in_field_102;
    wire data_in_field_125;
    wire data_in_field_73;
    wire \c0.n18_adj_1618 ;
    wire data_in_field_54;
    wire data_in_field_69;
    wire \c0.n8998 ;
    wire \c0.n16_adj_1591 ;
    wire rand_data_20;
    wire data_in_field_124;
    wire data_in_field_116;
    wire data_in_field_56;
    wire data_in_field_101;
    wire rand_data_16;
    wire \c0.n8788 ;
    wire \c0.n8828 ;
    wire \c0.n8855 ;
    wire \c0.n35 ;
    wire data_in_field_84;
    wire data_in_field_92;
    wire \c0.n9560 ;
    wire data_in_field_108;
    wire data_in_field_100;
    wire \c0.n8927 ;
    wire \c0.n8837 ;
    wire data_in_field_41;
    wire \c0.n16_adj_1629 ;
    wire \c0.n8977 ;
    wire \c0.n17_adj_1630 ;
    wire \c0.data_in_frame_19_4 ;
    wire \c0.data_in_frame_20_4 ;
    wire data_in_field_68;
    wire data_in_field_76;
    wire \c0.n9566 ;
    wire \c0.n9171 ;
    wire \c0.n9168_cascade_ ;
    wire \c0.n9165 ;
    wire \c0.n9162 ;
    wire \c0.n9554 ;
    wire \c0.n22_adj_1679 ;
    wire \c0.n9557_cascade_ ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire n5185_cascade_;
    wire data_in_field_150;
    wire data_in_field_52;
    wire data_in_field_151;
    wire data_in_field_86;
    wire \c0.n8915 ;
    wire n9077;
    wire n5185;
    wire r_Bit_Index_0_adj_1733;
    wire r_Bit_Index_1_adj_1732;
    wire n4_adj_1724;
    wire data_in_field_134;
    wire data_in_field_119;
    wire \c0.n8883 ;
    wire \c0.n8770 ;
    wire \c0.n8810 ;
    wire \c0.n8899 ;
    wire \c0.n16_adj_1657 ;
    wire \c0.n22_adj_1655_cascade_ ;
    wire data_in_field_37;
    wire \c0.n24_adj_1658 ;
    wire \c0.n8939 ;
    wire \c0.n20_adj_1659 ;
    wire \c0.data_in_frame_19_0 ;
    wire data_in_field_136;
    wire \c0.n9536_cascade_ ;
    wire data_in_field_128;
    wire \c0.n9539_cascade_ ;
    wire rand_data_18;
    wire data_in_field_114;
    wire data_in_field_144;
    wire \c0.n8971 ;
    wire \c0.n6_adj_1628 ;
    wire rand_data_0;
    wire \c0.n8918 ;
    wire \c0.n8840_cascade_ ;
    wire \c0.n4511 ;
    wire \c0.n4309 ;
    wire rand_data_11;
    wire data_in_field_123;
    wire data_in_field_146;
    wire data_in_field_130;
    wire \c0.n9698_cascade_ ;
    wire data_in_field_138;
    wire \c0.n9701_cascade_ ;
    wire data_in_field_142;
    wire data_in_field_78;
    wire \c0.n4215 ;
    wire \c0.n8912 ;
    wire \c0.n8954 ;
    wire \c0.n8819_cascade_ ;
    wire \c0.n4365 ;
    wire \c0.n21_adj_1644_cascade_ ;
    wire \c0.n19_adj_1643 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.n8782 ;
    wire \c0.n8807 ;
    wire data_in_field_110;
    wire \c0.n8819 ;
    wire \c0.n8893 ;
    wire \c0.n8427 ;
    wire \c0.n28_adj_1612 ;
    wire \c0.n26_adj_1613 ;
    wire \c0.n27_cascade_ ;
    wire \c0.n25_adj_1614 ;
    wire \c0.data_in_frame_20_0 ;
    wire \c0.n8995 ;
    wire \c0.n8834 ;
    wire \c0.n8924 ;
    wire \c0.n8852 ;
    wire \c0.n9013 ;
    wire data_in_field_70;
    wire \c0.n12_cascade_ ;
    wire data_in_field_112;
    wire \c0.data_in_frame_20_2 ;
    wire data_in_5_2;
    wire data_in_4_2;
    wire r_SM_Main_2_adj_1738;
    wire \c0.tx2.n4880 ;
    wire \c0.n4525 ;
    wire \c0.n4244 ;
    wire data_in_field_50;
    wire \c0.n20_adj_1642 ;
    wire n12_adj_1753_cascade_;
    wire r_SM_Main_2_N_1537_2_cascade_;
    wire \c0.rx.n4090 ;
    wire \c0.rx.n7393 ;
    wire data_in_field_122;
    wire \c0.n4537 ;
    wire \c0.rx.r_SM_Main_2_N_1543_0_cascade_ ;
    wire n6_adj_1751_cascade_;
    wire n30_cascade_;
    wire data_in_field_97;
    wire data_in_field_95;
    wire data_in_field_96;
    wire \c0.n4296 ;
    wire \c0.rx.n12 ;
    wire tx_enable;
    wire n2185;
    wire r_Bit_Index_2_adj_1731;
    wire n7415_cascade_;
    wire n9301_cascade_;
    wire n1;
    wire r_Rx_Data;
    wire \c0.rx.r_SM_Main_2_N_1543_0 ;
    wire n9300;
    wire \c0.data_in_field_24 ;
    wire \c0.data_in_field_16 ;
    wire \c0.data_in_field_8 ;
    wire \c0.data_in_field_0 ;
    wire \c0.n9446_cascade_ ;
    wire \c0.n9228 ;
    wire \c0.n9449_cascade_ ;
    wire data_in_field_80;
    wire data_in_field_72;
    wire \c0.n9740_cascade_ ;
    wire data_in_field_64;
    wire \c0.n9234 ;
    wire \c0.n9231_cascade_ ;
    wire \c0.n9728 ;
    wire \c0.n22_adj_1661 ;
    wire \c0.n9731 ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire rx_data_ready;
    wire data_in_19_0;
    wire data_in_18_0;
    wire rand_data_12;
    wire n4806;
    wire data_in_field_88;
    wire \c0.n4292 ;
    wire \c0.n8957 ;
    wire \c0.data_in_field_27 ;
    wire \c0.data_in_field_25 ;
    wire \c0.n8871 ;
    wire n26;
    wire bfn_11_27_0_;
    wire n25_adj_1722;
    wire n8130;
    wire n24;
    wire n8131;
    wire n23;
    wire n8132;
    wire n22;
    wire n8133;
    wire n21;
    wire n8134;
    wire n20;
    wire n8135;
    wire n19;
    wire n8136;
    wire n8137;
    wire n18;
    wire bfn_11_28_0_;
    wire n17;
    wire n8138;
    wire n16;
    wire n8139;
    wire n15;
    wire n8140;
    wire n14;
    wire n8141;
    wire n13;
    wire n8142;
    wire n12;
    wire n8143;
    wire n11;
    wire n8144;
    wire n8145;
    wire n10;
    wire bfn_11_29_0_;
    wire n9;
    wire n8146;
    wire n8;
    wire n8147;
    wire n7;
    wire n8148;
    wire n6;
    wire n8149;
    wire blink_counter_21;
    wire n8150;
    wire blink_counter_22;
    wire n8151;
    wire blink_counter_23;
    wire n8152;
    wire n8153;
    wire blink_counter_24;
    wire bfn_11_30_0_;
    wire n8154;
    wire blink_counter_25;
    wire r_SM_Main_1_adj_1735;
    wire n9246;
    wire r_SM_Main_0_adj_1736;
    wire n44_cascade_;
    wire r_SM_Main_2_adj_1734;
    wire r_SM_Main_2_N_1537_2;
    wire n9245;
    wire r_Clock_Count_0_adj_1730;
    wire n226;
    wire bfn_11_31_0_;
    wire r_Clock_Count_1;
    wire n225;
    wire \c0.rx.n8098 ;
    wire r_Clock_Count_2;
    wire n224;
    wire \c0.rx.n8099 ;
    wire r_Clock_Count_3;
    wire n223;
    wire \c0.rx.n8100 ;
    wire \c0.rx.n8101 ;
    wire \c0.rx.n8102 ;
    wire r_Clock_Count_6_adj_1728;
    wire n220;
    wire \c0.rx.n8103 ;
    wire r_Clock_Count_7_adj_1727;
    wire \c0.rx.n8104 ;
    wire n219;
    wire n4084;
    wire n221;
    wire r_Clock_Count_5;
    wire n30;
    wire n222;
    wire n44;
    wire r_Clock_Count_4_adj_1729;
    wire \c0.n9192 ;
    wire \c0.n9195 ;
    wire \c0.n22_adj_1681 ;
    wire \c0.n9491_cascade_ ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.tx2.n3760 ;
    wire data_in_field_82;
    wire data_in_field_90;
    wire \c0.byte_transmit_counter2_0 ;
    wire data_in_field_66;
    wire data_in_field_74;
    wire \c0.n9500 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.n9198_cascade_ ;
    wire \c0.n9488 ;
    wire data_in_field_98;
    wire \c0.n9494 ;
    wire data_in_field_106;
    wire \c0.n9201 ;
    wire \c0.n3056 ;
    wire \c0.n9671 ;
    wire \c0.data_in_frame_20_6 ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n22_adj_1677 ;
    wire bfn_13_26_0_;
    wire \c0.n8083 ;
    wire \c0.n8084 ;
    wire \c0.n8085 ;
    wire \c0.n8086 ;
    wire \c0.n8087 ;
    wire \c0.n8088 ;
    wire \c0.n8089 ;
    wire \c0.n11_cascade_ ;
    wire tx_data_3_N_keep_cascade_;
    wire tx_data_0_N_keep;
    wire data_in_field_133;
    wire data_in_field_103;
    wire data_in_field_148;
    wire \c0.n8986 ;
    wire \c0.n45_adj_1656 ;
    wire tx_data_5_N_keep_cascade_;
    wire \c0.n11 ;
    wire tx_data_2_N_keep_cascade_;
    wire tx_data_6_N_keep;
    wire n8705_cascade_;
    wire r_Tx_Data_6;
    wire r_Tx_Data_2;
    wire data_in_field_132;
    wire \c0.n9680 ;
    wire data_in_field_140;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.n9683 ;
    wire \c0.n17_adj_1663_cascade_ ;
    wire \c0.n123_cascade_ ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.data_out_6_7_N_965_3 ;
    wire \c0.data_out_6_7_N_965_2 ;
    wire \c0.data_out_6_7_N_965_0 ;
    wire \c0.data_out_6_7_N_965_6 ;
    wire \c0.data_out_6_7_N_965_4 ;
    wire \c0.data_out_6_7_N_965_7 ;
    wire \c0.n7_cascade_ ;
    wire \c0.n8 ;
    wire \c0.n7814_cascade_ ;
    wire data_out_6_7_N_965_5;
    wire n7204_cascade_;
    wire byte_transmit_counter_5;
    wire \c0.data_out_6_7_N_965_1 ;
    wire n7204;
    wire tx_data_1_N_keep_cascade_;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n7779_cascade_ ;
    wire tx_data_1_N_keep;
    wire \c0.data_out_6__7__N_973 ;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.byte_transmit_counter_4 ;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.byte_transmit_counter_3 ;
    wire \c0.n9291 ;
    wire r_Tx_Data_3;
    wire tx_data_7_N_keep;
    wire r_Tx_Data_7;
    wire r_Tx_Data_1;
    wire r_Tx_Data_5;
    wire n9710;
    wire n9713_cascade_;
    wire n5_cascade_;
    wire n3_cascade_;
    wire tx_o_adj_1726;
    wire n9452;
    wire r_Tx_Data_0;
    wire n9455;
    wire tx_data_4_N_keep;
    wire r_Tx_Data_4;
    wire n9073;
    wire r_Bit_Index_0;
    wire n5062;
    wire n9073_cascade_;
    wire r_Bit_Index_1;
    wire n3892;
    wire \c0.n18_adj_1662 ;
    wire \c0.n19_adj_1664 ;
    wire \c0.n123 ;
    wire \c0.n7814 ;
    wire \c0.n117 ;
    wire n3747;
    wire \c0.tx_active_prev ;
    wire n8749_cascade_;
    wire tx_active;
    wire \c0.tx.n8_cascade_ ;
    wire \c0.tx.n9059 ;
    wire n28;
    wire \c0.tx_transmit ;
    wire n3151_cascade_;
    wire n11_adj_1752;
    wire \c0.tx.n5_cascade_ ;
    wire r_SM_Main_0;
    wire \c0.tx.n23_cascade_ ;
    wire r_SM_Main_1;
    wire n9259;
    wire \c0.tx.n9027 ;
    wire bfn_15_30_0_;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.tx.n9290 ;
    wire \c0.tx.n8090 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n9313 ;
    wire \c0.tx.n8091 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.n9281 ;
    wire \c0.tx.n8092 ;
    wire \c0.tx.n8093 ;
    wire \c0.tx.n8094 ;
    wire r_Clock_Count_6;
    wire n9304;
    wire \c0.tx.n8095 ;
    wire \c0.tx.n8096 ;
    wire \c0.tx.n8097 ;
    wire \c0.tx.n7916 ;
    wire bfn_15_31_0_;
    wire n9249;
    wire r_Clock_Count_0;
    wire n9266;
    wire \c0.n900 ;
    wire \c0.n22 ;
    wire \c0.delay_counter_0 ;
    wire bfn_16_25_0_;
    wire \c0.n21_adj_1653 ;
    wire \c0.delay_counter_1 ;
    wire \c0.n8120 ;
    wire \c0.n20_adj_1652 ;
    wire \c0.delay_counter_2 ;
    wire \c0.n8121 ;
    wire \c0.n19_adj_1651 ;
    wire \c0.delay_counter_3 ;
    wire \c0.n8122 ;
    wire \c0.n18_adj_1650 ;
    wire \c0.delay_counter_4 ;
    wire \c0.n8123 ;
    wire \c0.n17_adj_1649 ;
    wire \c0.delay_counter_5 ;
    wire \c0.n8124 ;
    wire \c0.n16_adj_1641 ;
    wire \c0.delay_counter_6 ;
    wire \c0.n8125 ;
    wire \c0.n15 ;
    wire \c0.delay_counter_7 ;
    wire \c0.n8126 ;
    wire \c0.n8127 ;
    wire \c0.n14_adj_1639 ;
    wire \c0.delay_counter_8 ;
    wire bfn_16_26_0_;
    wire \c0.n13 ;
    wire \c0.delay_counter_9 ;
    wire \c0.n8128 ;
    wire \c0.n12_adj_1634 ;
    wire \c0.n8129 ;
    wire \c0.delay_counter_10 ;
    wire UART_TRANSMITTER_state_0;
    wire r_SM_Main_2_N_1480_1;
    wire \c0.tx.n23 ;
    wire r_Clock_Count_8;
    wire r_Bit_Index_2;
    wire \c0.tx.n9310 ;
    wire n9305;
    wire r_Clock_Count_4;
    wire \c0.tx.n9314 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire r_SM_Main_2;
    wire n9303;
    wire r_Clock_Count_7;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__35917),
            .DIN(N__35916),
            .DOUT(N__35915),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__35917),
            .PADOUT(N__35916),
            .PADIN(N__35915),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19242),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__35908),
            .DIN(N__35907),
            .DOUT(N__35906),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__35908),
            .PADOUT(N__35907),
            .PADIN(N__35906),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__35899),
            .DIN(N__35898),
            .DOUT(N__35897),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__35899),
            .PADOUT(N__35898),
            .PADIN(N__35897),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__35382),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__35890),
            .DIN(N__35889),
            .DOUT(N__35888),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__35890),
            .PADOUT(N__35889),
            .PADIN(N__35888),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15786),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13179));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__35881),
            .DIN(N__35880),
            .DOUT(N__35879),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__35881),
            .PADOUT(N__35880),
            .PADIN(N__35879),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34119),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__27585));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__35872),
            .DIN(N__35871),
            .DOUT(N__35870),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__35872),
            .PADOUT(N__35871),
            .PADIN(N__35870),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__8861 (
            .O(N__35853),
            .I(\c0.n8129 ));
    InMux I__8860 (
            .O(N__35850),
            .I(N__35847));
    LocalMux I__8859 (
            .O(N__35847),
            .I(N__35843));
    InMux I__8858 (
            .O(N__35846),
            .I(N__35840));
    Span4Mux_h I__8857 (
            .O(N__35843),
            .I(N__35837));
    LocalMux I__8856 (
            .O(N__35840),
            .I(\c0.delay_counter_10 ));
    Odrv4 I__8855 (
            .O(N__35837),
            .I(\c0.delay_counter_10 ));
    CEMux I__8854 (
            .O(N__35832),
            .I(N__35828));
    CEMux I__8853 (
            .O(N__35831),
            .I(N__35824));
    LocalMux I__8852 (
            .O(N__35828),
            .I(N__35821));
    CascadeMux I__8851 (
            .O(N__35827),
            .I(N__35818));
    LocalMux I__8850 (
            .O(N__35824),
            .I(N__35809));
    Span4Mux_h I__8849 (
            .O(N__35821),
            .I(N__35806));
    InMux I__8848 (
            .O(N__35818),
            .I(N__35799));
    InMux I__8847 (
            .O(N__35817),
            .I(N__35799));
    InMux I__8846 (
            .O(N__35816),
            .I(N__35799));
    CascadeMux I__8845 (
            .O(N__35815),
            .I(N__35796));
    CascadeMux I__8844 (
            .O(N__35814),
            .I(N__35793));
    CascadeMux I__8843 (
            .O(N__35813),
            .I(N__35790));
    CascadeMux I__8842 (
            .O(N__35812),
            .I(N__35787));
    Span4Mux_h I__8841 (
            .O(N__35809),
            .I(N__35781));
    Sp12to4 I__8840 (
            .O(N__35806),
            .I(N__35778));
    LocalMux I__8839 (
            .O(N__35799),
            .I(N__35775));
    InMux I__8838 (
            .O(N__35796),
            .I(N__35772));
    InMux I__8837 (
            .O(N__35793),
            .I(N__35769));
    InMux I__8836 (
            .O(N__35790),
            .I(N__35758));
    InMux I__8835 (
            .O(N__35787),
            .I(N__35758));
    InMux I__8834 (
            .O(N__35786),
            .I(N__35758));
    InMux I__8833 (
            .O(N__35785),
            .I(N__35758));
    InMux I__8832 (
            .O(N__35784),
            .I(N__35758));
    Odrv4 I__8831 (
            .O(N__35781),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__8830 (
            .O(N__35778),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__8829 (
            .O(N__35775),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__8828 (
            .O(N__35772),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__8827 (
            .O(N__35769),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__8826 (
            .O(N__35758),
            .I(UART_TRANSMITTER_state_0));
    InMux I__8825 (
            .O(N__35745),
            .I(N__35741));
    CascadeMux I__8824 (
            .O(N__35744),
            .I(N__35738));
    LocalMux I__8823 (
            .O(N__35741),
            .I(N__35732));
    InMux I__8822 (
            .O(N__35738),
            .I(N__35725));
    InMux I__8821 (
            .O(N__35737),
            .I(N__35725));
    InMux I__8820 (
            .O(N__35736),
            .I(N__35725));
    InMux I__8819 (
            .O(N__35735),
            .I(N__35722));
    Span4Mux_v I__8818 (
            .O(N__35732),
            .I(N__35719));
    LocalMux I__8817 (
            .O(N__35725),
            .I(r_SM_Main_2_N_1480_1));
    LocalMux I__8816 (
            .O(N__35722),
            .I(r_SM_Main_2_N_1480_1));
    Odrv4 I__8815 (
            .O(N__35719),
            .I(r_SM_Main_2_N_1480_1));
    InMux I__8814 (
            .O(N__35712),
            .I(N__35704));
    InMux I__8813 (
            .O(N__35711),
            .I(N__35704));
    InMux I__8812 (
            .O(N__35710),
            .I(N__35699));
    InMux I__8811 (
            .O(N__35709),
            .I(N__35699));
    LocalMux I__8810 (
            .O(N__35704),
            .I(\c0.tx.n23 ));
    LocalMux I__8809 (
            .O(N__35699),
            .I(\c0.tx.n23 ));
    CascadeMux I__8808 (
            .O(N__35694),
            .I(N__35691));
    InMux I__8807 (
            .O(N__35691),
            .I(N__35684));
    InMux I__8806 (
            .O(N__35690),
            .I(N__35684));
    InMux I__8805 (
            .O(N__35689),
            .I(N__35678));
    LocalMux I__8804 (
            .O(N__35684),
            .I(N__35675));
    InMux I__8803 (
            .O(N__35683),
            .I(N__35672));
    InMux I__8802 (
            .O(N__35682),
            .I(N__35669));
    InMux I__8801 (
            .O(N__35681),
            .I(N__35666));
    LocalMux I__8800 (
            .O(N__35678),
            .I(N__35661));
    Span4Mux_h I__8799 (
            .O(N__35675),
            .I(N__35661));
    LocalMux I__8798 (
            .O(N__35672),
            .I(N__35658));
    LocalMux I__8797 (
            .O(N__35669),
            .I(r_Clock_Count_8));
    LocalMux I__8796 (
            .O(N__35666),
            .I(r_Clock_Count_8));
    Odrv4 I__8795 (
            .O(N__35661),
            .I(r_Clock_Count_8));
    Odrv12 I__8794 (
            .O(N__35658),
            .I(r_Clock_Count_8));
    InMux I__8793 (
            .O(N__35649),
            .I(N__35646));
    LocalMux I__8792 (
            .O(N__35646),
            .I(N__35642));
    InMux I__8791 (
            .O(N__35645),
            .I(N__35639));
    Span4Mux_v I__8790 (
            .O(N__35642),
            .I(N__35633));
    LocalMux I__8789 (
            .O(N__35639),
            .I(N__35633));
    InMux I__8788 (
            .O(N__35638),
            .I(N__35627));
    Span4Mux_h I__8787 (
            .O(N__35633),
            .I(N__35624));
    InMux I__8786 (
            .O(N__35632),
            .I(N__35617));
    InMux I__8785 (
            .O(N__35631),
            .I(N__35617));
    InMux I__8784 (
            .O(N__35630),
            .I(N__35617));
    LocalMux I__8783 (
            .O(N__35627),
            .I(r_Bit_Index_2));
    Odrv4 I__8782 (
            .O(N__35624),
            .I(r_Bit_Index_2));
    LocalMux I__8781 (
            .O(N__35617),
            .I(r_Bit_Index_2));
    InMux I__8780 (
            .O(N__35610),
            .I(N__35607));
    LocalMux I__8779 (
            .O(N__35607),
            .I(\c0.tx.n9310 ));
    InMux I__8778 (
            .O(N__35604),
            .I(N__35601));
    LocalMux I__8777 (
            .O(N__35601),
            .I(n9305));
    InMux I__8776 (
            .O(N__35598),
            .I(N__35593));
    InMux I__8775 (
            .O(N__35597),
            .I(N__35590));
    InMux I__8774 (
            .O(N__35596),
            .I(N__35587));
    LocalMux I__8773 (
            .O(N__35593),
            .I(r_Clock_Count_4));
    LocalMux I__8772 (
            .O(N__35590),
            .I(r_Clock_Count_4));
    LocalMux I__8771 (
            .O(N__35587),
            .I(r_Clock_Count_4));
    InMux I__8770 (
            .O(N__35580),
            .I(N__35577));
    LocalMux I__8769 (
            .O(N__35577),
            .I(\c0.tx.n9314 ));
    InMux I__8768 (
            .O(N__35574),
            .I(N__35569));
    InMux I__8767 (
            .O(N__35573),
            .I(N__35566));
    InMux I__8766 (
            .O(N__35572),
            .I(N__35563));
    LocalMux I__8765 (
            .O(N__35569),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__8764 (
            .O(N__35566),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__8763 (
            .O(N__35563),
            .I(\c0.tx.r_Clock_Count_5 ));
    CascadeMux I__8762 (
            .O(N__35556),
            .I(N__35547));
    InMux I__8761 (
            .O(N__35555),
            .I(N__35540));
    InMux I__8760 (
            .O(N__35554),
            .I(N__35540));
    InMux I__8759 (
            .O(N__35553),
            .I(N__35531));
    InMux I__8758 (
            .O(N__35552),
            .I(N__35526));
    InMux I__8757 (
            .O(N__35551),
            .I(N__35526));
    InMux I__8756 (
            .O(N__35550),
            .I(N__35517));
    InMux I__8755 (
            .O(N__35547),
            .I(N__35517));
    InMux I__8754 (
            .O(N__35546),
            .I(N__35517));
    InMux I__8753 (
            .O(N__35545),
            .I(N__35517));
    LocalMux I__8752 (
            .O(N__35540),
            .I(N__35509));
    InMux I__8751 (
            .O(N__35539),
            .I(N__35506));
    InMux I__8750 (
            .O(N__35538),
            .I(N__35503));
    InMux I__8749 (
            .O(N__35537),
            .I(N__35498));
    InMux I__8748 (
            .O(N__35536),
            .I(N__35498));
    InMux I__8747 (
            .O(N__35535),
            .I(N__35493));
    InMux I__8746 (
            .O(N__35534),
            .I(N__35493));
    LocalMux I__8745 (
            .O(N__35531),
            .I(N__35486));
    LocalMux I__8744 (
            .O(N__35526),
            .I(N__35486));
    LocalMux I__8743 (
            .O(N__35517),
            .I(N__35486));
    InMux I__8742 (
            .O(N__35516),
            .I(N__35475));
    InMux I__8741 (
            .O(N__35515),
            .I(N__35475));
    InMux I__8740 (
            .O(N__35514),
            .I(N__35475));
    InMux I__8739 (
            .O(N__35513),
            .I(N__35475));
    InMux I__8738 (
            .O(N__35512),
            .I(N__35475));
    Odrv4 I__8737 (
            .O(N__35509),
            .I(r_SM_Main_2));
    LocalMux I__8736 (
            .O(N__35506),
            .I(r_SM_Main_2));
    LocalMux I__8735 (
            .O(N__35503),
            .I(r_SM_Main_2));
    LocalMux I__8734 (
            .O(N__35498),
            .I(r_SM_Main_2));
    LocalMux I__8733 (
            .O(N__35493),
            .I(r_SM_Main_2));
    Odrv4 I__8732 (
            .O(N__35486),
            .I(r_SM_Main_2));
    LocalMux I__8731 (
            .O(N__35475),
            .I(r_SM_Main_2));
    InMux I__8730 (
            .O(N__35460),
            .I(N__35457));
    LocalMux I__8729 (
            .O(N__35457),
            .I(n9303));
    InMux I__8728 (
            .O(N__35454),
            .I(N__35449));
    InMux I__8727 (
            .O(N__35453),
            .I(N__35446));
    InMux I__8726 (
            .O(N__35452),
            .I(N__35443));
    LocalMux I__8725 (
            .O(N__35449),
            .I(r_Clock_Count_7));
    LocalMux I__8724 (
            .O(N__35446),
            .I(r_Clock_Count_7));
    LocalMux I__8723 (
            .O(N__35443),
            .I(r_Clock_Count_7));
    ClkMux I__8722 (
            .O(N__35436),
            .I(N__34995));
    ClkMux I__8721 (
            .O(N__35435),
            .I(N__34995));
    ClkMux I__8720 (
            .O(N__35434),
            .I(N__34995));
    ClkMux I__8719 (
            .O(N__35433),
            .I(N__34995));
    ClkMux I__8718 (
            .O(N__35432),
            .I(N__34995));
    ClkMux I__8717 (
            .O(N__35431),
            .I(N__34995));
    ClkMux I__8716 (
            .O(N__35430),
            .I(N__34995));
    ClkMux I__8715 (
            .O(N__35429),
            .I(N__34995));
    ClkMux I__8714 (
            .O(N__35428),
            .I(N__34995));
    ClkMux I__8713 (
            .O(N__35427),
            .I(N__34995));
    ClkMux I__8712 (
            .O(N__35426),
            .I(N__34995));
    ClkMux I__8711 (
            .O(N__35425),
            .I(N__34995));
    ClkMux I__8710 (
            .O(N__35424),
            .I(N__34995));
    ClkMux I__8709 (
            .O(N__35423),
            .I(N__34995));
    ClkMux I__8708 (
            .O(N__35422),
            .I(N__34995));
    ClkMux I__8707 (
            .O(N__35421),
            .I(N__34995));
    ClkMux I__8706 (
            .O(N__35420),
            .I(N__34995));
    ClkMux I__8705 (
            .O(N__35419),
            .I(N__34995));
    ClkMux I__8704 (
            .O(N__35418),
            .I(N__34995));
    ClkMux I__8703 (
            .O(N__35417),
            .I(N__34995));
    ClkMux I__8702 (
            .O(N__35416),
            .I(N__34995));
    ClkMux I__8701 (
            .O(N__35415),
            .I(N__34995));
    ClkMux I__8700 (
            .O(N__35414),
            .I(N__34995));
    ClkMux I__8699 (
            .O(N__35413),
            .I(N__34995));
    ClkMux I__8698 (
            .O(N__35412),
            .I(N__34995));
    ClkMux I__8697 (
            .O(N__35411),
            .I(N__34995));
    ClkMux I__8696 (
            .O(N__35410),
            .I(N__34995));
    ClkMux I__8695 (
            .O(N__35409),
            .I(N__34995));
    ClkMux I__8694 (
            .O(N__35408),
            .I(N__34995));
    ClkMux I__8693 (
            .O(N__35407),
            .I(N__34995));
    ClkMux I__8692 (
            .O(N__35406),
            .I(N__34995));
    ClkMux I__8691 (
            .O(N__35405),
            .I(N__34995));
    ClkMux I__8690 (
            .O(N__35404),
            .I(N__34995));
    ClkMux I__8689 (
            .O(N__35403),
            .I(N__34995));
    ClkMux I__8688 (
            .O(N__35402),
            .I(N__34995));
    ClkMux I__8687 (
            .O(N__35401),
            .I(N__34995));
    ClkMux I__8686 (
            .O(N__35400),
            .I(N__34995));
    ClkMux I__8685 (
            .O(N__35399),
            .I(N__34995));
    ClkMux I__8684 (
            .O(N__35398),
            .I(N__34995));
    ClkMux I__8683 (
            .O(N__35397),
            .I(N__34995));
    ClkMux I__8682 (
            .O(N__35396),
            .I(N__34995));
    ClkMux I__8681 (
            .O(N__35395),
            .I(N__34995));
    ClkMux I__8680 (
            .O(N__35394),
            .I(N__34995));
    ClkMux I__8679 (
            .O(N__35393),
            .I(N__34995));
    ClkMux I__8678 (
            .O(N__35392),
            .I(N__34995));
    ClkMux I__8677 (
            .O(N__35391),
            .I(N__34995));
    ClkMux I__8676 (
            .O(N__35390),
            .I(N__34995));
    ClkMux I__8675 (
            .O(N__35389),
            .I(N__34995));
    ClkMux I__8674 (
            .O(N__35388),
            .I(N__34995));
    ClkMux I__8673 (
            .O(N__35387),
            .I(N__34995));
    ClkMux I__8672 (
            .O(N__35386),
            .I(N__34995));
    ClkMux I__8671 (
            .O(N__35385),
            .I(N__34995));
    ClkMux I__8670 (
            .O(N__35384),
            .I(N__34995));
    ClkMux I__8669 (
            .O(N__35383),
            .I(N__34995));
    ClkMux I__8668 (
            .O(N__35382),
            .I(N__34995));
    ClkMux I__8667 (
            .O(N__35381),
            .I(N__34995));
    ClkMux I__8666 (
            .O(N__35380),
            .I(N__34995));
    ClkMux I__8665 (
            .O(N__35379),
            .I(N__34995));
    ClkMux I__8664 (
            .O(N__35378),
            .I(N__34995));
    ClkMux I__8663 (
            .O(N__35377),
            .I(N__34995));
    ClkMux I__8662 (
            .O(N__35376),
            .I(N__34995));
    ClkMux I__8661 (
            .O(N__35375),
            .I(N__34995));
    ClkMux I__8660 (
            .O(N__35374),
            .I(N__34995));
    ClkMux I__8659 (
            .O(N__35373),
            .I(N__34995));
    ClkMux I__8658 (
            .O(N__35372),
            .I(N__34995));
    ClkMux I__8657 (
            .O(N__35371),
            .I(N__34995));
    ClkMux I__8656 (
            .O(N__35370),
            .I(N__34995));
    ClkMux I__8655 (
            .O(N__35369),
            .I(N__34995));
    ClkMux I__8654 (
            .O(N__35368),
            .I(N__34995));
    ClkMux I__8653 (
            .O(N__35367),
            .I(N__34995));
    ClkMux I__8652 (
            .O(N__35366),
            .I(N__34995));
    ClkMux I__8651 (
            .O(N__35365),
            .I(N__34995));
    ClkMux I__8650 (
            .O(N__35364),
            .I(N__34995));
    ClkMux I__8649 (
            .O(N__35363),
            .I(N__34995));
    ClkMux I__8648 (
            .O(N__35362),
            .I(N__34995));
    ClkMux I__8647 (
            .O(N__35361),
            .I(N__34995));
    ClkMux I__8646 (
            .O(N__35360),
            .I(N__34995));
    ClkMux I__8645 (
            .O(N__35359),
            .I(N__34995));
    ClkMux I__8644 (
            .O(N__35358),
            .I(N__34995));
    ClkMux I__8643 (
            .O(N__35357),
            .I(N__34995));
    ClkMux I__8642 (
            .O(N__35356),
            .I(N__34995));
    ClkMux I__8641 (
            .O(N__35355),
            .I(N__34995));
    ClkMux I__8640 (
            .O(N__35354),
            .I(N__34995));
    ClkMux I__8639 (
            .O(N__35353),
            .I(N__34995));
    ClkMux I__8638 (
            .O(N__35352),
            .I(N__34995));
    ClkMux I__8637 (
            .O(N__35351),
            .I(N__34995));
    ClkMux I__8636 (
            .O(N__35350),
            .I(N__34995));
    ClkMux I__8635 (
            .O(N__35349),
            .I(N__34995));
    ClkMux I__8634 (
            .O(N__35348),
            .I(N__34995));
    ClkMux I__8633 (
            .O(N__35347),
            .I(N__34995));
    ClkMux I__8632 (
            .O(N__35346),
            .I(N__34995));
    ClkMux I__8631 (
            .O(N__35345),
            .I(N__34995));
    ClkMux I__8630 (
            .O(N__35344),
            .I(N__34995));
    ClkMux I__8629 (
            .O(N__35343),
            .I(N__34995));
    ClkMux I__8628 (
            .O(N__35342),
            .I(N__34995));
    ClkMux I__8627 (
            .O(N__35341),
            .I(N__34995));
    ClkMux I__8626 (
            .O(N__35340),
            .I(N__34995));
    ClkMux I__8625 (
            .O(N__35339),
            .I(N__34995));
    ClkMux I__8624 (
            .O(N__35338),
            .I(N__34995));
    ClkMux I__8623 (
            .O(N__35337),
            .I(N__34995));
    ClkMux I__8622 (
            .O(N__35336),
            .I(N__34995));
    ClkMux I__8621 (
            .O(N__35335),
            .I(N__34995));
    ClkMux I__8620 (
            .O(N__35334),
            .I(N__34995));
    ClkMux I__8619 (
            .O(N__35333),
            .I(N__34995));
    ClkMux I__8618 (
            .O(N__35332),
            .I(N__34995));
    ClkMux I__8617 (
            .O(N__35331),
            .I(N__34995));
    ClkMux I__8616 (
            .O(N__35330),
            .I(N__34995));
    ClkMux I__8615 (
            .O(N__35329),
            .I(N__34995));
    ClkMux I__8614 (
            .O(N__35328),
            .I(N__34995));
    ClkMux I__8613 (
            .O(N__35327),
            .I(N__34995));
    ClkMux I__8612 (
            .O(N__35326),
            .I(N__34995));
    ClkMux I__8611 (
            .O(N__35325),
            .I(N__34995));
    ClkMux I__8610 (
            .O(N__35324),
            .I(N__34995));
    ClkMux I__8609 (
            .O(N__35323),
            .I(N__34995));
    ClkMux I__8608 (
            .O(N__35322),
            .I(N__34995));
    ClkMux I__8607 (
            .O(N__35321),
            .I(N__34995));
    ClkMux I__8606 (
            .O(N__35320),
            .I(N__34995));
    ClkMux I__8605 (
            .O(N__35319),
            .I(N__34995));
    ClkMux I__8604 (
            .O(N__35318),
            .I(N__34995));
    ClkMux I__8603 (
            .O(N__35317),
            .I(N__34995));
    ClkMux I__8602 (
            .O(N__35316),
            .I(N__34995));
    ClkMux I__8601 (
            .O(N__35315),
            .I(N__34995));
    ClkMux I__8600 (
            .O(N__35314),
            .I(N__34995));
    ClkMux I__8599 (
            .O(N__35313),
            .I(N__34995));
    ClkMux I__8598 (
            .O(N__35312),
            .I(N__34995));
    ClkMux I__8597 (
            .O(N__35311),
            .I(N__34995));
    ClkMux I__8596 (
            .O(N__35310),
            .I(N__34995));
    ClkMux I__8595 (
            .O(N__35309),
            .I(N__34995));
    ClkMux I__8594 (
            .O(N__35308),
            .I(N__34995));
    ClkMux I__8593 (
            .O(N__35307),
            .I(N__34995));
    ClkMux I__8592 (
            .O(N__35306),
            .I(N__34995));
    ClkMux I__8591 (
            .O(N__35305),
            .I(N__34995));
    ClkMux I__8590 (
            .O(N__35304),
            .I(N__34995));
    ClkMux I__8589 (
            .O(N__35303),
            .I(N__34995));
    ClkMux I__8588 (
            .O(N__35302),
            .I(N__34995));
    ClkMux I__8587 (
            .O(N__35301),
            .I(N__34995));
    ClkMux I__8586 (
            .O(N__35300),
            .I(N__34995));
    ClkMux I__8585 (
            .O(N__35299),
            .I(N__34995));
    ClkMux I__8584 (
            .O(N__35298),
            .I(N__34995));
    ClkMux I__8583 (
            .O(N__35297),
            .I(N__34995));
    ClkMux I__8582 (
            .O(N__35296),
            .I(N__34995));
    ClkMux I__8581 (
            .O(N__35295),
            .I(N__34995));
    ClkMux I__8580 (
            .O(N__35294),
            .I(N__34995));
    ClkMux I__8579 (
            .O(N__35293),
            .I(N__34995));
    ClkMux I__8578 (
            .O(N__35292),
            .I(N__34995));
    ClkMux I__8577 (
            .O(N__35291),
            .I(N__34995));
    ClkMux I__8576 (
            .O(N__35290),
            .I(N__34995));
    GlobalMux I__8575 (
            .O(N__34995),
            .I(N__34992));
    gio2CtrlBuf I__8574 (
            .O(N__34992),
            .I(CLK_c));
    InMux I__8573 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__8572 (
            .O(N__34986),
            .I(\c0.n19_adj_1651 ));
    InMux I__8571 (
            .O(N__34983),
            .I(N__34979));
    InMux I__8570 (
            .O(N__34982),
            .I(N__34976));
    LocalMux I__8569 (
            .O(N__34979),
            .I(N__34973));
    LocalMux I__8568 (
            .O(N__34976),
            .I(\c0.delay_counter_3 ));
    Odrv12 I__8567 (
            .O(N__34973),
            .I(\c0.delay_counter_3 ));
    InMux I__8566 (
            .O(N__34968),
            .I(\c0.n8122 ));
    InMux I__8565 (
            .O(N__34965),
            .I(N__34962));
    LocalMux I__8564 (
            .O(N__34962),
            .I(\c0.n18_adj_1650 ));
    CascadeMux I__8563 (
            .O(N__34959),
            .I(N__34955));
    InMux I__8562 (
            .O(N__34958),
            .I(N__34950));
    InMux I__8561 (
            .O(N__34955),
            .I(N__34950));
    LocalMux I__8560 (
            .O(N__34950),
            .I(\c0.delay_counter_4 ));
    InMux I__8559 (
            .O(N__34947),
            .I(\c0.n8123 ));
    InMux I__8558 (
            .O(N__34944),
            .I(N__34941));
    LocalMux I__8557 (
            .O(N__34941),
            .I(\c0.n17_adj_1649 ));
    InMux I__8556 (
            .O(N__34938),
            .I(N__34934));
    InMux I__8555 (
            .O(N__34937),
            .I(N__34931));
    LocalMux I__8554 (
            .O(N__34934),
            .I(\c0.delay_counter_5 ));
    LocalMux I__8553 (
            .O(N__34931),
            .I(\c0.delay_counter_5 ));
    InMux I__8552 (
            .O(N__34926),
            .I(\c0.n8124 ));
    InMux I__8551 (
            .O(N__34923),
            .I(N__34920));
    LocalMux I__8550 (
            .O(N__34920),
            .I(\c0.n16_adj_1641 ));
    InMux I__8549 (
            .O(N__34917),
            .I(N__34913));
    InMux I__8548 (
            .O(N__34916),
            .I(N__34910));
    LocalMux I__8547 (
            .O(N__34913),
            .I(N__34907));
    LocalMux I__8546 (
            .O(N__34910),
            .I(\c0.delay_counter_6 ));
    Odrv12 I__8545 (
            .O(N__34907),
            .I(\c0.delay_counter_6 ));
    InMux I__8544 (
            .O(N__34902),
            .I(\c0.n8125 ));
    InMux I__8543 (
            .O(N__34899),
            .I(N__34896));
    LocalMux I__8542 (
            .O(N__34896),
            .I(\c0.n15 ));
    InMux I__8541 (
            .O(N__34893),
            .I(N__34887));
    InMux I__8540 (
            .O(N__34892),
            .I(N__34887));
    LocalMux I__8539 (
            .O(N__34887),
            .I(\c0.delay_counter_7 ));
    InMux I__8538 (
            .O(N__34884),
            .I(\c0.n8126 ));
    InMux I__8537 (
            .O(N__34881),
            .I(N__34878));
    LocalMux I__8536 (
            .O(N__34878),
            .I(\c0.n14_adj_1639 ));
    InMux I__8535 (
            .O(N__34875),
            .I(N__34871));
    InMux I__8534 (
            .O(N__34874),
            .I(N__34868));
    LocalMux I__8533 (
            .O(N__34871),
            .I(\c0.delay_counter_8 ));
    LocalMux I__8532 (
            .O(N__34868),
            .I(\c0.delay_counter_8 ));
    InMux I__8531 (
            .O(N__34863),
            .I(bfn_16_26_0_));
    InMux I__8530 (
            .O(N__34860),
            .I(N__34857));
    LocalMux I__8529 (
            .O(N__34857),
            .I(\c0.n13 ));
    CascadeMux I__8528 (
            .O(N__34854),
            .I(N__34850));
    InMux I__8527 (
            .O(N__34853),
            .I(N__34847));
    InMux I__8526 (
            .O(N__34850),
            .I(N__34844));
    LocalMux I__8525 (
            .O(N__34847),
            .I(\c0.delay_counter_9 ));
    LocalMux I__8524 (
            .O(N__34844),
            .I(\c0.delay_counter_9 ));
    InMux I__8523 (
            .O(N__34839),
            .I(\c0.n8128 ));
    InMux I__8522 (
            .O(N__34836),
            .I(N__34833));
    LocalMux I__8521 (
            .O(N__34833),
            .I(\c0.n12_adj_1634 ));
    InMux I__8520 (
            .O(N__34830),
            .I(\c0.tx.n8094 ));
    InMux I__8519 (
            .O(N__34827),
            .I(N__34822));
    InMux I__8518 (
            .O(N__34826),
            .I(N__34817));
    InMux I__8517 (
            .O(N__34825),
            .I(N__34817));
    LocalMux I__8516 (
            .O(N__34822),
            .I(r_Clock_Count_6));
    LocalMux I__8515 (
            .O(N__34817),
            .I(r_Clock_Count_6));
    InMux I__8514 (
            .O(N__34812),
            .I(N__34809));
    LocalMux I__8513 (
            .O(N__34809),
            .I(n9304));
    InMux I__8512 (
            .O(N__34806),
            .I(\c0.tx.n8095 ));
    InMux I__8511 (
            .O(N__34803),
            .I(\c0.tx.n8096 ));
    InMux I__8510 (
            .O(N__34800),
            .I(N__34789));
    InMux I__8509 (
            .O(N__34799),
            .I(N__34780));
    InMux I__8508 (
            .O(N__34798),
            .I(N__34780));
    InMux I__8507 (
            .O(N__34797),
            .I(N__34780));
    InMux I__8506 (
            .O(N__34796),
            .I(N__34780));
    InMux I__8505 (
            .O(N__34795),
            .I(N__34771));
    InMux I__8504 (
            .O(N__34794),
            .I(N__34771));
    InMux I__8503 (
            .O(N__34793),
            .I(N__34771));
    InMux I__8502 (
            .O(N__34792),
            .I(N__34771));
    LocalMux I__8501 (
            .O(N__34789),
            .I(N__34768));
    LocalMux I__8500 (
            .O(N__34780),
            .I(\c0.tx.n7916 ));
    LocalMux I__8499 (
            .O(N__34771),
            .I(\c0.tx.n7916 ));
    Odrv4 I__8498 (
            .O(N__34768),
            .I(\c0.tx.n7916 ));
    InMux I__8497 (
            .O(N__34761),
            .I(bfn_15_31_0_));
    InMux I__8496 (
            .O(N__34758),
            .I(N__34755));
    LocalMux I__8495 (
            .O(N__34755),
            .I(n9249));
    InMux I__8494 (
            .O(N__34752),
            .I(N__34748));
    InMux I__8493 (
            .O(N__34751),
            .I(N__34745));
    LocalMux I__8492 (
            .O(N__34748),
            .I(r_Clock_Count_0));
    LocalMux I__8491 (
            .O(N__34745),
            .I(r_Clock_Count_0));
    InMux I__8490 (
            .O(N__34740),
            .I(N__34737));
    LocalMux I__8489 (
            .O(N__34737),
            .I(n9266));
    InMux I__8488 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__8487 (
            .O(N__34731),
            .I(\c0.n900 ));
    CascadeMux I__8486 (
            .O(N__34728),
            .I(N__34725));
    InMux I__8485 (
            .O(N__34725),
            .I(N__34722));
    LocalMux I__8484 (
            .O(N__34722),
            .I(\c0.n22 ));
    InMux I__8483 (
            .O(N__34719),
            .I(N__34715));
    InMux I__8482 (
            .O(N__34718),
            .I(N__34712));
    LocalMux I__8481 (
            .O(N__34715),
            .I(N__34709));
    LocalMux I__8480 (
            .O(N__34712),
            .I(\c0.delay_counter_0 ));
    Odrv4 I__8479 (
            .O(N__34709),
            .I(\c0.delay_counter_0 ));
    InMux I__8478 (
            .O(N__34704),
            .I(N__34701));
    LocalMux I__8477 (
            .O(N__34701),
            .I(\c0.n21_adj_1653 ));
    InMux I__8476 (
            .O(N__34698),
            .I(N__34692));
    InMux I__8475 (
            .O(N__34697),
            .I(N__34692));
    LocalMux I__8474 (
            .O(N__34692),
            .I(\c0.delay_counter_1 ));
    InMux I__8473 (
            .O(N__34689),
            .I(\c0.n8120 ));
    InMux I__8472 (
            .O(N__34686),
            .I(N__34683));
    LocalMux I__8471 (
            .O(N__34683),
            .I(\c0.n20_adj_1652 ));
    InMux I__8470 (
            .O(N__34680),
            .I(N__34674));
    InMux I__8469 (
            .O(N__34679),
            .I(N__34674));
    LocalMux I__8468 (
            .O(N__34674),
            .I(\c0.delay_counter_2 ));
    InMux I__8467 (
            .O(N__34671),
            .I(\c0.n8121 ));
    InMux I__8466 (
            .O(N__34668),
            .I(N__34665));
    LocalMux I__8465 (
            .O(N__34665),
            .I(\c0.tx.n9027 ));
    InMux I__8464 (
            .O(N__34662),
            .I(bfn_15_30_0_));
    CascadeMux I__8463 (
            .O(N__34659),
            .I(N__34654));
    InMux I__8462 (
            .O(N__34658),
            .I(N__34651));
    InMux I__8461 (
            .O(N__34657),
            .I(N__34648));
    InMux I__8460 (
            .O(N__34654),
            .I(N__34645));
    LocalMux I__8459 (
            .O(N__34651),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__8458 (
            .O(N__34648),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__8457 (
            .O(N__34645),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__8456 (
            .O(N__34638),
            .I(N__34635));
    LocalMux I__8455 (
            .O(N__34635),
            .I(\c0.tx.n9290 ));
    InMux I__8454 (
            .O(N__34632),
            .I(\c0.tx.n8090 ));
    InMux I__8453 (
            .O(N__34629),
            .I(N__34624));
    InMux I__8452 (
            .O(N__34628),
            .I(N__34619));
    InMux I__8451 (
            .O(N__34627),
            .I(N__34619));
    LocalMux I__8450 (
            .O(N__34624),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__8449 (
            .O(N__34619),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__8448 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__8447 (
            .O(N__34611),
            .I(\c0.tx.n9313 ));
    InMux I__8446 (
            .O(N__34608),
            .I(\c0.tx.n8091 ));
    InMux I__8445 (
            .O(N__34605),
            .I(N__34600));
    InMux I__8444 (
            .O(N__34604),
            .I(N__34595));
    InMux I__8443 (
            .O(N__34603),
            .I(N__34595));
    LocalMux I__8442 (
            .O(N__34600),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__8441 (
            .O(N__34595),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__8440 (
            .O(N__34590),
            .I(N__34587));
    LocalMux I__8439 (
            .O(N__34587),
            .I(\c0.tx.n9281 ));
    InMux I__8438 (
            .O(N__34584),
            .I(\c0.tx.n8092 ));
    InMux I__8437 (
            .O(N__34581),
            .I(\c0.tx.n8093 ));
    InMux I__8436 (
            .O(N__34578),
            .I(N__34575));
    LocalMux I__8435 (
            .O(N__34575),
            .I(\c0.tx.n9059 ));
    CascadeMux I__8434 (
            .O(N__34572),
            .I(N__34569));
    InMux I__8433 (
            .O(N__34569),
            .I(N__34565));
    CascadeMux I__8432 (
            .O(N__34568),
            .I(N__34562));
    LocalMux I__8431 (
            .O(N__34565),
            .I(N__34559));
    InMux I__8430 (
            .O(N__34562),
            .I(N__34556));
    Span4Mux_h I__8429 (
            .O(N__34559),
            .I(N__34551));
    LocalMux I__8428 (
            .O(N__34556),
            .I(N__34551));
    Odrv4 I__8427 (
            .O(N__34551),
            .I(n28));
    InMux I__8426 (
            .O(N__34548),
            .I(N__34544));
    InMux I__8425 (
            .O(N__34547),
            .I(N__34537));
    LocalMux I__8424 (
            .O(N__34544),
            .I(N__34534));
    InMux I__8423 (
            .O(N__34543),
            .I(N__34531));
    InMux I__8422 (
            .O(N__34542),
            .I(N__34524));
    InMux I__8421 (
            .O(N__34541),
            .I(N__34524));
    InMux I__8420 (
            .O(N__34540),
            .I(N__34524));
    LocalMux I__8419 (
            .O(N__34537),
            .I(\c0.tx_transmit ));
    Odrv4 I__8418 (
            .O(N__34534),
            .I(\c0.tx_transmit ));
    LocalMux I__8417 (
            .O(N__34531),
            .I(\c0.tx_transmit ));
    LocalMux I__8416 (
            .O(N__34524),
            .I(\c0.tx_transmit ));
    CascadeMux I__8415 (
            .O(N__34515),
            .I(n3151_cascade_));
    InMux I__8414 (
            .O(N__34512),
            .I(N__34509));
    LocalMux I__8413 (
            .O(N__34509),
            .I(n11_adj_1752));
    CascadeMux I__8412 (
            .O(N__34506),
            .I(\c0.tx.n5_cascade_ ));
    CascadeMux I__8411 (
            .O(N__34503),
            .I(N__34496));
    CascadeMux I__8410 (
            .O(N__34502),
            .I(N__34493));
    InMux I__8409 (
            .O(N__34501),
            .I(N__34490));
    CascadeMux I__8408 (
            .O(N__34500),
            .I(N__34487));
    CascadeMux I__8407 (
            .O(N__34499),
            .I(N__34480));
    InMux I__8406 (
            .O(N__34496),
            .I(N__34474));
    InMux I__8405 (
            .O(N__34493),
            .I(N__34474));
    LocalMux I__8404 (
            .O(N__34490),
            .I(N__34471));
    InMux I__8403 (
            .O(N__34487),
            .I(N__34468));
    InMux I__8402 (
            .O(N__34486),
            .I(N__34463));
    InMux I__8401 (
            .O(N__34485),
            .I(N__34463));
    InMux I__8400 (
            .O(N__34484),
            .I(N__34454));
    InMux I__8399 (
            .O(N__34483),
            .I(N__34454));
    InMux I__8398 (
            .O(N__34480),
            .I(N__34454));
    InMux I__8397 (
            .O(N__34479),
            .I(N__34454));
    LocalMux I__8396 (
            .O(N__34474),
            .I(r_SM_Main_0));
    Odrv4 I__8395 (
            .O(N__34471),
            .I(r_SM_Main_0));
    LocalMux I__8394 (
            .O(N__34468),
            .I(r_SM_Main_0));
    LocalMux I__8393 (
            .O(N__34463),
            .I(r_SM_Main_0));
    LocalMux I__8392 (
            .O(N__34454),
            .I(r_SM_Main_0));
    CascadeMux I__8391 (
            .O(N__34443),
            .I(\c0.tx.n23_cascade_ ));
    CascadeMux I__8390 (
            .O(N__34440),
            .I(N__34436));
    InMux I__8389 (
            .O(N__34439),
            .I(N__34433));
    InMux I__8388 (
            .O(N__34436),
            .I(N__34430));
    LocalMux I__8387 (
            .O(N__34433),
            .I(N__34414));
    LocalMux I__8386 (
            .O(N__34430),
            .I(N__34414));
    CascadeMux I__8385 (
            .O(N__34429),
            .I(N__34411));
    InMux I__8384 (
            .O(N__34428),
            .I(N__34407));
    InMux I__8383 (
            .O(N__34427),
            .I(N__34404));
    InMux I__8382 (
            .O(N__34426),
            .I(N__34397));
    InMux I__8381 (
            .O(N__34425),
            .I(N__34397));
    InMux I__8380 (
            .O(N__34424),
            .I(N__34397));
    InMux I__8379 (
            .O(N__34423),
            .I(N__34394));
    InMux I__8378 (
            .O(N__34422),
            .I(N__34389));
    InMux I__8377 (
            .O(N__34421),
            .I(N__34389));
    InMux I__8376 (
            .O(N__34420),
            .I(N__34384));
    InMux I__8375 (
            .O(N__34419),
            .I(N__34384));
    Span4Mux_h I__8374 (
            .O(N__34414),
            .I(N__34381));
    InMux I__8373 (
            .O(N__34411),
            .I(N__34376));
    InMux I__8372 (
            .O(N__34410),
            .I(N__34376));
    LocalMux I__8371 (
            .O(N__34407),
            .I(r_SM_Main_1));
    LocalMux I__8370 (
            .O(N__34404),
            .I(r_SM_Main_1));
    LocalMux I__8369 (
            .O(N__34397),
            .I(r_SM_Main_1));
    LocalMux I__8368 (
            .O(N__34394),
            .I(r_SM_Main_1));
    LocalMux I__8367 (
            .O(N__34389),
            .I(r_SM_Main_1));
    LocalMux I__8366 (
            .O(N__34384),
            .I(r_SM_Main_1));
    Odrv4 I__8365 (
            .O(N__34381),
            .I(r_SM_Main_1));
    LocalMux I__8364 (
            .O(N__34376),
            .I(r_SM_Main_1));
    InMux I__8363 (
            .O(N__34359),
            .I(N__34356));
    LocalMux I__8362 (
            .O(N__34356),
            .I(n9259));
    CascadeMux I__8361 (
            .O(N__34353),
            .I(N__34344));
    CascadeMux I__8360 (
            .O(N__34352),
            .I(N__34341));
    InMux I__8359 (
            .O(N__34351),
            .I(N__34329));
    InMux I__8358 (
            .O(N__34350),
            .I(N__34322));
    InMux I__8357 (
            .O(N__34349),
            .I(N__34322));
    InMux I__8356 (
            .O(N__34348),
            .I(N__34322));
    InMux I__8355 (
            .O(N__34347),
            .I(N__34319));
    InMux I__8354 (
            .O(N__34344),
            .I(N__34308));
    InMux I__8353 (
            .O(N__34341),
            .I(N__34308));
    InMux I__8352 (
            .O(N__34340),
            .I(N__34308));
    InMux I__8351 (
            .O(N__34339),
            .I(N__34308));
    InMux I__8350 (
            .O(N__34338),
            .I(N__34308));
    InMux I__8349 (
            .O(N__34337),
            .I(N__34295));
    InMux I__8348 (
            .O(N__34336),
            .I(N__34295));
    InMux I__8347 (
            .O(N__34335),
            .I(N__34295));
    InMux I__8346 (
            .O(N__34334),
            .I(N__34295));
    InMux I__8345 (
            .O(N__34333),
            .I(N__34295));
    InMux I__8344 (
            .O(N__34332),
            .I(N__34295));
    LocalMux I__8343 (
            .O(N__34329),
            .I(\c0.n123 ));
    LocalMux I__8342 (
            .O(N__34322),
            .I(\c0.n123 ));
    LocalMux I__8341 (
            .O(N__34319),
            .I(\c0.n123 ));
    LocalMux I__8340 (
            .O(N__34308),
            .I(\c0.n123 ));
    LocalMux I__8339 (
            .O(N__34295),
            .I(\c0.n123 ));
    InMux I__8338 (
            .O(N__34284),
            .I(N__34268));
    InMux I__8337 (
            .O(N__34283),
            .I(N__34265));
    InMux I__8336 (
            .O(N__34282),
            .I(N__34254));
    InMux I__8335 (
            .O(N__34281),
            .I(N__34254));
    InMux I__8334 (
            .O(N__34280),
            .I(N__34254));
    InMux I__8333 (
            .O(N__34279),
            .I(N__34254));
    InMux I__8332 (
            .O(N__34278),
            .I(N__34254));
    InMux I__8331 (
            .O(N__34277),
            .I(N__34239));
    InMux I__8330 (
            .O(N__34276),
            .I(N__34239));
    InMux I__8329 (
            .O(N__34275),
            .I(N__34239));
    InMux I__8328 (
            .O(N__34274),
            .I(N__34239));
    InMux I__8327 (
            .O(N__34273),
            .I(N__34239));
    InMux I__8326 (
            .O(N__34272),
            .I(N__34239));
    InMux I__8325 (
            .O(N__34271),
            .I(N__34239));
    LocalMux I__8324 (
            .O(N__34268),
            .I(\c0.n7814 ));
    LocalMux I__8323 (
            .O(N__34265),
            .I(\c0.n7814 ));
    LocalMux I__8322 (
            .O(N__34254),
            .I(\c0.n7814 ));
    LocalMux I__8321 (
            .O(N__34239),
            .I(\c0.n7814 ));
    InMux I__8320 (
            .O(N__34230),
            .I(N__34227));
    LocalMux I__8319 (
            .O(N__34227),
            .I(N__34224));
    Odrv4 I__8318 (
            .O(N__34224),
            .I(\c0.n117 ));
    InMux I__8317 (
            .O(N__34221),
            .I(N__34213));
    InMux I__8316 (
            .O(N__34220),
            .I(N__34213));
    InMux I__8315 (
            .O(N__34219),
            .I(N__34208));
    InMux I__8314 (
            .O(N__34218),
            .I(N__34208));
    LocalMux I__8313 (
            .O(N__34213),
            .I(N__34204));
    LocalMux I__8312 (
            .O(N__34208),
            .I(N__34201));
    InMux I__8311 (
            .O(N__34207),
            .I(N__34197));
    Span4Mux_v I__8310 (
            .O(N__34204),
            .I(N__34192));
    Span4Mux_h I__8309 (
            .O(N__34201),
            .I(N__34189));
    InMux I__8308 (
            .O(N__34200),
            .I(N__34186));
    LocalMux I__8307 (
            .O(N__34197),
            .I(N__34183));
    InMux I__8306 (
            .O(N__34196),
            .I(N__34178));
    InMux I__8305 (
            .O(N__34195),
            .I(N__34178));
    Odrv4 I__8304 (
            .O(N__34192),
            .I(n3747));
    Odrv4 I__8303 (
            .O(N__34189),
            .I(n3747));
    LocalMux I__8302 (
            .O(N__34186),
            .I(n3747));
    Odrv4 I__8301 (
            .O(N__34183),
            .I(n3747));
    LocalMux I__8300 (
            .O(N__34178),
            .I(n3747));
    InMux I__8299 (
            .O(N__34167),
            .I(N__34164));
    LocalMux I__8298 (
            .O(N__34164),
            .I(\c0.tx_active_prev ));
    CascadeMux I__8297 (
            .O(N__34161),
            .I(n8749_cascade_));
    InMux I__8296 (
            .O(N__34158),
            .I(N__34150));
    InMux I__8295 (
            .O(N__34157),
            .I(N__34147));
    InMux I__8294 (
            .O(N__34156),
            .I(N__34140));
    InMux I__8293 (
            .O(N__34155),
            .I(N__34140));
    InMux I__8292 (
            .O(N__34154),
            .I(N__34140));
    InMux I__8291 (
            .O(N__34153),
            .I(N__34137));
    LocalMux I__8290 (
            .O(N__34150),
            .I(tx_active));
    LocalMux I__8289 (
            .O(N__34147),
            .I(tx_active));
    LocalMux I__8288 (
            .O(N__34140),
            .I(tx_active));
    LocalMux I__8287 (
            .O(N__34137),
            .I(tx_active));
    CascadeMux I__8286 (
            .O(N__34128),
            .I(\c0.tx.n8_cascade_ ));
    InMux I__8285 (
            .O(N__34125),
            .I(N__34122));
    LocalMux I__8284 (
            .O(N__34122),
            .I(\c0.n19_adj_1664 ));
    IoInMux I__8283 (
            .O(N__34119),
            .I(N__34116));
    LocalMux I__8282 (
            .O(N__34116),
            .I(N__34113));
    Span4Mux_s0_v I__8281 (
            .O(N__34113),
            .I(N__34109));
    InMux I__8280 (
            .O(N__34112),
            .I(N__34106));
    Span4Mux_h I__8279 (
            .O(N__34109),
            .I(N__34101));
    LocalMux I__8278 (
            .O(N__34106),
            .I(N__34101));
    Span4Mux_h I__8277 (
            .O(N__34101),
            .I(N__34098));
    Span4Mux_v I__8276 (
            .O(N__34098),
            .I(N__34094));
    InMux I__8275 (
            .O(N__34097),
            .I(N__34091));
    Odrv4 I__8274 (
            .O(N__34094),
            .I(tx_o_adj_1726));
    LocalMux I__8273 (
            .O(N__34091),
            .I(tx_o_adj_1726));
    InMux I__8272 (
            .O(N__34086),
            .I(N__34083));
    LocalMux I__8271 (
            .O(N__34083),
            .I(n9452));
    CascadeMux I__8270 (
            .O(N__34080),
            .I(N__34076));
    InMux I__8269 (
            .O(N__34079),
            .I(N__34073));
    InMux I__8268 (
            .O(N__34076),
            .I(N__34070));
    LocalMux I__8267 (
            .O(N__34073),
            .I(r_Tx_Data_0));
    LocalMux I__8266 (
            .O(N__34070),
            .I(r_Tx_Data_0));
    InMux I__8265 (
            .O(N__34065),
            .I(N__34062));
    LocalMux I__8264 (
            .O(N__34062),
            .I(n9455));
    InMux I__8263 (
            .O(N__34059),
            .I(N__34056));
    LocalMux I__8262 (
            .O(N__34056),
            .I(tx_data_4_N_keep));
    InMux I__8261 (
            .O(N__34053),
            .I(N__34047));
    InMux I__8260 (
            .O(N__34052),
            .I(N__34047));
    LocalMux I__8259 (
            .O(N__34047),
            .I(r_Tx_Data_4));
    InMux I__8258 (
            .O(N__34044),
            .I(N__34038));
    InMux I__8257 (
            .O(N__34043),
            .I(N__34038));
    LocalMux I__8256 (
            .O(N__34038),
            .I(n9073));
    InMux I__8255 (
            .O(N__34035),
            .I(N__34028));
    InMux I__8254 (
            .O(N__34034),
            .I(N__34025));
    InMux I__8253 (
            .O(N__34033),
            .I(N__34022));
    InMux I__8252 (
            .O(N__34032),
            .I(N__34017));
    InMux I__8251 (
            .O(N__34031),
            .I(N__34017));
    LocalMux I__8250 (
            .O(N__34028),
            .I(r_Bit_Index_0));
    LocalMux I__8249 (
            .O(N__34025),
            .I(r_Bit_Index_0));
    LocalMux I__8248 (
            .O(N__34022),
            .I(r_Bit_Index_0));
    LocalMux I__8247 (
            .O(N__34017),
            .I(r_Bit_Index_0));
    InMux I__8246 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__8245 (
            .O(N__34005),
            .I(N__34000));
    InMux I__8244 (
            .O(N__34004),
            .I(N__33995));
    InMux I__8243 (
            .O(N__34003),
            .I(N__33995));
    Odrv4 I__8242 (
            .O(N__34000),
            .I(n5062));
    LocalMux I__8241 (
            .O(N__33995),
            .I(n5062));
    CascadeMux I__8240 (
            .O(N__33990),
            .I(n9073_cascade_));
    CascadeMux I__8239 (
            .O(N__33987),
            .I(N__33981));
    InMux I__8238 (
            .O(N__33986),
            .I(N__33977));
    InMux I__8237 (
            .O(N__33985),
            .I(N__33974));
    InMux I__8236 (
            .O(N__33984),
            .I(N__33969));
    InMux I__8235 (
            .O(N__33981),
            .I(N__33966));
    InMux I__8234 (
            .O(N__33980),
            .I(N__33963));
    LocalMux I__8233 (
            .O(N__33977),
            .I(N__33958));
    LocalMux I__8232 (
            .O(N__33974),
            .I(N__33958));
    InMux I__8231 (
            .O(N__33973),
            .I(N__33953));
    InMux I__8230 (
            .O(N__33972),
            .I(N__33953));
    LocalMux I__8229 (
            .O(N__33969),
            .I(N__33950));
    LocalMux I__8228 (
            .O(N__33966),
            .I(N__33947));
    LocalMux I__8227 (
            .O(N__33963),
            .I(r_Bit_Index_1));
    Odrv4 I__8226 (
            .O(N__33958),
            .I(r_Bit_Index_1));
    LocalMux I__8225 (
            .O(N__33953),
            .I(r_Bit_Index_1));
    Odrv4 I__8224 (
            .O(N__33950),
            .I(r_Bit_Index_1));
    Odrv4 I__8223 (
            .O(N__33947),
            .I(r_Bit_Index_1));
    CascadeMux I__8222 (
            .O(N__33936),
            .I(N__33933));
    InMux I__8221 (
            .O(N__33933),
            .I(N__33930));
    LocalMux I__8220 (
            .O(N__33930),
            .I(n3892));
    InMux I__8219 (
            .O(N__33927),
            .I(N__33924));
    LocalMux I__8218 (
            .O(N__33924),
            .I(\c0.n18_adj_1662 ));
    CascadeMux I__8217 (
            .O(N__33921),
            .I(N__33914));
    InMux I__8216 (
            .O(N__33920),
            .I(N__33907));
    InMux I__8215 (
            .O(N__33919),
            .I(N__33900));
    InMux I__8214 (
            .O(N__33918),
            .I(N__33900));
    InMux I__8213 (
            .O(N__33917),
            .I(N__33900));
    InMux I__8212 (
            .O(N__33914),
            .I(N__33897));
    InMux I__8211 (
            .O(N__33913),
            .I(N__33893));
    InMux I__8210 (
            .O(N__33912),
            .I(N__33890));
    InMux I__8209 (
            .O(N__33911),
            .I(N__33885));
    InMux I__8208 (
            .O(N__33910),
            .I(N__33885));
    LocalMux I__8207 (
            .O(N__33907),
            .I(N__33878));
    LocalMux I__8206 (
            .O(N__33900),
            .I(N__33878));
    LocalMux I__8205 (
            .O(N__33897),
            .I(N__33878));
    InMux I__8204 (
            .O(N__33896),
            .I(N__33875));
    LocalMux I__8203 (
            .O(N__33893),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__8202 (
            .O(N__33890),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__8201 (
            .O(N__33885),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__8200 (
            .O(N__33878),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__8199 (
            .O(N__33875),
            .I(\c0.byte_transmit_counter_1 ));
    CascadeMux I__8198 (
            .O(N__33864),
            .I(\c0.n7779_cascade_ ));
    InMux I__8197 (
            .O(N__33861),
            .I(N__33857));
    InMux I__8196 (
            .O(N__33860),
            .I(N__33854));
    LocalMux I__8195 (
            .O(N__33857),
            .I(tx_data_1_N_keep));
    LocalMux I__8194 (
            .O(N__33854),
            .I(tx_data_1_N_keep));
    InMux I__8193 (
            .O(N__33849),
            .I(N__33846));
    LocalMux I__8192 (
            .O(N__33846),
            .I(\c0.data_out_6__7__N_973 ));
    InMux I__8191 (
            .O(N__33843),
            .I(N__33839));
    CascadeMux I__8190 (
            .O(N__33842),
            .I(N__33832));
    LocalMux I__8189 (
            .O(N__33839),
            .I(N__33829));
    InMux I__8188 (
            .O(N__33838),
            .I(N__33824));
    InMux I__8187 (
            .O(N__33837),
            .I(N__33824));
    CascadeMux I__8186 (
            .O(N__33836),
            .I(N__33817));
    InMux I__8185 (
            .O(N__33835),
            .I(N__33814));
    InMux I__8184 (
            .O(N__33832),
            .I(N__33811));
    Span4Mux_v I__8183 (
            .O(N__33829),
            .I(N__33806));
    LocalMux I__8182 (
            .O(N__33824),
            .I(N__33806));
    InMux I__8181 (
            .O(N__33823),
            .I(N__33801));
    InMux I__8180 (
            .O(N__33822),
            .I(N__33801));
    InMux I__8179 (
            .O(N__33821),
            .I(N__33796));
    InMux I__8178 (
            .O(N__33820),
            .I(N__33796));
    InMux I__8177 (
            .O(N__33817),
            .I(N__33793));
    LocalMux I__8176 (
            .O(N__33814),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8175 (
            .O(N__33811),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__8174 (
            .O(N__33806),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8173 (
            .O(N__33801),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8172 (
            .O(N__33796),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8171 (
            .O(N__33793),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__8170 (
            .O(N__33780),
            .I(N__33771));
    InMux I__8169 (
            .O(N__33779),
            .I(N__33771));
    InMux I__8168 (
            .O(N__33778),
            .I(N__33767));
    InMux I__8167 (
            .O(N__33777),
            .I(N__33762));
    InMux I__8166 (
            .O(N__33776),
            .I(N__33762));
    LocalMux I__8165 (
            .O(N__33771),
            .I(N__33759));
    InMux I__8164 (
            .O(N__33770),
            .I(N__33755));
    LocalMux I__8163 (
            .O(N__33767),
            .I(N__33750));
    LocalMux I__8162 (
            .O(N__33762),
            .I(N__33750));
    Span4Mux_v I__8161 (
            .O(N__33759),
            .I(N__33747));
    InMux I__8160 (
            .O(N__33758),
            .I(N__33744));
    LocalMux I__8159 (
            .O(N__33755),
            .I(\c0.byte_transmit_counter_4 ));
    Odrv4 I__8158 (
            .O(N__33750),
            .I(\c0.byte_transmit_counter_4 ));
    Odrv4 I__8157 (
            .O(N__33747),
            .I(\c0.byte_transmit_counter_4 ));
    LocalMux I__8156 (
            .O(N__33744),
            .I(\c0.byte_transmit_counter_4 ));
    CascadeMux I__8155 (
            .O(N__33735),
            .I(N__33732));
    InMux I__8154 (
            .O(N__33732),
            .I(N__33728));
    CascadeMux I__8153 (
            .O(N__33731),
            .I(N__33720));
    LocalMux I__8152 (
            .O(N__33728),
            .I(N__33716));
    InMux I__8151 (
            .O(N__33727),
            .I(N__33713));
    InMux I__8150 (
            .O(N__33726),
            .I(N__33706));
    InMux I__8149 (
            .O(N__33725),
            .I(N__33706));
    InMux I__8148 (
            .O(N__33724),
            .I(N__33706));
    InMux I__8147 (
            .O(N__33723),
            .I(N__33701));
    InMux I__8146 (
            .O(N__33720),
            .I(N__33701));
    InMux I__8145 (
            .O(N__33719),
            .I(N__33697));
    Span4Mux_v I__8144 (
            .O(N__33716),
            .I(N__33688));
    LocalMux I__8143 (
            .O(N__33713),
            .I(N__33688));
    LocalMux I__8142 (
            .O(N__33706),
            .I(N__33688));
    LocalMux I__8141 (
            .O(N__33701),
            .I(N__33688));
    InMux I__8140 (
            .O(N__33700),
            .I(N__33685));
    LocalMux I__8139 (
            .O(N__33697),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__8138 (
            .O(N__33688),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__8137 (
            .O(N__33685),
            .I(\c0.byte_transmit_counter_2 ));
    InMux I__8136 (
            .O(N__33678),
            .I(N__33666));
    InMux I__8135 (
            .O(N__33677),
            .I(N__33666));
    InMux I__8134 (
            .O(N__33676),
            .I(N__33666));
    InMux I__8133 (
            .O(N__33675),
            .I(N__33661));
    InMux I__8132 (
            .O(N__33674),
            .I(N__33661));
    InMux I__8131 (
            .O(N__33673),
            .I(N__33657));
    LocalMux I__8130 (
            .O(N__33666),
            .I(N__33654));
    LocalMux I__8129 (
            .O(N__33661),
            .I(N__33651));
    InMux I__8128 (
            .O(N__33660),
            .I(N__33648));
    LocalMux I__8127 (
            .O(N__33657),
            .I(\c0.byte_transmit_counter_3 ));
    Odrv4 I__8126 (
            .O(N__33654),
            .I(\c0.byte_transmit_counter_3 ));
    Odrv4 I__8125 (
            .O(N__33651),
            .I(\c0.byte_transmit_counter_3 ));
    LocalMux I__8124 (
            .O(N__33648),
            .I(\c0.byte_transmit_counter_3 ));
    InMux I__8123 (
            .O(N__33639),
            .I(N__33636));
    LocalMux I__8122 (
            .O(N__33636),
            .I(\c0.n9291 ));
    InMux I__8121 (
            .O(N__33633),
            .I(N__33629));
    InMux I__8120 (
            .O(N__33632),
            .I(N__33626));
    LocalMux I__8119 (
            .O(N__33629),
            .I(N__33623));
    LocalMux I__8118 (
            .O(N__33626),
            .I(r_Tx_Data_3));
    Odrv4 I__8117 (
            .O(N__33623),
            .I(r_Tx_Data_3));
    InMux I__8116 (
            .O(N__33618),
            .I(N__33615));
    LocalMux I__8115 (
            .O(N__33615),
            .I(tx_data_7_N_keep));
    CascadeMux I__8114 (
            .O(N__33612),
            .I(N__33608));
    InMux I__8113 (
            .O(N__33611),
            .I(N__33603));
    InMux I__8112 (
            .O(N__33608),
            .I(N__33603));
    LocalMux I__8111 (
            .O(N__33603),
            .I(r_Tx_Data_7));
    InMux I__8110 (
            .O(N__33600),
            .I(N__33596));
    InMux I__8109 (
            .O(N__33599),
            .I(N__33593));
    LocalMux I__8108 (
            .O(N__33596),
            .I(N__33590));
    LocalMux I__8107 (
            .O(N__33593),
            .I(r_Tx_Data_1));
    Odrv4 I__8106 (
            .O(N__33590),
            .I(r_Tx_Data_1));
    CascadeMux I__8105 (
            .O(N__33585),
            .I(N__33581));
    InMux I__8104 (
            .O(N__33584),
            .I(N__33578));
    InMux I__8103 (
            .O(N__33581),
            .I(N__33575));
    LocalMux I__8102 (
            .O(N__33578),
            .I(r_Tx_Data_5));
    LocalMux I__8101 (
            .O(N__33575),
            .I(r_Tx_Data_5));
    InMux I__8100 (
            .O(N__33570),
            .I(N__33567));
    LocalMux I__8099 (
            .O(N__33567),
            .I(n9710));
    CascadeMux I__8098 (
            .O(N__33564),
            .I(n9713_cascade_));
    CascadeMux I__8097 (
            .O(N__33561),
            .I(n5_cascade_));
    CascadeMux I__8096 (
            .O(N__33558),
            .I(n3_cascade_));
    InMux I__8095 (
            .O(N__33555),
            .I(N__33551));
    InMux I__8094 (
            .O(N__33554),
            .I(N__33548));
    LocalMux I__8093 (
            .O(N__33551),
            .I(\c0.data_out_6_7_N_965_6 ));
    LocalMux I__8092 (
            .O(N__33548),
            .I(\c0.data_out_6_7_N_965_6 ));
    InMux I__8091 (
            .O(N__33543),
            .I(N__33539));
    InMux I__8090 (
            .O(N__33542),
            .I(N__33536));
    LocalMux I__8089 (
            .O(N__33539),
            .I(\c0.data_out_6_7_N_965_4 ));
    LocalMux I__8088 (
            .O(N__33536),
            .I(\c0.data_out_6_7_N_965_4 ));
    InMux I__8087 (
            .O(N__33531),
            .I(N__33527));
    InMux I__8086 (
            .O(N__33530),
            .I(N__33524));
    LocalMux I__8085 (
            .O(N__33527),
            .I(\c0.data_out_6_7_N_965_7 ));
    LocalMux I__8084 (
            .O(N__33524),
            .I(\c0.data_out_6_7_N_965_7 ));
    CascadeMux I__8083 (
            .O(N__33519),
            .I(\c0.n7_cascade_ ));
    InMux I__8082 (
            .O(N__33516),
            .I(N__33513));
    LocalMux I__8081 (
            .O(N__33513),
            .I(\c0.n8 ));
    CascadeMux I__8080 (
            .O(N__33510),
            .I(\c0.n7814_cascade_ ));
    InMux I__8079 (
            .O(N__33507),
            .I(N__33501));
    InMux I__8078 (
            .O(N__33506),
            .I(N__33501));
    LocalMux I__8077 (
            .O(N__33501),
            .I(data_out_6_7_N_965_5));
    CascadeMux I__8076 (
            .O(N__33498),
            .I(n7204_cascade_));
    InMux I__8075 (
            .O(N__33495),
            .I(N__33491));
    InMux I__8074 (
            .O(N__33494),
            .I(N__33488));
    LocalMux I__8073 (
            .O(N__33491),
            .I(byte_transmit_counter_5));
    LocalMux I__8072 (
            .O(N__33488),
            .I(byte_transmit_counter_5));
    InMux I__8071 (
            .O(N__33483),
            .I(N__33477));
    InMux I__8070 (
            .O(N__33482),
            .I(N__33477));
    LocalMux I__8069 (
            .O(N__33477),
            .I(\c0.data_out_6_7_N_965_1 ));
    CascadeMux I__8068 (
            .O(N__33474),
            .I(N__33470));
    InMux I__8067 (
            .O(N__33473),
            .I(N__33466));
    InMux I__8066 (
            .O(N__33470),
            .I(N__33461));
    InMux I__8065 (
            .O(N__33469),
            .I(N__33461));
    LocalMux I__8064 (
            .O(N__33466),
            .I(n7204));
    LocalMux I__8063 (
            .O(N__33461),
            .I(n7204));
    CascadeMux I__8062 (
            .O(N__33456),
            .I(tx_data_1_N_keep_cascade_));
    CascadeMux I__8061 (
            .O(N__33453),
            .I(\c0.n17_adj_1663_cascade_ ));
    CascadeMux I__8060 (
            .O(N__33450),
            .I(\c0.n123_cascade_ ));
    CascadeMux I__8059 (
            .O(N__33447),
            .I(N__33444));
    InMux I__8058 (
            .O(N__33444),
            .I(N__33440));
    InMux I__8057 (
            .O(N__33443),
            .I(N__33437));
    LocalMux I__8056 (
            .O(N__33440),
            .I(\c0.byte_transmit_counter_6 ));
    LocalMux I__8055 (
            .O(N__33437),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__8054 (
            .O(N__33432),
            .I(N__33428));
    InMux I__8053 (
            .O(N__33431),
            .I(N__33425));
    LocalMux I__8052 (
            .O(N__33428),
            .I(\c0.byte_transmit_counter_7 ));
    LocalMux I__8051 (
            .O(N__33425),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__8050 (
            .O(N__33420),
            .I(N__33416));
    InMux I__8049 (
            .O(N__33419),
            .I(N__33413));
    LocalMux I__8048 (
            .O(N__33416),
            .I(\c0.data_out_6_7_N_965_3 ));
    LocalMux I__8047 (
            .O(N__33413),
            .I(\c0.data_out_6_7_N_965_3 ));
    InMux I__8046 (
            .O(N__33408),
            .I(N__33404));
    InMux I__8045 (
            .O(N__33407),
            .I(N__33401));
    LocalMux I__8044 (
            .O(N__33404),
            .I(\c0.data_out_6_7_N_965_2 ));
    LocalMux I__8043 (
            .O(N__33401),
            .I(\c0.data_out_6_7_N_965_2 ));
    CascadeMux I__8042 (
            .O(N__33396),
            .I(N__33392));
    InMux I__8041 (
            .O(N__33395),
            .I(N__33387));
    InMux I__8040 (
            .O(N__33392),
            .I(N__33387));
    LocalMux I__8039 (
            .O(N__33387),
            .I(\c0.data_out_6_7_N_965_0 ));
    CascadeMux I__8038 (
            .O(N__33384),
            .I(tx_data_5_N_keep_cascade_));
    InMux I__8037 (
            .O(N__33381),
            .I(N__33376));
    CascadeMux I__8036 (
            .O(N__33380),
            .I(N__33372));
    CascadeMux I__8035 (
            .O(N__33379),
            .I(N__33369));
    LocalMux I__8034 (
            .O(N__33376),
            .I(N__33366));
    InMux I__8033 (
            .O(N__33375),
            .I(N__33363));
    InMux I__8032 (
            .O(N__33372),
            .I(N__33358));
    InMux I__8031 (
            .O(N__33369),
            .I(N__33358));
    Odrv12 I__8030 (
            .O(N__33366),
            .I(\c0.n11 ));
    LocalMux I__8029 (
            .O(N__33363),
            .I(\c0.n11 ));
    LocalMux I__8028 (
            .O(N__33358),
            .I(\c0.n11 ));
    CascadeMux I__8027 (
            .O(N__33351),
            .I(tx_data_2_N_keep_cascade_));
    InMux I__8026 (
            .O(N__33348),
            .I(N__33345));
    LocalMux I__8025 (
            .O(N__33345),
            .I(tx_data_6_N_keep));
    CascadeMux I__8024 (
            .O(N__33342),
            .I(n8705_cascade_));
    InMux I__8023 (
            .O(N__33339),
            .I(N__33333));
    InMux I__8022 (
            .O(N__33338),
            .I(N__33333));
    LocalMux I__8021 (
            .O(N__33333),
            .I(r_Tx_Data_6));
    InMux I__8020 (
            .O(N__33330),
            .I(N__33324));
    InMux I__8019 (
            .O(N__33329),
            .I(N__33324));
    LocalMux I__8018 (
            .O(N__33324),
            .I(r_Tx_Data_2));
    InMux I__8017 (
            .O(N__33321),
            .I(N__33318));
    LocalMux I__8016 (
            .O(N__33318),
            .I(N__33315));
    Span4Mux_s2_v I__8015 (
            .O(N__33315),
            .I(N__33310));
    InMux I__8014 (
            .O(N__33314),
            .I(N__33307));
    InMux I__8013 (
            .O(N__33313),
            .I(N__33304));
    Span4Mux_h I__8012 (
            .O(N__33310),
            .I(N__33297));
    LocalMux I__8011 (
            .O(N__33307),
            .I(N__33297));
    LocalMux I__8010 (
            .O(N__33304),
            .I(N__33294));
    InMux I__8009 (
            .O(N__33303),
            .I(N__33291));
    InMux I__8008 (
            .O(N__33302),
            .I(N__33288));
    Span4Mux_v I__8007 (
            .O(N__33297),
            .I(N__33285));
    Span4Mux_h I__8006 (
            .O(N__33294),
            .I(N__33280));
    LocalMux I__8005 (
            .O(N__33291),
            .I(N__33280));
    LocalMux I__8004 (
            .O(N__33288),
            .I(data_in_field_132));
    Odrv4 I__8003 (
            .O(N__33285),
            .I(data_in_field_132));
    Odrv4 I__8002 (
            .O(N__33280),
            .I(data_in_field_132));
    InMux I__8001 (
            .O(N__33273),
            .I(N__33270));
    LocalMux I__8000 (
            .O(N__33270),
            .I(N__33267));
    Span4Mux_s2_v I__7999 (
            .O(N__33267),
            .I(N__33264));
    Odrv4 I__7998 (
            .O(N__33264),
            .I(\c0.n9680 ));
    CascadeMux I__7997 (
            .O(N__33261),
            .I(N__33258));
    InMux I__7996 (
            .O(N__33258),
            .I(N__33254));
    CascadeMux I__7995 (
            .O(N__33257),
            .I(N__33251));
    LocalMux I__7994 (
            .O(N__33254),
            .I(N__33248));
    InMux I__7993 (
            .O(N__33251),
            .I(N__33244));
    Span4Mux_h I__7992 (
            .O(N__33248),
            .I(N__33241));
    InMux I__7991 (
            .O(N__33247),
            .I(N__33238));
    LocalMux I__7990 (
            .O(N__33244),
            .I(N__33235));
    Span4Mux_v I__7989 (
            .O(N__33241),
            .I(N__33228));
    LocalMux I__7988 (
            .O(N__33238),
            .I(N__33228));
    Span4Mux_v I__7987 (
            .O(N__33235),
            .I(N__33225));
    InMux I__7986 (
            .O(N__33234),
            .I(N__33220));
    InMux I__7985 (
            .O(N__33233),
            .I(N__33220));
    Span4Mux_h I__7984 (
            .O(N__33228),
            .I(N__33217));
    Odrv4 I__7983 (
            .O(N__33225),
            .I(data_in_field_140));
    LocalMux I__7982 (
            .O(N__33220),
            .I(data_in_field_140));
    Odrv4 I__7981 (
            .O(N__33217),
            .I(data_in_field_140));
    CascadeMux I__7980 (
            .O(N__33210),
            .I(N__33205));
    InMux I__7979 (
            .O(N__33209),
            .I(N__33194));
    InMux I__7978 (
            .O(N__33208),
            .I(N__33194));
    InMux I__7977 (
            .O(N__33205),
            .I(N__33186));
    CascadeMux I__7976 (
            .O(N__33204),
            .I(N__33183));
    CascadeMux I__7975 (
            .O(N__33203),
            .I(N__33178));
    InMux I__7974 (
            .O(N__33202),
            .I(N__33164));
    InMux I__7973 (
            .O(N__33201),
            .I(N__33164));
    InMux I__7972 (
            .O(N__33200),
            .I(N__33164));
    InMux I__7971 (
            .O(N__33199),
            .I(N__33164));
    LocalMux I__7970 (
            .O(N__33194),
            .I(N__33161));
    InMux I__7969 (
            .O(N__33193),
            .I(N__33152));
    InMux I__7968 (
            .O(N__33192),
            .I(N__33152));
    InMux I__7967 (
            .O(N__33191),
            .I(N__33152));
    InMux I__7966 (
            .O(N__33190),
            .I(N__33152));
    InMux I__7965 (
            .O(N__33189),
            .I(N__33145));
    LocalMux I__7964 (
            .O(N__33186),
            .I(N__33142));
    InMux I__7963 (
            .O(N__33183),
            .I(N__33139));
    InMux I__7962 (
            .O(N__33182),
            .I(N__33130));
    InMux I__7961 (
            .O(N__33181),
            .I(N__33130));
    InMux I__7960 (
            .O(N__33178),
            .I(N__33125));
    InMux I__7959 (
            .O(N__33177),
            .I(N__33125));
    InMux I__7958 (
            .O(N__33176),
            .I(N__33122));
    CascadeMux I__7957 (
            .O(N__33175),
            .I(N__33117));
    CascadeMux I__7956 (
            .O(N__33174),
            .I(N__33112));
    InMux I__7955 (
            .O(N__33173),
            .I(N__33109));
    LocalMux I__7954 (
            .O(N__33164),
            .I(N__33102));
    Span4Mux_v I__7953 (
            .O(N__33161),
            .I(N__33102));
    LocalMux I__7952 (
            .O(N__33152),
            .I(N__33102));
    InMux I__7951 (
            .O(N__33151),
            .I(N__33099));
    CascadeMux I__7950 (
            .O(N__33150),
            .I(N__33092));
    InMux I__7949 (
            .O(N__33149),
            .I(N__33085));
    InMux I__7948 (
            .O(N__33148),
            .I(N__33085));
    LocalMux I__7947 (
            .O(N__33145),
            .I(N__33082));
    Span4Mux_h I__7946 (
            .O(N__33142),
            .I(N__33077));
    LocalMux I__7945 (
            .O(N__33139),
            .I(N__33077));
    InMux I__7944 (
            .O(N__33138),
            .I(N__33074));
    InMux I__7943 (
            .O(N__33137),
            .I(N__33071));
    CascadeMux I__7942 (
            .O(N__33136),
            .I(N__33068));
    CascadeMux I__7941 (
            .O(N__33135),
            .I(N__33065));
    LocalMux I__7940 (
            .O(N__33130),
            .I(N__33057));
    LocalMux I__7939 (
            .O(N__33125),
            .I(N__33057));
    LocalMux I__7938 (
            .O(N__33122),
            .I(N__33057));
    InMux I__7937 (
            .O(N__33121),
            .I(N__33054));
    InMux I__7936 (
            .O(N__33120),
            .I(N__33047));
    InMux I__7935 (
            .O(N__33117),
            .I(N__33047));
    InMux I__7934 (
            .O(N__33116),
            .I(N__33047));
    InMux I__7933 (
            .O(N__33115),
            .I(N__33042));
    InMux I__7932 (
            .O(N__33112),
            .I(N__33042));
    LocalMux I__7931 (
            .O(N__33109),
            .I(N__33035));
    Span4Mux_v I__7930 (
            .O(N__33102),
            .I(N__33035));
    LocalMux I__7929 (
            .O(N__33099),
            .I(N__33035));
    CascadeMux I__7928 (
            .O(N__33098),
            .I(N__33025));
    InMux I__7927 (
            .O(N__33097),
            .I(N__33020));
    InMux I__7926 (
            .O(N__33096),
            .I(N__33015));
    InMux I__7925 (
            .O(N__33095),
            .I(N__33009));
    InMux I__7924 (
            .O(N__33092),
            .I(N__33009));
    InMux I__7923 (
            .O(N__33091),
            .I(N__33006));
    CascadeMux I__7922 (
            .O(N__33090),
            .I(N__33003));
    LocalMux I__7921 (
            .O(N__33085),
            .I(N__33000));
    Span4Mux_h I__7920 (
            .O(N__33082),
            .I(N__32995));
    Span4Mux_h I__7919 (
            .O(N__33077),
            .I(N__32995));
    LocalMux I__7918 (
            .O(N__33074),
            .I(N__32992));
    LocalMux I__7917 (
            .O(N__33071),
            .I(N__32989));
    InMux I__7916 (
            .O(N__33068),
            .I(N__32982));
    InMux I__7915 (
            .O(N__33065),
            .I(N__32979));
    InMux I__7914 (
            .O(N__33064),
            .I(N__32975));
    Span4Mux_v I__7913 (
            .O(N__33057),
            .I(N__32966));
    LocalMux I__7912 (
            .O(N__33054),
            .I(N__32966));
    LocalMux I__7911 (
            .O(N__33047),
            .I(N__32966));
    LocalMux I__7910 (
            .O(N__33042),
            .I(N__32966));
    Span4Mux_v I__7909 (
            .O(N__33035),
            .I(N__32963));
    InMux I__7908 (
            .O(N__33034),
            .I(N__32958));
    InMux I__7907 (
            .O(N__33033),
            .I(N__32958));
    CascadeMux I__7906 (
            .O(N__33032),
            .I(N__32952));
    CascadeMux I__7905 (
            .O(N__33031),
            .I(N__32949));
    InMux I__7904 (
            .O(N__33030),
            .I(N__32936));
    InMux I__7903 (
            .O(N__33029),
            .I(N__32936));
    InMux I__7902 (
            .O(N__33028),
            .I(N__32936));
    InMux I__7901 (
            .O(N__33025),
            .I(N__32936));
    CascadeMux I__7900 (
            .O(N__33024),
            .I(N__32933));
    InMux I__7899 (
            .O(N__33023),
            .I(N__32930));
    LocalMux I__7898 (
            .O(N__33020),
            .I(N__32927));
    InMux I__7897 (
            .O(N__33019),
            .I(N__32922));
    InMux I__7896 (
            .O(N__33018),
            .I(N__32922));
    LocalMux I__7895 (
            .O(N__33015),
            .I(N__32919));
    CascadeMux I__7894 (
            .O(N__33014),
            .I(N__32915));
    LocalMux I__7893 (
            .O(N__33009),
            .I(N__32912));
    LocalMux I__7892 (
            .O(N__33006),
            .I(N__32909));
    InMux I__7891 (
            .O(N__33003),
            .I(N__32906));
    Span4Mux_h I__7890 (
            .O(N__33000),
            .I(N__32899));
    Span4Mux_v I__7889 (
            .O(N__32995),
            .I(N__32899));
    Span4Mux_h I__7888 (
            .O(N__32992),
            .I(N__32899));
    Span4Mux_s3_h I__7887 (
            .O(N__32989),
            .I(N__32896));
    InMux I__7886 (
            .O(N__32988),
            .I(N__32893));
    CascadeMux I__7885 (
            .O(N__32987),
            .I(N__32886));
    InMux I__7884 (
            .O(N__32986),
            .I(N__32878));
    InMux I__7883 (
            .O(N__32985),
            .I(N__32878));
    LocalMux I__7882 (
            .O(N__32982),
            .I(N__32873));
    LocalMux I__7881 (
            .O(N__32979),
            .I(N__32873));
    InMux I__7880 (
            .O(N__32978),
            .I(N__32867));
    LocalMux I__7879 (
            .O(N__32975),
            .I(N__32860));
    Span4Mux_v I__7878 (
            .O(N__32966),
            .I(N__32860));
    IoSpan4Mux I__7877 (
            .O(N__32963),
            .I(N__32860));
    LocalMux I__7876 (
            .O(N__32958),
            .I(N__32857));
    InMux I__7875 (
            .O(N__32957),
            .I(N__32852));
    InMux I__7874 (
            .O(N__32956),
            .I(N__32852));
    InMux I__7873 (
            .O(N__32955),
            .I(N__32843));
    InMux I__7872 (
            .O(N__32952),
            .I(N__32843));
    InMux I__7871 (
            .O(N__32949),
            .I(N__32840));
    InMux I__7870 (
            .O(N__32948),
            .I(N__32835));
    InMux I__7869 (
            .O(N__32947),
            .I(N__32835));
    InMux I__7868 (
            .O(N__32946),
            .I(N__32832));
    InMux I__7867 (
            .O(N__32945),
            .I(N__32829));
    LocalMux I__7866 (
            .O(N__32936),
            .I(N__32826));
    InMux I__7865 (
            .O(N__32933),
            .I(N__32823));
    LocalMux I__7864 (
            .O(N__32930),
            .I(N__32820));
    Span4Mux_h I__7863 (
            .O(N__32927),
            .I(N__32815));
    LocalMux I__7862 (
            .O(N__32922),
            .I(N__32815));
    Span4Mux_h I__7861 (
            .O(N__32919),
            .I(N__32812));
    InMux I__7860 (
            .O(N__32918),
            .I(N__32807));
    InMux I__7859 (
            .O(N__32915),
            .I(N__32807));
    Span4Mux_v I__7858 (
            .O(N__32912),
            .I(N__32799));
    Span4Mux_v I__7857 (
            .O(N__32909),
            .I(N__32799));
    LocalMux I__7856 (
            .O(N__32906),
            .I(N__32799));
    IoSpan4Mux I__7855 (
            .O(N__32899),
            .I(N__32796));
    Span4Mux_h I__7854 (
            .O(N__32896),
            .I(N__32791));
    LocalMux I__7853 (
            .O(N__32893),
            .I(N__32791));
    InMux I__7852 (
            .O(N__32892),
            .I(N__32786));
    InMux I__7851 (
            .O(N__32891),
            .I(N__32783));
    InMux I__7850 (
            .O(N__32890),
            .I(N__32780));
    InMux I__7849 (
            .O(N__32889),
            .I(N__32775));
    InMux I__7848 (
            .O(N__32886),
            .I(N__32775));
    InMux I__7847 (
            .O(N__32885),
            .I(N__32770));
    InMux I__7846 (
            .O(N__32884),
            .I(N__32770));
    InMux I__7845 (
            .O(N__32883),
            .I(N__32767));
    LocalMux I__7844 (
            .O(N__32878),
            .I(N__32764));
    Span4Mux_h I__7843 (
            .O(N__32873),
            .I(N__32761));
    InMux I__7842 (
            .O(N__32872),
            .I(N__32758));
    InMux I__7841 (
            .O(N__32871),
            .I(N__32755));
    InMux I__7840 (
            .O(N__32870),
            .I(N__32752));
    LocalMux I__7839 (
            .O(N__32867),
            .I(N__32749));
    Span4Mux_s2_h I__7838 (
            .O(N__32860),
            .I(N__32742));
    Span4Mux_s2_h I__7837 (
            .O(N__32857),
            .I(N__32742));
    LocalMux I__7836 (
            .O(N__32852),
            .I(N__32742));
    InMux I__7835 (
            .O(N__32851),
            .I(N__32733));
    InMux I__7834 (
            .O(N__32850),
            .I(N__32733));
    InMux I__7833 (
            .O(N__32849),
            .I(N__32733));
    InMux I__7832 (
            .O(N__32848),
            .I(N__32733));
    LocalMux I__7831 (
            .O(N__32843),
            .I(N__32728));
    LocalMux I__7830 (
            .O(N__32840),
            .I(N__32728));
    LocalMux I__7829 (
            .O(N__32835),
            .I(N__32709));
    LocalMux I__7828 (
            .O(N__32832),
            .I(N__32709));
    LocalMux I__7827 (
            .O(N__32829),
            .I(N__32709));
    Span4Mux_s1_v I__7826 (
            .O(N__32826),
            .I(N__32709));
    LocalMux I__7825 (
            .O(N__32823),
            .I(N__32709));
    Span4Mux_h I__7824 (
            .O(N__32820),
            .I(N__32709));
    Span4Mux_h I__7823 (
            .O(N__32815),
            .I(N__32709));
    Span4Mux_h I__7822 (
            .O(N__32812),
            .I(N__32709));
    LocalMux I__7821 (
            .O(N__32807),
            .I(N__32709));
    InMux I__7820 (
            .O(N__32806),
            .I(N__32706));
    Span4Mux_h I__7819 (
            .O(N__32799),
            .I(N__32699));
    Span4Mux_s2_v I__7818 (
            .O(N__32796),
            .I(N__32699));
    Span4Mux_h I__7817 (
            .O(N__32791),
            .I(N__32699));
    InMux I__7816 (
            .O(N__32790),
            .I(N__32696));
    InMux I__7815 (
            .O(N__32789),
            .I(N__32693));
    LocalMux I__7814 (
            .O(N__32786),
            .I(N__32678));
    LocalMux I__7813 (
            .O(N__32783),
            .I(N__32678));
    LocalMux I__7812 (
            .O(N__32780),
            .I(N__32678));
    LocalMux I__7811 (
            .O(N__32775),
            .I(N__32678));
    LocalMux I__7810 (
            .O(N__32770),
            .I(N__32678));
    LocalMux I__7809 (
            .O(N__32767),
            .I(N__32678));
    Span12Mux_s1_h I__7808 (
            .O(N__32764),
            .I(N__32678));
    Span4Mux_v I__7807 (
            .O(N__32761),
            .I(N__32675));
    LocalMux I__7806 (
            .O(N__32758),
            .I(N__32668));
    LocalMux I__7805 (
            .O(N__32755),
            .I(N__32668));
    LocalMux I__7804 (
            .O(N__32752),
            .I(N__32668));
    Span4Mux_h I__7803 (
            .O(N__32749),
            .I(N__32663));
    Span4Mux_h I__7802 (
            .O(N__32742),
            .I(N__32663));
    LocalMux I__7801 (
            .O(N__32733),
            .I(N__32656));
    Span12Mux_s6_h I__7800 (
            .O(N__32728),
            .I(N__32656));
    Sp12to4 I__7799 (
            .O(N__32709),
            .I(N__32656));
    LocalMux I__7798 (
            .O(N__32706),
            .I(N__32653));
    Span4Mux_v I__7797 (
            .O(N__32699),
            .I(N__32650));
    LocalMux I__7796 (
            .O(N__32696),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__7795 (
            .O(N__32693),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__7794 (
            .O(N__32678),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7793 (
            .O(N__32675),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7792 (
            .O(N__32668),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7791 (
            .O(N__32663),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__7790 (
            .O(N__32656),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7789 (
            .O(N__32653),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7788 (
            .O(N__32650),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__7787 (
            .O(N__32631),
            .I(N__32628));
    LocalMux I__7786 (
            .O(N__32628),
            .I(N__32625));
    Span4Mux_h I__7785 (
            .O(N__32625),
            .I(N__32622));
    Odrv4 I__7784 (
            .O(N__32622),
            .I(\c0.n9683 ));
    CascadeMux I__7783 (
            .O(N__32619),
            .I(\c0.n11_cascade_ ));
    CascadeMux I__7782 (
            .O(N__32616),
            .I(tx_data_3_N_keep_cascade_));
    InMux I__7781 (
            .O(N__32613),
            .I(N__32610));
    LocalMux I__7780 (
            .O(N__32610),
            .I(tx_data_0_N_keep));
    InMux I__7779 (
            .O(N__32607),
            .I(N__32603));
    InMux I__7778 (
            .O(N__32606),
            .I(N__32600));
    LocalMux I__7777 (
            .O(N__32603),
            .I(N__32595));
    LocalMux I__7776 (
            .O(N__32600),
            .I(N__32592));
    InMux I__7775 (
            .O(N__32599),
            .I(N__32587));
    InMux I__7774 (
            .O(N__32598),
            .I(N__32587));
    Span4Mux_h I__7773 (
            .O(N__32595),
            .I(N__32583));
    Span4Mux_h I__7772 (
            .O(N__32592),
            .I(N__32580));
    LocalMux I__7771 (
            .O(N__32587),
            .I(N__32577));
    InMux I__7770 (
            .O(N__32586),
            .I(N__32574));
    Span4Mux_h I__7769 (
            .O(N__32583),
            .I(N__32571));
    Span4Mux_v I__7768 (
            .O(N__32580),
            .I(N__32568));
    Span4Mux_h I__7767 (
            .O(N__32577),
            .I(N__32565));
    LocalMux I__7766 (
            .O(N__32574),
            .I(data_in_field_133));
    Odrv4 I__7765 (
            .O(N__32571),
            .I(data_in_field_133));
    Odrv4 I__7764 (
            .O(N__32568),
            .I(data_in_field_133));
    Odrv4 I__7763 (
            .O(N__32565),
            .I(data_in_field_133));
    InMux I__7762 (
            .O(N__32556),
            .I(N__32551));
    CascadeMux I__7761 (
            .O(N__32555),
            .I(N__32548));
    InMux I__7760 (
            .O(N__32554),
            .I(N__32545));
    LocalMux I__7759 (
            .O(N__32551),
            .I(N__32542));
    InMux I__7758 (
            .O(N__32548),
            .I(N__32539));
    LocalMux I__7757 (
            .O(N__32545),
            .I(N__32533));
    Span4Mux_h I__7756 (
            .O(N__32542),
            .I(N__32533));
    LocalMux I__7755 (
            .O(N__32539),
            .I(N__32530));
    InMux I__7754 (
            .O(N__32538),
            .I(N__32527));
    Span4Mux_h I__7753 (
            .O(N__32533),
            .I(N__32524));
    Span4Mux_h I__7752 (
            .O(N__32530),
            .I(N__32521));
    LocalMux I__7751 (
            .O(N__32527),
            .I(data_in_field_103));
    Odrv4 I__7750 (
            .O(N__32524),
            .I(data_in_field_103));
    Odrv4 I__7749 (
            .O(N__32521),
            .I(data_in_field_103));
    InMux I__7748 (
            .O(N__32514),
            .I(N__32510));
    InMux I__7747 (
            .O(N__32513),
            .I(N__32504));
    LocalMux I__7746 (
            .O(N__32510),
            .I(N__32501));
    InMux I__7745 (
            .O(N__32509),
            .I(N__32498));
    InMux I__7744 (
            .O(N__32508),
            .I(N__32494));
    InMux I__7743 (
            .O(N__32507),
            .I(N__32491));
    LocalMux I__7742 (
            .O(N__32504),
            .I(N__32488));
    Span4Mux_h I__7741 (
            .O(N__32501),
            .I(N__32485));
    LocalMux I__7740 (
            .O(N__32498),
            .I(N__32482));
    InMux I__7739 (
            .O(N__32497),
            .I(N__32479));
    LocalMux I__7738 (
            .O(N__32494),
            .I(N__32474));
    LocalMux I__7737 (
            .O(N__32491),
            .I(N__32474));
    Span4Mux_h I__7736 (
            .O(N__32488),
            .I(N__32471));
    Span4Mux_v I__7735 (
            .O(N__32485),
            .I(N__32466));
    Span4Mux_h I__7734 (
            .O(N__32482),
            .I(N__32466));
    LocalMux I__7733 (
            .O(N__32479),
            .I(data_in_field_148));
    Odrv12 I__7732 (
            .O(N__32474),
            .I(data_in_field_148));
    Odrv4 I__7731 (
            .O(N__32471),
            .I(data_in_field_148));
    Odrv4 I__7730 (
            .O(N__32466),
            .I(data_in_field_148));
    InMux I__7729 (
            .O(N__32457),
            .I(N__32454));
    LocalMux I__7728 (
            .O(N__32454),
            .I(N__32451));
    Span4Mux_v I__7727 (
            .O(N__32451),
            .I(N__32448));
    Span4Mux_h I__7726 (
            .O(N__32448),
            .I(N__32444));
    InMux I__7725 (
            .O(N__32447),
            .I(N__32441));
    Span4Mux_h I__7724 (
            .O(N__32444),
            .I(N__32436));
    LocalMux I__7723 (
            .O(N__32441),
            .I(N__32436));
    Span4Mux_v I__7722 (
            .O(N__32436),
            .I(N__32433));
    Odrv4 I__7721 (
            .O(N__32433),
            .I(\c0.n8986 ));
    InMux I__7720 (
            .O(N__32430),
            .I(N__32427));
    LocalMux I__7719 (
            .O(N__32427),
            .I(\c0.n45_adj_1656 ));
    InMux I__7718 (
            .O(N__32424),
            .I(\c0.n8083 ));
    InMux I__7717 (
            .O(N__32421),
            .I(\c0.n8084 ));
    InMux I__7716 (
            .O(N__32418),
            .I(\c0.n8085 ));
    InMux I__7715 (
            .O(N__32415),
            .I(\c0.n8086 ));
    InMux I__7714 (
            .O(N__32412),
            .I(\c0.n8087 ));
    InMux I__7713 (
            .O(N__32409),
            .I(\c0.n8088 ));
    InMux I__7712 (
            .O(N__32406),
            .I(\c0.n8089 ));
    InMux I__7711 (
            .O(N__32403),
            .I(N__32400));
    LocalMux I__7710 (
            .O(N__32400),
            .I(N__32397));
    Span4Mux_h I__7709 (
            .O(N__32397),
            .I(N__32394));
    Odrv4 I__7708 (
            .O(N__32394),
            .I(\c0.n22_adj_1681 ));
    CascadeMux I__7707 (
            .O(N__32391),
            .I(\c0.n9491_cascade_ ));
    InMux I__7706 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__7705 (
            .O(N__32385),
            .I(N__32378));
    InMux I__7704 (
            .O(N__32384),
            .I(N__32374));
    InMux I__7703 (
            .O(N__32383),
            .I(N__32371));
    InMux I__7702 (
            .O(N__32382),
            .I(N__32368));
    InMux I__7701 (
            .O(N__32381),
            .I(N__32365));
    Span4Mux_s3_v I__7700 (
            .O(N__32378),
            .I(N__32362));
    InMux I__7699 (
            .O(N__32377),
            .I(N__32359));
    LocalMux I__7698 (
            .O(N__32374),
            .I(N__32356));
    LocalMux I__7697 (
            .O(N__32371),
            .I(N__32353));
    LocalMux I__7696 (
            .O(N__32368),
            .I(N__32350));
    LocalMux I__7695 (
            .O(N__32365),
            .I(N__32345));
    Sp12to4 I__7694 (
            .O(N__32362),
            .I(N__32339));
    LocalMux I__7693 (
            .O(N__32359),
            .I(N__32339));
    Span4Mux_h I__7692 (
            .O(N__32356),
            .I(N__32332));
    Span4Mux_s1_v I__7691 (
            .O(N__32353),
            .I(N__32332));
    Span4Mux_h I__7690 (
            .O(N__32350),
            .I(N__32332));
    InMux I__7689 (
            .O(N__32349),
            .I(N__32329));
    InMux I__7688 (
            .O(N__32348),
            .I(N__32326));
    Span4Mux_v I__7687 (
            .O(N__32345),
            .I(N__32323));
    InMux I__7686 (
            .O(N__32344),
            .I(N__32320));
    Span12Mux_s6_h I__7685 (
            .O(N__32339),
            .I(N__32310));
    Sp12to4 I__7684 (
            .O(N__32332),
            .I(N__32310));
    LocalMux I__7683 (
            .O(N__32329),
            .I(N__32310));
    LocalMux I__7682 (
            .O(N__32326),
            .I(N__32310));
    Sp12to4 I__7681 (
            .O(N__32323),
            .I(N__32305));
    LocalMux I__7680 (
            .O(N__32320),
            .I(N__32305));
    InMux I__7679 (
            .O(N__32319),
            .I(N__32302));
    Span12Mux_s3_v I__7678 (
            .O(N__32310),
            .I(N__32299));
    Odrv12 I__7677 (
            .O(N__32305),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__7676 (
            .O(N__32302),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv12 I__7675 (
            .O(N__32299),
            .I(\c0.byte_transmit_counter2_4 ));
    InMux I__7674 (
            .O(N__32292),
            .I(N__32289));
    LocalMux I__7673 (
            .O(N__32289),
            .I(N__32286));
    Sp12to4 I__7672 (
            .O(N__32286),
            .I(N__32283));
    Span12Mux_s6_v I__7671 (
            .O(N__32283),
            .I(N__32280));
    Odrv12 I__7670 (
            .O(N__32280),
            .I(\c0.tx2.r_Tx_Data_2 ));
    CEMux I__7669 (
            .O(N__32277),
            .I(N__32274));
    LocalMux I__7668 (
            .O(N__32274),
            .I(N__32268));
    CEMux I__7667 (
            .O(N__32273),
            .I(N__32265));
    CEMux I__7666 (
            .O(N__32272),
            .I(N__32261));
    CEMux I__7665 (
            .O(N__32271),
            .I(N__32258));
    IoSpan4Mux I__7664 (
            .O(N__32268),
            .I(N__32255));
    LocalMux I__7663 (
            .O(N__32265),
            .I(N__32252));
    CEMux I__7662 (
            .O(N__32264),
            .I(N__32249));
    LocalMux I__7661 (
            .O(N__32261),
            .I(N__32246));
    LocalMux I__7660 (
            .O(N__32258),
            .I(N__32243));
    Span4Mux_s0_v I__7659 (
            .O(N__32255),
            .I(N__32240));
    Span4Mux_v I__7658 (
            .O(N__32252),
            .I(N__32237));
    LocalMux I__7657 (
            .O(N__32249),
            .I(N__32234));
    Span4Mux_v I__7656 (
            .O(N__32246),
            .I(N__32230));
    Span4Mux_v I__7655 (
            .O(N__32243),
            .I(N__32225));
    Span4Mux_h I__7654 (
            .O(N__32240),
            .I(N__32218));
    Span4Mux_s1_h I__7653 (
            .O(N__32237),
            .I(N__32218));
    Span4Mux_v I__7652 (
            .O(N__32234),
            .I(N__32218));
    CEMux I__7651 (
            .O(N__32233),
            .I(N__32215));
    Span4Mux_v I__7650 (
            .O(N__32230),
            .I(N__32212));
    CEMux I__7649 (
            .O(N__32229),
            .I(N__32209));
    CEMux I__7648 (
            .O(N__32228),
            .I(N__32206));
    Span4Mux_v I__7647 (
            .O(N__32225),
            .I(N__32203));
    Span4Mux_h I__7646 (
            .O(N__32218),
            .I(N__32198));
    LocalMux I__7645 (
            .O(N__32215),
            .I(N__32198));
    Span4Mux_h I__7644 (
            .O(N__32212),
            .I(N__32193));
    LocalMux I__7643 (
            .O(N__32209),
            .I(N__32193));
    LocalMux I__7642 (
            .O(N__32206),
            .I(N__32190));
    Sp12to4 I__7641 (
            .O(N__32203),
            .I(N__32185));
    Sp12to4 I__7640 (
            .O(N__32198),
            .I(N__32185));
    Span4Mux_h I__7639 (
            .O(N__32193),
            .I(N__32182));
    Sp12to4 I__7638 (
            .O(N__32190),
            .I(N__32179));
    Odrv12 I__7637 (
            .O(N__32185),
            .I(\c0.tx2.n3760 ));
    Odrv4 I__7636 (
            .O(N__32182),
            .I(\c0.tx2.n3760 ));
    Odrv12 I__7635 (
            .O(N__32179),
            .I(\c0.tx2.n3760 ));
    InMux I__7634 (
            .O(N__32172),
            .I(N__32168));
    InMux I__7633 (
            .O(N__32171),
            .I(N__32165));
    LocalMux I__7632 (
            .O(N__32168),
            .I(N__32161));
    LocalMux I__7631 (
            .O(N__32165),
            .I(N__32155));
    InMux I__7630 (
            .O(N__32164),
            .I(N__32152));
    Span4Mux_v I__7629 (
            .O(N__32161),
            .I(N__32149));
    InMux I__7628 (
            .O(N__32160),
            .I(N__32146));
    InMux I__7627 (
            .O(N__32159),
            .I(N__32143));
    InMux I__7626 (
            .O(N__32158),
            .I(N__32140));
    Span4Mux_h I__7625 (
            .O(N__32155),
            .I(N__32137));
    LocalMux I__7624 (
            .O(N__32152),
            .I(N__32128));
    Sp12to4 I__7623 (
            .O(N__32149),
            .I(N__32128));
    LocalMux I__7622 (
            .O(N__32146),
            .I(N__32128));
    LocalMux I__7621 (
            .O(N__32143),
            .I(N__32128));
    LocalMux I__7620 (
            .O(N__32140),
            .I(data_in_field_82));
    Odrv4 I__7619 (
            .O(N__32137),
            .I(data_in_field_82));
    Odrv12 I__7618 (
            .O(N__32128),
            .I(data_in_field_82));
    InMux I__7617 (
            .O(N__32121),
            .I(N__32113));
    CascadeMux I__7616 (
            .O(N__32120),
            .I(N__32110));
    InMux I__7615 (
            .O(N__32119),
            .I(N__32105));
    InMux I__7614 (
            .O(N__32118),
            .I(N__32105));
    InMux I__7613 (
            .O(N__32117),
            .I(N__32101));
    InMux I__7612 (
            .O(N__32116),
            .I(N__32098));
    LocalMux I__7611 (
            .O(N__32113),
            .I(N__32095));
    InMux I__7610 (
            .O(N__32110),
            .I(N__32092));
    LocalMux I__7609 (
            .O(N__32105),
            .I(N__32089));
    InMux I__7608 (
            .O(N__32104),
            .I(N__32086));
    LocalMux I__7607 (
            .O(N__32101),
            .I(N__32081));
    LocalMux I__7606 (
            .O(N__32098),
            .I(N__32081));
    Span4Mux_s2_v I__7605 (
            .O(N__32095),
            .I(N__32078));
    LocalMux I__7604 (
            .O(N__32092),
            .I(N__32075));
    Span4Mux_h I__7603 (
            .O(N__32089),
            .I(N__32072));
    LocalMux I__7602 (
            .O(N__32086),
            .I(N__32063));
    Span4Mux_v I__7601 (
            .O(N__32081),
            .I(N__32063));
    Span4Mux_v I__7600 (
            .O(N__32078),
            .I(N__32063));
    Span4Mux_h I__7599 (
            .O(N__32075),
            .I(N__32063));
    Odrv4 I__7598 (
            .O(N__32072),
            .I(data_in_field_90));
    Odrv4 I__7597 (
            .O(N__32063),
            .I(data_in_field_90));
    InMux I__7596 (
            .O(N__32058),
            .I(N__32047));
    InMux I__7595 (
            .O(N__32057),
            .I(N__32047));
    InMux I__7594 (
            .O(N__32056),
            .I(N__32027));
    InMux I__7593 (
            .O(N__32055),
            .I(N__32022));
    InMux I__7592 (
            .O(N__32054),
            .I(N__32022));
    InMux I__7591 (
            .O(N__32053),
            .I(N__32017));
    InMux I__7590 (
            .O(N__32052),
            .I(N__32017));
    LocalMux I__7589 (
            .O(N__32047),
            .I(N__32008));
    InMux I__7588 (
            .O(N__32046),
            .I(N__32004));
    InMux I__7587 (
            .O(N__32045),
            .I(N__32001));
    InMux I__7586 (
            .O(N__32044),
            .I(N__31997));
    InMux I__7585 (
            .O(N__32043),
            .I(N__31994));
    InMux I__7584 (
            .O(N__32042),
            .I(N__31987));
    InMux I__7583 (
            .O(N__32041),
            .I(N__31987));
    InMux I__7582 (
            .O(N__32040),
            .I(N__31984));
    InMux I__7581 (
            .O(N__32039),
            .I(N__31981));
    InMux I__7580 (
            .O(N__32038),
            .I(N__31978));
    InMux I__7579 (
            .O(N__32037),
            .I(N__31972));
    CascadeMux I__7578 (
            .O(N__32036),
            .I(N__31968));
    CascadeMux I__7577 (
            .O(N__32035),
            .I(N__31964));
    InMux I__7576 (
            .O(N__32034),
            .I(N__31961));
    InMux I__7575 (
            .O(N__32033),
            .I(N__31956));
    InMux I__7574 (
            .O(N__32032),
            .I(N__31956));
    InMux I__7573 (
            .O(N__32031),
            .I(N__31953));
    InMux I__7572 (
            .O(N__32030),
            .I(N__31949));
    LocalMux I__7571 (
            .O(N__32027),
            .I(N__31946));
    LocalMux I__7570 (
            .O(N__32022),
            .I(N__31943));
    LocalMux I__7569 (
            .O(N__32017),
            .I(N__31940));
    InMux I__7568 (
            .O(N__32016),
            .I(N__31937));
    InMux I__7567 (
            .O(N__32015),
            .I(N__31934));
    InMux I__7566 (
            .O(N__32014),
            .I(N__31931));
    InMux I__7565 (
            .O(N__32013),
            .I(N__31928));
    InMux I__7564 (
            .O(N__32012),
            .I(N__31923));
    InMux I__7563 (
            .O(N__32011),
            .I(N__31923));
    Span4Mux_s3_v I__7562 (
            .O(N__32008),
            .I(N__31920));
    InMux I__7561 (
            .O(N__32007),
            .I(N__31917));
    LocalMux I__7560 (
            .O(N__32004),
            .I(N__31914));
    LocalMux I__7559 (
            .O(N__32001),
            .I(N__31911));
    InMux I__7558 (
            .O(N__32000),
            .I(N__31907));
    LocalMux I__7557 (
            .O(N__31997),
            .I(N__31904));
    LocalMux I__7556 (
            .O(N__31994),
            .I(N__31901));
    InMux I__7555 (
            .O(N__31993),
            .I(N__31898));
    InMux I__7554 (
            .O(N__31992),
            .I(N__31894));
    LocalMux I__7553 (
            .O(N__31987),
            .I(N__31889));
    LocalMux I__7552 (
            .O(N__31984),
            .I(N__31889));
    LocalMux I__7551 (
            .O(N__31981),
            .I(N__31884));
    LocalMux I__7550 (
            .O(N__31978),
            .I(N__31884));
    InMux I__7549 (
            .O(N__31977),
            .I(N__31881));
    InMux I__7548 (
            .O(N__31976),
            .I(N__31878));
    InMux I__7547 (
            .O(N__31975),
            .I(N__31875));
    LocalMux I__7546 (
            .O(N__31972),
            .I(N__31872));
    CascadeMux I__7545 (
            .O(N__31971),
            .I(N__31869));
    InMux I__7544 (
            .O(N__31968),
            .I(N__31866));
    InMux I__7543 (
            .O(N__31967),
            .I(N__31863));
    InMux I__7542 (
            .O(N__31964),
            .I(N__31860));
    LocalMux I__7541 (
            .O(N__31961),
            .I(N__31853));
    LocalMux I__7540 (
            .O(N__31956),
            .I(N__31853));
    LocalMux I__7539 (
            .O(N__31953),
            .I(N__31853));
    InMux I__7538 (
            .O(N__31952),
            .I(N__31850));
    LocalMux I__7537 (
            .O(N__31949),
            .I(N__31837));
    Span4Mux_h I__7536 (
            .O(N__31946),
            .I(N__31837));
    Span4Mux_s1_v I__7535 (
            .O(N__31943),
            .I(N__31837));
    Span4Mux_s1_v I__7534 (
            .O(N__31940),
            .I(N__31837));
    LocalMux I__7533 (
            .O(N__31937),
            .I(N__31837));
    LocalMux I__7532 (
            .O(N__31934),
            .I(N__31837));
    LocalMux I__7531 (
            .O(N__31931),
            .I(N__31834));
    LocalMux I__7530 (
            .O(N__31928),
            .I(N__31829));
    LocalMux I__7529 (
            .O(N__31923),
            .I(N__31829));
    Span4Mux_h I__7528 (
            .O(N__31920),
            .I(N__31820));
    LocalMux I__7527 (
            .O(N__31917),
            .I(N__31820));
    Span4Mux_s3_v I__7526 (
            .O(N__31914),
            .I(N__31820));
    Span4Mux_s3_v I__7525 (
            .O(N__31911),
            .I(N__31820));
    InMux I__7524 (
            .O(N__31910),
            .I(N__31817));
    LocalMux I__7523 (
            .O(N__31907),
            .I(N__31814));
    Span4Mux_v I__7522 (
            .O(N__31904),
            .I(N__31807));
    Span4Mux_h I__7521 (
            .O(N__31901),
            .I(N__31807));
    LocalMux I__7520 (
            .O(N__31898),
            .I(N__31807));
    InMux I__7519 (
            .O(N__31897),
            .I(N__31804));
    LocalMux I__7518 (
            .O(N__31894),
            .I(N__31797));
    Span4Mux_v I__7517 (
            .O(N__31889),
            .I(N__31797));
    Span4Mux_v I__7516 (
            .O(N__31884),
            .I(N__31797));
    LocalMux I__7515 (
            .O(N__31881),
            .I(N__31788));
    LocalMux I__7514 (
            .O(N__31878),
            .I(N__31788));
    LocalMux I__7513 (
            .O(N__31875),
            .I(N__31788));
    Span4Mux_s3_v I__7512 (
            .O(N__31872),
            .I(N__31788));
    InMux I__7511 (
            .O(N__31869),
            .I(N__31785));
    LocalMux I__7510 (
            .O(N__31866),
            .I(N__31776));
    LocalMux I__7509 (
            .O(N__31863),
            .I(N__31776));
    LocalMux I__7508 (
            .O(N__31860),
            .I(N__31776));
    Span12Mux_s7_v I__7507 (
            .O(N__31853),
            .I(N__31776));
    LocalMux I__7506 (
            .O(N__31850),
            .I(N__31773));
    Span4Mux_v I__7505 (
            .O(N__31837),
            .I(N__31770));
    Span4Mux_h I__7504 (
            .O(N__31834),
            .I(N__31763));
    Span4Mux_v I__7503 (
            .O(N__31829),
            .I(N__31763));
    Span4Mux_v I__7502 (
            .O(N__31820),
            .I(N__31763));
    LocalMux I__7501 (
            .O(N__31817),
            .I(N__31754));
    Span4Mux_h I__7500 (
            .O(N__31814),
            .I(N__31754));
    Span4Mux_h I__7499 (
            .O(N__31807),
            .I(N__31754));
    LocalMux I__7498 (
            .O(N__31804),
            .I(N__31754));
    Span4Mux_h I__7497 (
            .O(N__31797),
            .I(N__31749));
    Span4Mux_v I__7496 (
            .O(N__31788),
            .I(N__31749));
    LocalMux I__7495 (
            .O(N__31785),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__7494 (
            .O(N__31776),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7493 (
            .O(N__31773),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7492 (
            .O(N__31770),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7491 (
            .O(N__31763),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7490 (
            .O(N__31754),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7489 (
            .O(N__31749),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__7488 (
            .O(N__31734),
            .I(N__31726));
    InMux I__7487 (
            .O(N__31733),
            .I(N__31726));
    InMux I__7486 (
            .O(N__31732),
            .I(N__31723));
    InMux I__7485 (
            .O(N__31731),
            .I(N__31719));
    LocalMux I__7484 (
            .O(N__31726),
            .I(N__31716));
    LocalMux I__7483 (
            .O(N__31723),
            .I(N__31713));
    InMux I__7482 (
            .O(N__31722),
            .I(N__31709));
    LocalMux I__7481 (
            .O(N__31719),
            .I(N__31706));
    Span12Mux_s3_h I__7480 (
            .O(N__31716),
            .I(N__31703));
    Span4Mux_h I__7479 (
            .O(N__31713),
            .I(N__31700));
    InMux I__7478 (
            .O(N__31712),
            .I(N__31697));
    LocalMux I__7477 (
            .O(N__31709),
            .I(data_in_field_66));
    Odrv4 I__7476 (
            .O(N__31706),
            .I(data_in_field_66));
    Odrv12 I__7475 (
            .O(N__31703),
            .I(data_in_field_66));
    Odrv4 I__7474 (
            .O(N__31700),
            .I(data_in_field_66));
    LocalMux I__7473 (
            .O(N__31697),
            .I(data_in_field_66));
    CascadeMux I__7472 (
            .O(N__31686),
            .I(N__31682));
    InMux I__7471 (
            .O(N__31685),
            .I(N__31679));
    InMux I__7470 (
            .O(N__31682),
            .I(N__31675));
    LocalMux I__7469 (
            .O(N__31679),
            .I(N__31670));
    InMux I__7468 (
            .O(N__31678),
            .I(N__31667));
    LocalMux I__7467 (
            .O(N__31675),
            .I(N__31664));
    InMux I__7466 (
            .O(N__31674),
            .I(N__31661));
    InMux I__7465 (
            .O(N__31673),
            .I(N__31658));
    Span12Mux_s8_h I__7464 (
            .O(N__31670),
            .I(N__31655));
    LocalMux I__7463 (
            .O(N__31667),
            .I(N__31652));
    Span4Mux_v I__7462 (
            .O(N__31664),
            .I(N__31647));
    LocalMux I__7461 (
            .O(N__31661),
            .I(N__31647));
    LocalMux I__7460 (
            .O(N__31658),
            .I(data_in_field_74));
    Odrv12 I__7459 (
            .O(N__31655),
            .I(data_in_field_74));
    Odrv4 I__7458 (
            .O(N__31652),
            .I(data_in_field_74));
    Odrv4 I__7457 (
            .O(N__31647),
            .I(data_in_field_74));
    InMux I__7456 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__7455 (
            .O(N__31635),
            .I(\c0.n9500 ));
    InMux I__7454 (
            .O(N__31632),
            .I(N__31620));
    InMux I__7453 (
            .O(N__31631),
            .I(N__31620));
    InMux I__7452 (
            .O(N__31630),
            .I(N__31620));
    InMux I__7451 (
            .O(N__31629),
            .I(N__31607));
    InMux I__7450 (
            .O(N__31628),
            .I(N__31607));
    InMux I__7449 (
            .O(N__31627),
            .I(N__31607));
    LocalMux I__7448 (
            .O(N__31620),
            .I(N__31601));
    InMux I__7447 (
            .O(N__31619),
            .I(N__31594));
    InMux I__7446 (
            .O(N__31618),
            .I(N__31594));
    InMux I__7445 (
            .O(N__31617),
            .I(N__31594));
    InMux I__7444 (
            .O(N__31616),
            .I(N__31587));
    InMux I__7443 (
            .O(N__31615),
            .I(N__31587));
    InMux I__7442 (
            .O(N__31614),
            .I(N__31587));
    LocalMux I__7441 (
            .O(N__31607),
            .I(N__31580));
    InMux I__7440 (
            .O(N__31606),
            .I(N__31573));
    InMux I__7439 (
            .O(N__31605),
            .I(N__31573));
    InMux I__7438 (
            .O(N__31604),
            .I(N__31573));
    Span4Mux_s3_v I__7437 (
            .O(N__31601),
            .I(N__31564));
    LocalMux I__7436 (
            .O(N__31594),
            .I(N__31564));
    LocalMux I__7435 (
            .O(N__31587),
            .I(N__31561));
    InMux I__7434 (
            .O(N__31586),
            .I(N__31556));
    InMux I__7433 (
            .O(N__31585),
            .I(N__31556));
    InMux I__7432 (
            .O(N__31584),
            .I(N__31553));
    InMux I__7431 (
            .O(N__31583),
            .I(N__31548));
    Span4Mux_v I__7430 (
            .O(N__31580),
            .I(N__31543));
    LocalMux I__7429 (
            .O(N__31573),
            .I(N__31543));
    InMux I__7428 (
            .O(N__31572),
            .I(N__31536));
    InMux I__7427 (
            .O(N__31571),
            .I(N__31536));
    InMux I__7426 (
            .O(N__31570),
            .I(N__31536));
    InMux I__7425 (
            .O(N__31569),
            .I(N__31533));
    Span4Mux_v I__7424 (
            .O(N__31564),
            .I(N__31529));
    Span4Mux_s3_v I__7423 (
            .O(N__31561),
            .I(N__31526));
    LocalMux I__7422 (
            .O(N__31556),
            .I(N__31521));
    LocalMux I__7421 (
            .O(N__31553),
            .I(N__31521));
    InMux I__7420 (
            .O(N__31552),
            .I(N__31516));
    InMux I__7419 (
            .O(N__31551),
            .I(N__31516));
    LocalMux I__7418 (
            .O(N__31548),
            .I(N__31513));
    Span4Mux_h I__7417 (
            .O(N__31543),
            .I(N__31506));
    LocalMux I__7416 (
            .O(N__31536),
            .I(N__31506));
    LocalMux I__7415 (
            .O(N__31533),
            .I(N__31506));
    InMux I__7414 (
            .O(N__31532),
            .I(N__31503));
    Span4Mux_h I__7413 (
            .O(N__31529),
            .I(N__31498));
    Span4Mux_v I__7412 (
            .O(N__31526),
            .I(N__31498));
    Span12Mux_s7_v I__7411 (
            .O(N__31521),
            .I(N__31493));
    LocalMux I__7410 (
            .O(N__31516),
            .I(N__31493));
    Span4Mux_h I__7409 (
            .O(N__31513),
            .I(N__31488));
    Span4Mux_v I__7408 (
            .O(N__31506),
            .I(N__31488));
    LocalMux I__7407 (
            .O(N__31503),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__7406 (
            .O(N__31498),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__7405 (
            .O(N__31493),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__7404 (
            .O(N__31488),
            .I(\c0.byte_transmit_counter2_3 ));
    CascadeMux I__7403 (
            .O(N__31479),
            .I(\c0.n9198_cascade_ ));
    InMux I__7402 (
            .O(N__31476),
            .I(N__31473));
    LocalMux I__7401 (
            .O(N__31473),
            .I(\c0.n9488 ));
    InMux I__7400 (
            .O(N__31470),
            .I(N__31466));
    InMux I__7399 (
            .O(N__31469),
            .I(N__31463));
    LocalMux I__7398 (
            .O(N__31466),
            .I(N__31457));
    LocalMux I__7397 (
            .O(N__31463),
            .I(N__31454));
    InMux I__7396 (
            .O(N__31462),
            .I(N__31451));
    InMux I__7395 (
            .O(N__31461),
            .I(N__31446));
    InMux I__7394 (
            .O(N__31460),
            .I(N__31446));
    Span12Mux_h I__7393 (
            .O(N__31457),
            .I(N__31443));
    Span4Mux_h I__7392 (
            .O(N__31454),
            .I(N__31436));
    LocalMux I__7391 (
            .O(N__31451),
            .I(N__31436));
    LocalMux I__7390 (
            .O(N__31446),
            .I(N__31436));
    Odrv12 I__7389 (
            .O(N__31443),
            .I(data_in_field_98));
    Odrv4 I__7388 (
            .O(N__31436),
            .I(data_in_field_98));
    InMux I__7387 (
            .O(N__31431),
            .I(N__31428));
    LocalMux I__7386 (
            .O(N__31428),
            .I(N__31425));
    Span4Mux_h I__7385 (
            .O(N__31425),
            .I(N__31422));
    Odrv4 I__7384 (
            .O(N__31422),
            .I(\c0.n9494 ));
    InMux I__7383 (
            .O(N__31419),
            .I(N__31416));
    LocalMux I__7382 (
            .O(N__31416),
            .I(N__31411));
    InMux I__7381 (
            .O(N__31415),
            .I(N__31408));
    InMux I__7380 (
            .O(N__31414),
            .I(N__31404));
    Span12Mux_s4_v I__7379 (
            .O(N__31411),
            .I(N__31399));
    LocalMux I__7378 (
            .O(N__31408),
            .I(N__31399));
    InMux I__7377 (
            .O(N__31407),
            .I(N__31396));
    LocalMux I__7376 (
            .O(N__31404),
            .I(data_in_field_106));
    Odrv12 I__7375 (
            .O(N__31399),
            .I(data_in_field_106));
    LocalMux I__7374 (
            .O(N__31396),
            .I(data_in_field_106));
    InMux I__7373 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__7372 (
            .O(N__31386),
            .I(\c0.n9201 ));
    InMux I__7371 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__7370 (
            .O(N__31380),
            .I(N__31373));
    InMux I__7369 (
            .O(N__31379),
            .I(N__31370));
    InMux I__7368 (
            .O(N__31378),
            .I(N__31367));
    InMux I__7367 (
            .O(N__31377),
            .I(N__31364));
    InMux I__7366 (
            .O(N__31376),
            .I(N__31361));
    Span4Mux_v I__7365 (
            .O(N__31373),
            .I(N__31355));
    LocalMux I__7364 (
            .O(N__31370),
            .I(N__31355));
    LocalMux I__7363 (
            .O(N__31367),
            .I(N__31352));
    LocalMux I__7362 (
            .O(N__31364),
            .I(N__31347));
    LocalMux I__7361 (
            .O(N__31361),
            .I(N__31347));
    InMux I__7360 (
            .O(N__31360),
            .I(N__31344));
    Span4Mux_v I__7359 (
            .O(N__31355),
            .I(N__31340));
    Span4Mux_v I__7358 (
            .O(N__31352),
            .I(N__31337));
    Span4Mux_v I__7357 (
            .O(N__31347),
            .I(N__31334));
    LocalMux I__7356 (
            .O(N__31344),
            .I(N__31331));
    InMux I__7355 (
            .O(N__31343),
            .I(N__31328));
    Span4Mux_s2_v I__7354 (
            .O(N__31340),
            .I(N__31325));
    Span4Mux_v I__7353 (
            .O(N__31337),
            .I(N__31322));
    Span4Mux_v I__7352 (
            .O(N__31334),
            .I(N__31319));
    Span4Mux_h I__7351 (
            .O(N__31331),
            .I(N__31314));
    LocalMux I__7350 (
            .O(N__31328),
            .I(N__31314));
    Span4Mux_h I__7349 (
            .O(N__31325),
            .I(N__31311));
    Span4Mux_s0_v I__7348 (
            .O(N__31322),
            .I(N__31308));
    Span4Mux_h I__7347 (
            .O(N__31319),
            .I(N__31303));
    Span4Mux_v I__7346 (
            .O(N__31314),
            .I(N__31303));
    Odrv4 I__7345 (
            .O(N__31311),
            .I(\c0.n3056 ));
    Odrv4 I__7344 (
            .O(N__31308),
            .I(\c0.n3056 ));
    Odrv4 I__7343 (
            .O(N__31303),
            .I(\c0.n3056 ));
    InMux I__7342 (
            .O(N__31296),
            .I(N__31293));
    LocalMux I__7341 (
            .O(N__31293),
            .I(N__31290));
    Span4Mux_v I__7340 (
            .O(N__31290),
            .I(N__31287));
    Span4Mux_h I__7339 (
            .O(N__31287),
            .I(N__31284));
    Odrv4 I__7338 (
            .O(N__31284),
            .I(\c0.n9671 ));
    CascadeMux I__7337 (
            .O(N__31281),
            .I(N__31278));
    InMux I__7336 (
            .O(N__31278),
            .I(N__31275));
    LocalMux I__7335 (
            .O(N__31275),
            .I(N__31272));
    Span4Mux_h I__7334 (
            .O(N__31272),
            .I(N__31269));
    Span4Mux_h I__7333 (
            .O(N__31269),
            .I(N__31266));
    Odrv4 I__7332 (
            .O(N__31266),
            .I(\c0.data_in_frame_20_6 ));
    InMux I__7331 (
            .O(N__31263),
            .I(N__31260));
    LocalMux I__7330 (
            .O(N__31260),
            .I(N__31256));
    InMux I__7329 (
            .O(N__31259),
            .I(N__31252));
    Span4Mux_s1_v I__7328 (
            .O(N__31256),
            .I(N__31249));
    InMux I__7327 (
            .O(N__31255),
            .I(N__31246));
    LocalMux I__7326 (
            .O(N__31252),
            .I(N__31239));
    Span4Mux_h I__7325 (
            .O(N__31249),
            .I(N__31234));
    LocalMux I__7324 (
            .O(N__31246),
            .I(N__31234));
    InMux I__7323 (
            .O(N__31245),
            .I(N__31226));
    InMux I__7322 (
            .O(N__31244),
            .I(N__31223));
    InMux I__7321 (
            .O(N__31243),
            .I(N__31220));
    InMux I__7320 (
            .O(N__31242),
            .I(N__31217));
    Span4Mux_v I__7319 (
            .O(N__31239),
            .I(N__31214));
    Span4Mux_v I__7318 (
            .O(N__31234),
            .I(N__31211));
    InMux I__7317 (
            .O(N__31233),
            .I(N__31208));
    InMux I__7316 (
            .O(N__31232),
            .I(N__31205));
    InMux I__7315 (
            .O(N__31231),
            .I(N__31200));
    InMux I__7314 (
            .O(N__31230),
            .I(N__31197));
    InMux I__7313 (
            .O(N__31229),
            .I(N__31194));
    LocalMux I__7312 (
            .O(N__31226),
            .I(N__31189));
    LocalMux I__7311 (
            .O(N__31223),
            .I(N__31186));
    LocalMux I__7310 (
            .O(N__31220),
            .I(N__31183));
    LocalMux I__7309 (
            .O(N__31217),
            .I(N__31180));
    Sp12to4 I__7308 (
            .O(N__31214),
            .I(N__31169));
    Sp12to4 I__7307 (
            .O(N__31211),
            .I(N__31169));
    LocalMux I__7306 (
            .O(N__31208),
            .I(N__31169));
    LocalMux I__7305 (
            .O(N__31205),
            .I(N__31169));
    InMux I__7304 (
            .O(N__31204),
            .I(N__31166));
    InMux I__7303 (
            .O(N__31203),
            .I(N__31163));
    LocalMux I__7302 (
            .O(N__31200),
            .I(N__31156));
    LocalMux I__7301 (
            .O(N__31197),
            .I(N__31156));
    LocalMux I__7300 (
            .O(N__31194),
            .I(N__31156));
    InMux I__7299 (
            .O(N__31193),
            .I(N__31153));
    InMux I__7298 (
            .O(N__31192),
            .I(N__31150));
    Span4Mux_h I__7297 (
            .O(N__31189),
            .I(N__31141));
    Span4Mux_h I__7296 (
            .O(N__31186),
            .I(N__31141));
    Span4Mux_s1_v I__7295 (
            .O(N__31183),
            .I(N__31141));
    Span4Mux_h I__7294 (
            .O(N__31180),
            .I(N__31141));
    InMux I__7293 (
            .O(N__31179),
            .I(N__31138));
    InMux I__7292 (
            .O(N__31178),
            .I(N__31135));
    Span12Mux_h I__7291 (
            .O(N__31169),
            .I(N__31132));
    LocalMux I__7290 (
            .O(N__31166),
            .I(N__31123));
    LocalMux I__7289 (
            .O(N__31163),
            .I(N__31123));
    Span12Mux_s7_v I__7288 (
            .O(N__31156),
            .I(N__31123));
    LocalMux I__7287 (
            .O(N__31153),
            .I(N__31123));
    LocalMux I__7286 (
            .O(N__31150),
            .I(N__31116));
    Sp12to4 I__7285 (
            .O(N__31141),
            .I(N__31116));
    LocalMux I__7284 (
            .O(N__31138),
            .I(N__31116));
    LocalMux I__7283 (
            .O(N__31135),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv12 I__7282 (
            .O(N__31132),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv12 I__7281 (
            .O(N__31123),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv12 I__7280 (
            .O(N__31116),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__7279 (
            .O(N__31107),
            .I(N__31104));
    LocalMux I__7278 (
            .O(N__31104),
            .I(N__31101));
    Span4Mux_s1_v I__7277 (
            .O(N__31101),
            .I(N__31098));
    Span4Mux_h I__7276 (
            .O(N__31098),
            .I(N__31095));
    Odrv4 I__7275 (
            .O(N__31095),
            .I(\c0.n22_adj_1677 ));
    InMux I__7274 (
            .O(N__31092),
            .I(\c0.rx.n8101 ));
    InMux I__7273 (
            .O(N__31089),
            .I(\c0.rx.n8102 ));
    InMux I__7272 (
            .O(N__31086),
            .I(N__31083));
    LocalMux I__7271 (
            .O(N__31083),
            .I(N__31080));
    Span4Mux_h I__7270 (
            .O(N__31080),
            .I(N__31077));
    Span4Mux_h I__7269 (
            .O(N__31077),
            .I(N__31069));
    InMux I__7268 (
            .O(N__31076),
            .I(N__31066));
    InMux I__7267 (
            .O(N__31075),
            .I(N__31063));
    InMux I__7266 (
            .O(N__31074),
            .I(N__31058));
    InMux I__7265 (
            .O(N__31073),
            .I(N__31058));
    InMux I__7264 (
            .O(N__31072),
            .I(N__31055));
    Odrv4 I__7263 (
            .O(N__31069),
            .I(r_Clock_Count_6_adj_1728));
    LocalMux I__7262 (
            .O(N__31066),
            .I(r_Clock_Count_6_adj_1728));
    LocalMux I__7261 (
            .O(N__31063),
            .I(r_Clock_Count_6_adj_1728));
    LocalMux I__7260 (
            .O(N__31058),
            .I(r_Clock_Count_6_adj_1728));
    LocalMux I__7259 (
            .O(N__31055),
            .I(r_Clock_Count_6_adj_1728));
    CascadeMux I__7258 (
            .O(N__31044),
            .I(N__31041));
    InMux I__7257 (
            .O(N__31041),
            .I(N__31038));
    LocalMux I__7256 (
            .O(N__31038),
            .I(n220));
    InMux I__7255 (
            .O(N__31035),
            .I(\c0.rx.n8103 ));
    CascadeMux I__7254 (
            .O(N__31032),
            .I(N__31029));
    InMux I__7253 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__7252 (
            .O(N__31026),
            .I(N__31023));
    Span4Mux_h I__7251 (
            .O(N__31023),
            .I(N__31017));
    CascadeMux I__7250 (
            .O(N__31022),
            .I(N__31013));
    CascadeMux I__7249 (
            .O(N__31021),
            .I(N__31009));
    InMux I__7248 (
            .O(N__31020),
            .I(N__31006));
    Span4Mux_v I__7247 (
            .O(N__31017),
            .I(N__31003));
    InMux I__7246 (
            .O(N__31016),
            .I(N__31000));
    InMux I__7245 (
            .O(N__31013),
            .I(N__30997));
    InMux I__7244 (
            .O(N__31012),
            .I(N__30992));
    InMux I__7243 (
            .O(N__31009),
            .I(N__30992));
    LocalMux I__7242 (
            .O(N__31006),
            .I(r_Clock_Count_7_adj_1727));
    Odrv4 I__7241 (
            .O(N__31003),
            .I(r_Clock_Count_7_adj_1727));
    LocalMux I__7240 (
            .O(N__31000),
            .I(r_Clock_Count_7_adj_1727));
    LocalMux I__7239 (
            .O(N__30997),
            .I(r_Clock_Count_7_adj_1727));
    LocalMux I__7238 (
            .O(N__30992),
            .I(r_Clock_Count_7_adj_1727));
    InMux I__7237 (
            .O(N__30981),
            .I(\c0.rx.n8104 ));
    InMux I__7236 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__7235 (
            .O(N__30975),
            .I(n219));
    InMux I__7234 (
            .O(N__30972),
            .I(N__30969));
    LocalMux I__7233 (
            .O(N__30969),
            .I(N__30966));
    Span4Mux_v I__7232 (
            .O(N__30966),
            .I(N__30960));
    InMux I__7231 (
            .O(N__30965),
            .I(N__30955));
    InMux I__7230 (
            .O(N__30964),
            .I(N__30955));
    InMux I__7229 (
            .O(N__30963),
            .I(N__30952));
    Span4Mux_h I__7228 (
            .O(N__30960),
            .I(N__30947));
    LocalMux I__7227 (
            .O(N__30955),
            .I(N__30947));
    LocalMux I__7226 (
            .O(N__30952),
            .I(n4084));
    Odrv4 I__7225 (
            .O(N__30947),
            .I(n4084));
    CascadeMux I__7224 (
            .O(N__30942),
            .I(N__30939));
    InMux I__7223 (
            .O(N__30939),
            .I(N__30936));
    LocalMux I__7222 (
            .O(N__30936),
            .I(N__30933));
    Odrv4 I__7221 (
            .O(N__30933),
            .I(n221));
    InMux I__7220 (
            .O(N__30930),
            .I(N__30925));
    InMux I__7219 (
            .O(N__30929),
            .I(N__30920));
    InMux I__7218 (
            .O(N__30928),
            .I(N__30920));
    LocalMux I__7217 (
            .O(N__30925),
            .I(r_Clock_Count_5));
    LocalMux I__7216 (
            .O(N__30920),
            .I(r_Clock_Count_5));
    InMux I__7215 (
            .O(N__30915),
            .I(N__30904));
    InMux I__7214 (
            .O(N__30914),
            .I(N__30904));
    InMux I__7213 (
            .O(N__30913),
            .I(N__30895));
    InMux I__7212 (
            .O(N__30912),
            .I(N__30895));
    InMux I__7211 (
            .O(N__30911),
            .I(N__30895));
    InMux I__7210 (
            .O(N__30910),
            .I(N__30895));
    InMux I__7209 (
            .O(N__30909),
            .I(N__30892));
    LocalMux I__7208 (
            .O(N__30904),
            .I(n30));
    LocalMux I__7207 (
            .O(N__30895),
            .I(n30));
    LocalMux I__7206 (
            .O(N__30892),
            .I(n30));
    CascadeMux I__7205 (
            .O(N__30885),
            .I(N__30882));
    InMux I__7204 (
            .O(N__30882),
            .I(N__30879));
    LocalMux I__7203 (
            .O(N__30879),
            .I(n222));
    CascadeMux I__7202 (
            .O(N__30876),
            .I(N__30870));
    InMux I__7201 (
            .O(N__30875),
            .I(N__30862));
    InMux I__7200 (
            .O(N__30874),
            .I(N__30862));
    InMux I__7199 (
            .O(N__30873),
            .I(N__30859));
    InMux I__7198 (
            .O(N__30870),
            .I(N__30856));
    InMux I__7197 (
            .O(N__30869),
            .I(N__30849));
    InMux I__7196 (
            .O(N__30868),
            .I(N__30849));
    InMux I__7195 (
            .O(N__30867),
            .I(N__30849));
    LocalMux I__7194 (
            .O(N__30862),
            .I(N__30846));
    LocalMux I__7193 (
            .O(N__30859),
            .I(n44));
    LocalMux I__7192 (
            .O(N__30856),
            .I(n44));
    LocalMux I__7191 (
            .O(N__30849),
            .I(n44));
    Odrv4 I__7190 (
            .O(N__30846),
            .I(n44));
    InMux I__7189 (
            .O(N__30837),
            .I(N__30832));
    InMux I__7188 (
            .O(N__30836),
            .I(N__30827));
    InMux I__7187 (
            .O(N__30835),
            .I(N__30827));
    LocalMux I__7186 (
            .O(N__30832),
            .I(r_Clock_Count_4_adj_1729));
    LocalMux I__7185 (
            .O(N__30827),
            .I(r_Clock_Count_4_adj_1729));
    InMux I__7184 (
            .O(N__30822),
            .I(N__30819));
    LocalMux I__7183 (
            .O(N__30819),
            .I(N__30816));
    Span4Mux_v I__7182 (
            .O(N__30816),
            .I(N__30813));
    Sp12to4 I__7181 (
            .O(N__30813),
            .I(N__30810));
    Odrv12 I__7180 (
            .O(N__30810),
            .I(\c0.n9192 ));
    CascadeMux I__7179 (
            .O(N__30807),
            .I(N__30804));
    InMux I__7178 (
            .O(N__30804),
            .I(N__30801));
    LocalMux I__7177 (
            .O(N__30801),
            .I(N__30798));
    Span12Mux_h I__7176 (
            .O(N__30798),
            .I(N__30795));
    Odrv12 I__7175 (
            .O(N__30795),
            .I(\c0.n9195 ));
    InMux I__7174 (
            .O(N__30792),
            .I(N__30778));
    InMux I__7173 (
            .O(N__30791),
            .I(N__30778));
    InMux I__7172 (
            .O(N__30790),
            .I(N__30771));
    InMux I__7171 (
            .O(N__30789),
            .I(N__30771));
    InMux I__7170 (
            .O(N__30788),
            .I(N__30771));
    InMux I__7169 (
            .O(N__30787),
            .I(N__30768));
    InMux I__7168 (
            .O(N__30786),
            .I(N__30765));
    InMux I__7167 (
            .O(N__30785),
            .I(N__30760));
    InMux I__7166 (
            .O(N__30784),
            .I(N__30760));
    InMux I__7165 (
            .O(N__30783),
            .I(N__30757));
    LocalMux I__7164 (
            .O(N__30778),
            .I(N__30752));
    LocalMux I__7163 (
            .O(N__30771),
            .I(N__30752));
    LocalMux I__7162 (
            .O(N__30768),
            .I(N__30747));
    LocalMux I__7161 (
            .O(N__30765),
            .I(N__30747));
    LocalMux I__7160 (
            .O(N__30760),
            .I(r_SM_Main_1_adj_1735));
    LocalMux I__7159 (
            .O(N__30757),
            .I(r_SM_Main_1_adj_1735));
    Odrv12 I__7158 (
            .O(N__30752),
            .I(r_SM_Main_1_adj_1735));
    Odrv4 I__7157 (
            .O(N__30747),
            .I(r_SM_Main_1_adj_1735));
    InMux I__7156 (
            .O(N__30738),
            .I(N__30735));
    LocalMux I__7155 (
            .O(N__30735),
            .I(n9246));
    CascadeMux I__7154 (
            .O(N__30732),
            .I(N__30729));
    InMux I__7153 (
            .O(N__30729),
            .I(N__30725));
    CascadeMux I__7152 (
            .O(N__30728),
            .I(N__30716));
    LocalMux I__7151 (
            .O(N__30725),
            .I(N__30711));
    InMux I__7150 (
            .O(N__30724),
            .I(N__30708));
    InMux I__7149 (
            .O(N__30723),
            .I(N__30703));
    InMux I__7148 (
            .O(N__30722),
            .I(N__30703));
    InMux I__7147 (
            .O(N__30721),
            .I(N__30700));
    InMux I__7146 (
            .O(N__30720),
            .I(N__30697));
    InMux I__7145 (
            .O(N__30719),
            .I(N__30690));
    InMux I__7144 (
            .O(N__30716),
            .I(N__30690));
    InMux I__7143 (
            .O(N__30715),
            .I(N__30690));
    InMux I__7142 (
            .O(N__30714),
            .I(N__30687));
    Span4Mux_v I__7141 (
            .O(N__30711),
            .I(N__30684));
    LocalMux I__7140 (
            .O(N__30708),
            .I(N__30679));
    LocalMux I__7139 (
            .O(N__30703),
            .I(N__30679));
    LocalMux I__7138 (
            .O(N__30700),
            .I(N__30676));
    LocalMux I__7137 (
            .O(N__30697),
            .I(r_SM_Main_0_adj_1736));
    LocalMux I__7136 (
            .O(N__30690),
            .I(r_SM_Main_0_adj_1736));
    LocalMux I__7135 (
            .O(N__30687),
            .I(r_SM_Main_0_adj_1736));
    Odrv4 I__7134 (
            .O(N__30684),
            .I(r_SM_Main_0_adj_1736));
    Odrv12 I__7133 (
            .O(N__30679),
            .I(r_SM_Main_0_adj_1736));
    Odrv4 I__7132 (
            .O(N__30676),
            .I(r_SM_Main_0_adj_1736));
    CascadeMux I__7131 (
            .O(N__30663),
            .I(n44_cascade_));
    InMux I__7130 (
            .O(N__30660),
            .I(N__30652));
    InMux I__7129 (
            .O(N__30659),
            .I(N__30652));
    InMux I__7128 (
            .O(N__30658),
            .I(N__30649));
    CascadeMux I__7127 (
            .O(N__30657),
            .I(N__30643));
    LocalMux I__7126 (
            .O(N__30652),
            .I(N__30636));
    LocalMux I__7125 (
            .O(N__30649),
            .I(N__30636));
    InMux I__7124 (
            .O(N__30648),
            .I(N__30629));
    InMux I__7123 (
            .O(N__30647),
            .I(N__30629));
    InMux I__7122 (
            .O(N__30646),
            .I(N__30629));
    InMux I__7121 (
            .O(N__30643),
            .I(N__30626));
    InMux I__7120 (
            .O(N__30642),
            .I(N__30623));
    InMux I__7119 (
            .O(N__30641),
            .I(N__30620));
    Span4Mux_s2_v I__7118 (
            .O(N__30636),
            .I(N__30617));
    LocalMux I__7117 (
            .O(N__30629),
            .I(N__30614));
    LocalMux I__7116 (
            .O(N__30626),
            .I(N__30611));
    LocalMux I__7115 (
            .O(N__30623),
            .I(N__30608));
    LocalMux I__7114 (
            .O(N__30620),
            .I(N__30605));
    Span4Mux_v I__7113 (
            .O(N__30617),
            .I(N__30602));
    Span4Mux_s2_v I__7112 (
            .O(N__30614),
            .I(N__30599));
    Span4Mux_s2_v I__7111 (
            .O(N__30611),
            .I(N__30592));
    Span4Mux_h I__7110 (
            .O(N__30608),
            .I(N__30592));
    Span4Mux_h I__7109 (
            .O(N__30605),
            .I(N__30592));
    Span4Mux_h I__7108 (
            .O(N__30602),
            .I(N__30589));
    Span4Mux_v I__7107 (
            .O(N__30599),
            .I(N__30584));
    Span4Mux_v I__7106 (
            .O(N__30592),
            .I(N__30584));
    Odrv4 I__7105 (
            .O(N__30589),
            .I(r_SM_Main_2_adj_1734));
    Odrv4 I__7104 (
            .O(N__30584),
            .I(r_SM_Main_2_adj_1734));
    CascadeMux I__7103 (
            .O(N__30579),
            .I(N__30576));
    InMux I__7102 (
            .O(N__30576),
            .I(N__30573));
    LocalMux I__7101 (
            .O(N__30573),
            .I(N__30570));
    Span4Mux_s2_v I__7100 (
            .O(N__30570),
            .I(N__30564));
    InMux I__7099 (
            .O(N__30569),
            .I(N__30558));
    InMux I__7098 (
            .O(N__30568),
            .I(N__30558));
    InMux I__7097 (
            .O(N__30567),
            .I(N__30555));
    Span4Mux_h I__7096 (
            .O(N__30564),
            .I(N__30552));
    InMux I__7095 (
            .O(N__30563),
            .I(N__30549));
    LocalMux I__7094 (
            .O(N__30558),
            .I(N__30544));
    LocalMux I__7093 (
            .O(N__30555),
            .I(N__30544));
    Odrv4 I__7092 (
            .O(N__30552),
            .I(r_SM_Main_2_N_1537_2));
    LocalMux I__7091 (
            .O(N__30549),
            .I(r_SM_Main_2_N_1537_2));
    Odrv4 I__7090 (
            .O(N__30544),
            .I(r_SM_Main_2_N_1537_2));
    InMux I__7089 (
            .O(N__30537),
            .I(N__30534));
    LocalMux I__7088 (
            .O(N__30534),
            .I(n9245));
    CascadeMux I__7087 (
            .O(N__30531),
            .I(N__30527));
    CascadeMux I__7086 (
            .O(N__30530),
            .I(N__30524));
    InMux I__7085 (
            .O(N__30527),
            .I(N__30519));
    InMux I__7084 (
            .O(N__30524),
            .I(N__30516));
    InMux I__7083 (
            .O(N__30523),
            .I(N__30511));
    InMux I__7082 (
            .O(N__30522),
            .I(N__30511));
    LocalMux I__7081 (
            .O(N__30519),
            .I(r_Clock_Count_0_adj_1730));
    LocalMux I__7080 (
            .O(N__30516),
            .I(r_Clock_Count_0_adj_1730));
    LocalMux I__7079 (
            .O(N__30511),
            .I(r_Clock_Count_0_adj_1730));
    InMux I__7078 (
            .O(N__30504),
            .I(N__30501));
    LocalMux I__7077 (
            .O(N__30501),
            .I(n226));
    InMux I__7076 (
            .O(N__30498),
            .I(bfn_11_31_0_));
    CascadeMux I__7075 (
            .O(N__30495),
            .I(N__30492));
    InMux I__7074 (
            .O(N__30492),
            .I(N__30485));
    InMux I__7073 (
            .O(N__30491),
            .I(N__30482));
    InMux I__7072 (
            .O(N__30490),
            .I(N__30479));
    InMux I__7071 (
            .O(N__30489),
            .I(N__30474));
    InMux I__7070 (
            .O(N__30488),
            .I(N__30474));
    LocalMux I__7069 (
            .O(N__30485),
            .I(r_Clock_Count_1));
    LocalMux I__7068 (
            .O(N__30482),
            .I(r_Clock_Count_1));
    LocalMux I__7067 (
            .O(N__30479),
            .I(r_Clock_Count_1));
    LocalMux I__7066 (
            .O(N__30474),
            .I(r_Clock_Count_1));
    InMux I__7065 (
            .O(N__30465),
            .I(N__30462));
    LocalMux I__7064 (
            .O(N__30462),
            .I(N__30459));
    Odrv4 I__7063 (
            .O(N__30459),
            .I(n225));
    InMux I__7062 (
            .O(N__30456),
            .I(\c0.rx.n8098 ));
    InMux I__7061 (
            .O(N__30453),
            .I(N__30446));
    InMux I__7060 (
            .O(N__30452),
            .I(N__30443));
    InMux I__7059 (
            .O(N__30451),
            .I(N__30440));
    InMux I__7058 (
            .O(N__30450),
            .I(N__30435));
    InMux I__7057 (
            .O(N__30449),
            .I(N__30435));
    LocalMux I__7056 (
            .O(N__30446),
            .I(r_Clock_Count_2));
    LocalMux I__7055 (
            .O(N__30443),
            .I(r_Clock_Count_2));
    LocalMux I__7054 (
            .O(N__30440),
            .I(r_Clock_Count_2));
    LocalMux I__7053 (
            .O(N__30435),
            .I(r_Clock_Count_2));
    CascadeMux I__7052 (
            .O(N__30426),
            .I(N__30423));
    InMux I__7051 (
            .O(N__30423),
            .I(N__30420));
    LocalMux I__7050 (
            .O(N__30420),
            .I(n224));
    InMux I__7049 (
            .O(N__30417),
            .I(\c0.rx.n8099 ));
    InMux I__7048 (
            .O(N__30414),
            .I(N__30407));
    InMux I__7047 (
            .O(N__30413),
            .I(N__30404));
    InMux I__7046 (
            .O(N__30412),
            .I(N__30401));
    InMux I__7045 (
            .O(N__30411),
            .I(N__30396));
    InMux I__7044 (
            .O(N__30410),
            .I(N__30396));
    LocalMux I__7043 (
            .O(N__30407),
            .I(r_Clock_Count_3));
    LocalMux I__7042 (
            .O(N__30404),
            .I(r_Clock_Count_3));
    LocalMux I__7041 (
            .O(N__30401),
            .I(r_Clock_Count_3));
    LocalMux I__7040 (
            .O(N__30396),
            .I(r_Clock_Count_3));
    InMux I__7039 (
            .O(N__30387),
            .I(N__30384));
    LocalMux I__7038 (
            .O(N__30384),
            .I(n223));
    InMux I__7037 (
            .O(N__30381),
            .I(\c0.rx.n8100 ));
    InMux I__7036 (
            .O(N__30378),
            .I(N__30375));
    LocalMux I__7035 (
            .O(N__30375),
            .I(n7));
    InMux I__7034 (
            .O(N__30372),
            .I(n8148));
    InMux I__7033 (
            .O(N__30369),
            .I(N__30366));
    LocalMux I__7032 (
            .O(N__30366),
            .I(n6));
    InMux I__7031 (
            .O(N__30363),
            .I(n8149));
    CascadeMux I__7030 (
            .O(N__30360),
            .I(N__30356));
    InMux I__7029 (
            .O(N__30359),
            .I(N__30351));
    InMux I__7028 (
            .O(N__30356),
            .I(N__30351));
    LocalMux I__7027 (
            .O(N__30351),
            .I(N__30348));
    Span4Mux_h I__7026 (
            .O(N__30348),
            .I(N__30345));
    Sp12to4 I__7025 (
            .O(N__30345),
            .I(N__30342));
    Span12Mux_v I__7024 (
            .O(N__30342),
            .I(N__30338));
    InMux I__7023 (
            .O(N__30341),
            .I(N__30335));
    Odrv12 I__7022 (
            .O(N__30338),
            .I(blink_counter_21));
    LocalMux I__7021 (
            .O(N__30335),
            .I(blink_counter_21));
    InMux I__7020 (
            .O(N__30330),
            .I(n8150));
    CascadeMux I__7019 (
            .O(N__30327),
            .I(N__30324));
    InMux I__7018 (
            .O(N__30324),
            .I(N__30318));
    InMux I__7017 (
            .O(N__30323),
            .I(N__30318));
    LocalMux I__7016 (
            .O(N__30318),
            .I(N__30315));
    Span4Mux_v I__7015 (
            .O(N__30315),
            .I(N__30312));
    Span4Mux_h I__7014 (
            .O(N__30312),
            .I(N__30308));
    InMux I__7013 (
            .O(N__30311),
            .I(N__30305));
    Odrv4 I__7012 (
            .O(N__30308),
            .I(blink_counter_22));
    LocalMux I__7011 (
            .O(N__30305),
            .I(blink_counter_22));
    InMux I__7010 (
            .O(N__30300),
            .I(n8151));
    InMux I__7009 (
            .O(N__30297),
            .I(N__30291));
    InMux I__7008 (
            .O(N__30296),
            .I(N__30291));
    LocalMux I__7007 (
            .O(N__30291),
            .I(N__30288));
    Span4Mux_h I__7006 (
            .O(N__30288),
            .I(N__30285));
    Span4Mux_h I__7005 (
            .O(N__30285),
            .I(N__30281));
    InMux I__7004 (
            .O(N__30284),
            .I(N__30278));
    Odrv4 I__7003 (
            .O(N__30281),
            .I(blink_counter_23));
    LocalMux I__7002 (
            .O(N__30278),
            .I(blink_counter_23));
    InMux I__7001 (
            .O(N__30273),
            .I(n8152));
    InMux I__7000 (
            .O(N__30270),
            .I(N__30264));
    InMux I__6999 (
            .O(N__30269),
            .I(N__30264));
    LocalMux I__6998 (
            .O(N__30264),
            .I(N__30261));
    Span12Mux_s10_h I__6997 (
            .O(N__30261),
            .I(N__30257));
    InMux I__6996 (
            .O(N__30260),
            .I(N__30254));
    Odrv12 I__6995 (
            .O(N__30257),
            .I(blink_counter_24));
    LocalMux I__6994 (
            .O(N__30254),
            .I(blink_counter_24));
    InMux I__6993 (
            .O(N__30249),
            .I(bfn_11_30_0_));
    InMux I__6992 (
            .O(N__30246),
            .I(n8154));
    InMux I__6991 (
            .O(N__30243),
            .I(N__30240));
    LocalMux I__6990 (
            .O(N__30240),
            .I(N__30237));
    Span12Mux_v I__6989 (
            .O(N__30237),
            .I(N__30233));
    InMux I__6988 (
            .O(N__30236),
            .I(N__30230));
    Odrv12 I__6987 (
            .O(N__30233),
            .I(blink_counter_25));
    LocalMux I__6986 (
            .O(N__30230),
            .I(blink_counter_25));
    InMux I__6985 (
            .O(N__30225),
            .I(N__30222));
    LocalMux I__6984 (
            .O(N__30222),
            .I(n15));
    InMux I__6983 (
            .O(N__30219),
            .I(n8140));
    InMux I__6982 (
            .O(N__30216),
            .I(N__30213));
    LocalMux I__6981 (
            .O(N__30213),
            .I(n14));
    InMux I__6980 (
            .O(N__30210),
            .I(n8141));
    InMux I__6979 (
            .O(N__30207),
            .I(N__30204));
    LocalMux I__6978 (
            .O(N__30204),
            .I(n13));
    InMux I__6977 (
            .O(N__30201),
            .I(n8142));
    InMux I__6976 (
            .O(N__30198),
            .I(N__30195));
    LocalMux I__6975 (
            .O(N__30195),
            .I(n12));
    InMux I__6974 (
            .O(N__30192),
            .I(n8143));
    InMux I__6973 (
            .O(N__30189),
            .I(N__30186));
    LocalMux I__6972 (
            .O(N__30186),
            .I(n11));
    InMux I__6971 (
            .O(N__30183),
            .I(n8144));
    InMux I__6970 (
            .O(N__30180),
            .I(N__30177));
    LocalMux I__6969 (
            .O(N__30177),
            .I(n10));
    InMux I__6968 (
            .O(N__30174),
            .I(bfn_11_29_0_));
    InMux I__6967 (
            .O(N__30171),
            .I(N__30168));
    LocalMux I__6966 (
            .O(N__30168),
            .I(n9));
    InMux I__6965 (
            .O(N__30165),
            .I(n8146));
    InMux I__6964 (
            .O(N__30162),
            .I(N__30159));
    LocalMux I__6963 (
            .O(N__30159),
            .I(n8));
    InMux I__6962 (
            .O(N__30156),
            .I(n8147));
    InMux I__6961 (
            .O(N__30153),
            .I(N__30150));
    LocalMux I__6960 (
            .O(N__30150),
            .I(n24));
    InMux I__6959 (
            .O(N__30147),
            .I(n8131));
    InMux I__6958 (
            .O(N__30144),
            .I(N__30141));
    LocalMux I__6957 (
            .O(N__30141),
            .I(n23));
    InMux I__6956 (
            .O(N__30138),
            .I(n8132));
    InMux I__6955 (
            .O(N__30135),
            .I(N__30132));
    LocalMux I__6954 (
            .O(N__30132),
            .I(n22));
    InMux I__6953 (
            .O(N__30129),
            .I(n8133));
    InMux I__6952 (
            .O(N__30126),
            .I(N__30123));
    LocalMux I__6951 (
            .O(N__30123),
            .I(n21));
    InMux I__6950 (
            .O(N__30120),
            .I(n8134));
    InMux I__6949 (
            .O(N__30117),
            .I(N__30114));
    LocalMux I__6948 (
            .O(N__30114),
            .I(n20));
    InMux I__6947 (
            .O(N__30111),
            .I(n8135));
    InMux I__6946 (
            .O(N__30108),
            .I(N__30105));
    LocalMux I__6945 (
            .O(N__30105),
            .I(n19));
    InMux I__6944 (
            .O(N__30102),
            .I(n8136));
    InMux I__6943 (
            .O(N__30099),
            .I(N__30096));
    LocalMux I__6942 (
            .O(N__30096),
            .I(n18));
    InMux I__6941 (
            .O(N__30093),
            .I(bfn_11_28_0_));
    InMux I__6940 (
            .O(N__30090),
            .I(N__30087));
    LocalMux I__6939 (
            .O(N__30087),
            .I(n17));
    InMux I__6938 (
            .O(N__30084),
            .I(n8138));
    InMux I__6937 (
            .O(N__30081),
            .I(N__30078));
    LocalMux I__6936 (
            .O(N__30078),
            .I(n16));
    InMux I__6935 (
            .O(N__30075),
            .I(n8139));
    CascadeMux I__6934 (
            .O(N__30072),
            .I(N__30069));
    InMux I__6933 (
            .O(N__30069),
            .I(N__30066));
    LocalMux I__6932 (
            .O(N__30066),
            .I(N__30063));
    Odrv4 I__6931 (
            .O(N__30063),
            .I(\c0.n22_adj_1661 ));
    InMux I__6930 (
            .O(N__30060),
            .I(N__30057));
    LocalMux I__6929 (
            .O(N__30057),
            .I(\c0.n9731 ));
    InMux I__6928 (
            .O(N__30054),
            .I(N__30051));
    LocalMux I__6927 (
            .O(N__30051),
            .I(N__30048));
    Span4Mux_h I__6926 (
            .O(N__30048),
            .I(N__30045));
    Span4Mux_h I__6925 (
            .O(N__30045),
            .I(N__30042));
    Span4Mux_v I__6924 (
            .O(N__30042),
            .I(N__30039));
    Odrv4 I__6923 (
            .O(N__30039),
            .I(\c0.tx2.r_Tx_Data_0 ));
    CascadeMux I__6922 (
            .O(N__30036),
            .I(N__30025));
    CascadeMux I__6921 (
            .O(N__30035),
            .I(N__30015));
    CascadeMux I__6920 (
            .O(N__30034),
            .I(N__30012));
    CascadeMux I__6919 (
            .O(N__30033),
            .I(N__30009));
    InMux I__6918 (
            .O(N__30032),
            .I(N__30002));
    CascadeMux I__6917 (
            .O(N__30031),
            .I(N__29999));
    CascadeMux I__6916 (
            .O(N__30030),
            .I(N__29996));
    CascadeMux I__6915 (
            .O(N__30029),
            .I(N__29961));
    CascadeMux I__6914 (
            .O(N__30028),
            .I(N__29958));
    InMux I__6913 (
            .O(N__30025),
            .I(N__29942));
    InMux I__6912 (
            .O(N__30024),
            .I(N__29942));
    InMux I__6911 (
            .O(N__30023),
            .I(N__29942));
    InMux I__6910 (
            .O(N__30022),
            .I(N__29942));
    InMux I__6909 (
            .O(N__30021),
            .I(N__29942));
    CascadeMux I__6908 (
            .O(N__30020),
            .I(N__29939));
    CascadeMux I__6907 (
            .O(N__30019),
            .I(N__29936));
    CascadeMux I__6906 (
            .O(N__30018),
            .I(N__29933));
    InMux I__6905 (
            .O(N__30015),
            .I(N__29908));
    InMux I__6904 (
            .O(N__30012),
            .I(N__29908));
    InMux I__6903 (
            .O(N__30009),
            .I(N__29908));
    InMux I__6902 (
            .O(N__30008),
            .I(N__29908));
    InMux I__6901 (
            .O(N__30007),
            .I(N__29908));
    InMux I__6900 (
            .O(N__30006),
            .I(N__29908));
    InMux I__6899 (
            .O(N__30005),
            .I(N__29908));
    LocalMux I__6898 (
            .O(N__30002),
            .I(N__29905));
    InMux I__6897 (
            .O(N__29999),
            .I(N__29894));
    InMux I__6896 (
            .O(N__29996),
            .I(N__29894));
    InMux I__6895 (
            .O(N__29995),
            .I(N__29894));
    InMux I__6894 (
            .O(N__29994),
            .I(N__29894));
    InMux I__6893 (
            .O(N__29993),
            .I(N__29894));
    InMux I__6892 (
            .O(N__29992),
            .I(N__29887));
    InMux I__6891 (
            .O(N__29991),
            .I(N__29887));
    InMux I__6890 (
            .O(N__29990),
            .I(N__29887));
    CascadeMux I__6889 (
            .O(N__29989),
            .I(N__29879));
    CascadeMux I__6888 (
            .O(N__29988),
            .I(N__29876));
    CascadeMux I__6887 (
            .O(N__29987),
            .I(N__29867));
    CascadeMux I__6886 (
            .O(N__29986),
            .I(N__29863));
    InMux I__6885 (
            .O(N__29985),
            .I(N__29846));
    InMux I__6884 (
            .O(N__29984),
            .I(N__29846));
    InMux I__6883 (
            .O(N__29983),
            .I(N__29846));
    InMux I__6882 (
            .O(N__29982),
            .I(N__29846));
    InMux I__6881 (
            .O(N__29981),
            .I(N__29846));
    InMux I__6880 (
            .O(N__29980),
            .I(N__29846));
    InMux I__6879 (
            .O(N__29979),
            .I(N__29830));
    InMux I__6878 (
            .O(N__29978),
            .I(N__29830));
    InMux I__6877 (
            .O(N__29977),
            .I(N__29830));
    InMux I__6876 (
            .O(N__29976),
            .I(N__29825));
    InMux I__6875 (
            .O(N__29975),
            .I(N__29825));
    InMux I__6874 (
            .O(N__29974),
            .I(N__29816));
    InMux I__6873 (
            .O(N__29973),
            .I(N__29816));
    InMux I__6872 (
            .O(N__29972),
            .I(N__29816));
    InMux I__6871 (
            .O(N__29971),
            .I(N__29816));
    InMux I__6870 (
            .O(N__29970),
            .I(N__29805));
    InMux I__6869 (
            .O(N__29969),
            .I(N__29805));
    InMux I__6868 (
            .O(N__29968),
            .I(N__29805));
    InMux I__6867 (
            .O(N__29967),
            .I(N__29805));
    InMux I__6866 (
            .O(N__29966),
            .I(N__29805));
    CascadeMux I__6865 (
            .O(N__29965),
            .I(N__29797));
    InMux I__6864 (
            .O(N__29964),
            .I(N__29782));
    InMux I__6863 (
            .O(N__29961),
            .I(N__29782));
    InMux I__6862 (
            .O(N__29958),
            .I(N__29782));
    InMux I__6861 (
            .O(N__29957),
            .I(N__29782));
    InMux I__6860 (
            .O(N__29956),
            .I(N__29782));
    CascadeMux I__6859 (
            .O(N__29955),
            .I(N__29771));
    InMux I__6858 (
            .O(N__29954),
            .I(N__29763));
    InMux I__6857 (
            .O(N__29953),
            .I(N__29760));
    LocalMux I__6856 (
            .O(N__29942),
            .I(N__29756));
    InMux I__6855 (
            .O(N__29939),
            .I(N__29743));
    InMux I__6854 (
            .O(N__29936),
            .I(N__29743));
    InMux I__6853 (
            .O(N__29933),
            .I(N__29743));
    InMux I__6852 (
            .O(N__29932),
            .I(N__29743));
    InMux I__6851 (
            .O(N__29931),
            .I(N__29743));
    InMux I__6850 (
            .O(N__29930),
            .I(N__29743));
    InMux I__6849 (
            .O(N__29929),
            .I(N__29740));
    InMux I__6848 (
            .O(N__29928),
            .I(N__29735));
    InMux I__6847 (
            .O(N__29927),
            .I(N__29735));
    InMux I__6846 (
            .O(N__29926),
            .I(N__29730));
    InMux I__6845 (
            .O(N__29925),
            .I(N__29730));
    InMux I__6844 (
            .O(N__29924),
            .I(N__29727));
    InMux I__6843 (
            .O(N__29923),
            .I(N__29724));
    LocalMux I__6842 (
            .O(N__29908),
            .I(N__29721));
    Span4Mux_h I__6841 (
            .O(N__29905),
            .I(N__29714));
    LocalMux I__6840 (
            .O(N__29894),
            .I(N__29714));
    LocalMux I__6839 (
            .O(N__29887),
            .I(N__29714));
    InMux I__6838 (
            .O(N__29886),
            .I(N__29705));
    InMux I__6837 (
            .O(N__29885),
            .I(N__29705));
    InMux I__6836 (
            .O(N__29884),
            .I(N__29705));
    InMux I__6835 (
            .O(N__29883),
            .I(N__29702));
    InMux I__6834 (
            .O(N__29882),
            .I(N__29694));
    InMux I__6833 (
            .O(N__29879),
            .I(N__29685));
    InMux I__6832 (
            .O(N__29876),
            .I(N__29685));
    InMux I__6831 (
            .O(N__29875),
            .I(N__29685));
    InMux I__6830 (
            .O(N__29874),
            .I(N__29685));
    InMux I__6829 (
            .O(N__29873),
            .I(N__29676));
    InMux I__6828 (
            .O(N__29872),
            .I(N__29676));
    InMux I__6827 (
            .O(N__29871),
            .I(N__29676));
    InMux I__6826 (
            .O(N__29870),
            .I(N__29676));
    InMux I__6825 (
            .O(N__29867),
            .I(N__29671));
    InMux I__6824 (
            .O(N__29866),
            .I(N__29671));
    InMux I__6823 (
            .O(N__29863),
            .I(N__29660));
    InMux I__6822 (
            .O(N__29862),
            .I(N__29660));
    InMux I__6821 (
            .O(N__29861),
            .I(N__29660));
    InMux I__6820 (
            .O(N__29860),
            .I(N__29660));
    InMux I__6819 (
            .O(N__29859),
            .I(N__29660));
    LocalMux I__6818 (
            .O(N__29846),
            .I(N__29657));
    CascadeMux I__6817 (
            .O(N__29845),
            .I(N__29639));
    CascadeMux I__6816 (
            .O(N__29844),
            .I(N__29636));
    CascadeMux I__6815 (
            .O(N__29843),
            .I(N__29628));
    InMux I__6814 (
            .O(N__29842),
            .I(N__29620));
    InMux I__6813 (
            .O(N__29841),
            .I(N__29617));
    InMux I__6812 (
            .O(N__29840),
            .I(N__29611));
    InMux I__6811 (
            .O(N__29839),
            .I(N__29604));
    InMux I__6810 (
            .O(N__29838),
            .I(N__29604));
    InMux I__6809 (
            .O(N__29837),
            .I(N__29604));
    LocalMux I__6808 (
            .O(N__29830),
            .I(N__29599));
    LocalMux I__6807 (
            .O(N__29825),
            .I(N__29599));
    LocalMux I__6806 (
            .O(N__29816),
            .I(N__29594));
    LocalMux I__6805 (
            .O(N__29805),
            .I(N__29594));
    InMux I__6804 (
            .O(N__29804),
            .I(N__29587));
    InMux I__6803 (
            .O(N__29803),
            .I(N__29587));
    InMux I__6802 (
            .O(N__29802),
            .I(N__29587));
    InMux I__6801 (
            .O(N__29801),
            .I(N__29572));
    InMux I__6800 (
            .O(N__29800),
            .I(N__29572));
    InMux I__6799 (
            .O(N__29797),
            .I(N__29572));
    InMux I__6798 (
            .O(N__29796),
            .I(N__29572));
    InMux I__6797 (
            .O(N__29795),
            .I(N__29572));
    InMux I__6796 (
            .O(N__29794),
            .I(N__29572));
    InMux I__6795 (
            .O(N__29793),
            .I(N__29572));
    LocalMux I__6794 (
            .O(N__29782),
            .I(N__29567));
    InMux I__6793 (
            .O(N__29781),
            .I(N__29560));
    InMux I__6792 (
            .O(N__29780),
            .I(N__29560));
    InMux I__6791 (
            .O(N__29779),
            .I(N__29560));
    InMux I__6790 (
            .O(N__29778),
            .I(N__29551));
    InMux I__6789 (
            .O(N__29777),
            .I(N__29551));
    InMux I__6788 (
            .O(N__29776),
            .I(N__29551));
    InMux I__6787 (
            .O(N__29775),
            .I(N__29551));
    InMux I__6786 (
            .O(N__29774),
            .I(N__29536));
    InMux I__6785 (
            .O(N__29771),
            .I(N__29536));
    InMux I__6784 (
            .O(N__29770),
            .I(N__29536));
    InMux I__6783 (
            .O(N__29769),
            .I(N__29536));
    InMux I__6782 (
            .O(N__29768),
            .I(N__29536));
    InMux I__6781 (
            .O(N__29767),
            .I(N__29536));
    InMux I__6780 (
            .O(N__29766),
            .I(N__29536));
    LocalMux I__6779 (
            .O(N__29763),
            .I(N__29531));
    LocalMux I__6778 (
            .O(N__29760),
            .I(N__29531));
    InMux I__6777 (
            .O(N__29759),
            .I(N__29528));
    Span4Mux_v I__6776 (
            .O(N__29756),
            .I(N__29521));
    LocalMux I__6775 (
            .O(N__29743),
            .I(N__29521));
    LocalMux I__6774 (
            .O(N__29740),
            .I(N__29521));
    LocalMux I__6773 (
            .O(N__29735),
            .I(N__29508));
    LocalMux I__6772 (
            .O(N__29730),
            .I(N__29508));
    LocalMux I__6771 (
            .O(N__29727),
            .I(N__29508));
    LocalMux I__6770 (
            .O(N__29724),
            .I(N__29508));
    Span4Mux_h I__6769 (
            .O(N__29721),
            .I(N__29508));
    Span4Mux_v I__6768 (
            .O(N__29714),
            .I(N__29508));
    InMux I__6767 (
            .O(N__29713),
            .I(N__29503));
    InMux I__6766 (
            .O(N__29712),
            .I(N__29503));
    LocalMux I__6765 (
            .O(N__29705),
            .I(N__29498));
    LocalMux I__6764 (
            .O(N__29702),
            .I(N__29498));
    CascadeMux I__6763 (
            .O(N__29701),
            .I(N__29494));
    CascadeMux I__6762 (
            .O(N__29700),
            .I(N__29489));
    InMux I__6761 (
            .O(N__29699),
            .I(N__29482));
    InMux I__6760 (
            .O(N__29698),
            .I(N__29477));
    InMux I__6759 (
            .O(N__29697),
            .I(N__29477));
    LocalMux I__6758 (
            .O(N__29694),
            .I(N__29472));
    LocalMux I__6757 (
            .O(N__29685),
            .I(N__29472));
    LocalMux I__6756 (
            .O(N__29676),
            .I(N__29467));
    LocalMux I__6755 (
            .O(N__29671),
            .I(N__29467));
    LocalMux I__6754 (
            .O(N__29660),
            .I(N__29464));
    Span4Mux_v I__6753 (
            .O(N__29657),
            .I(N__29461));
    InMux I__6752 (
            .O(N__29656),
            .I(N__29452));
    InMux I__6751 (
            .O(N__29655),
            .I(N__29452));
    InMux I__6750 (
            .O(N__29654),
            .I(N__29452));
    InMux I__6749 (
            .O(N__29653),
            .I(N__29452));
    InMux I__6748 (
            .O(N__29652),
            .I(N__29447));
    InMux I__6747 (
            .O(N__29651),
            .I(N__29447));
    InMux I__6746 (
            .O(N__29650),
            .I(N__29444));
    InMux I__6745 (
            .O(N__29649),
            .I(N__29437));
    InMux I__6744 (
            .O(N__29648),
            .I(N__29437));
    InMux I__6743 (
            .O(N__29647),
            .I(N__29437));
    InMux I__6742 (
            .O(N__29646),
            .I(N__29428));
    InMux I__6741 (
            .O(N__29645),
            .I(N__29428));
    InMux I__6740 (
            .O(N__29644),
            .I(N__29428));
    InMux I__6739 (
            .O(N__29643),
            .I(N__29428));
    InMux I__6738 (
            .O(N__29642),
            .I(N__29425));
    InMux I__6737 (
            .O(N__29639),
            .I(N__29414));
    InMux I__6736 (
            .O(N__29636),
            .I(N__29414));
    InMux I__6735 (
            .O(N__29635),
            .I(N__29414));
    InMux I__6734 (
            .O(N__29634),
            .I(N__29414));
    InMux I__6733 (
            .O(N__29633),
            .I(N__29414));
    InMux I__6732 (
            .O(N__29632),
            .I(N__29409));
    InMux I__6731 (
            .O(N__29631),
            .I(N__29409));
    InMux I__6730 (
            .O(N__29628),
            .I(N__29400));
    InMux I__6729 (
            .O(N__29627),
            .I(N__29400));
    InMux I__6728 (
            .O(N__29626),
            .I(N__29400));
    InMux I__6727 (
            .O(N__29625),
            .I(N__29400));
    InMux I__6726 (
            .O(N__29624),
            .I(N__29397));
    CascadeMux I__6725 (
            .O(N__29623),
            .I(N__29390));
    LocalMux I__6724 (
            .O(N__29620),
            .I(N__29384));
    LocalMux I__6723 (
            .O(N__29617),
            .I(N__29381));
    InMux I__6722 (
            .O(N__29616),
            .I(N__29375));
    InMux I__6721 (
            .O(N__29615),
            .I(N__29375));
    InMux I__6720 (
            .O(N__29614),
            .I(N__29372));
    LocalMux I__6719 (
            .O(N__29611),
            .I(N__29359));
    LocalMux I__6718 (
            .O(N__29604),
            .I(N__29359));
    Span4Mux_v I__6717 (
            .O(N__29599),
            .I(N__29359));
    Span4Mux_v I__6716 (
            .O(N__29594),
            .I(N__29359));
    LocalMux I__6715 (
            .O(N__29587),
            .I(N__29359));
    LocalMux I__6714 (
            .O(N__29572),
            .I(N__29359));
    InMux I__6713 (
            .O(N__29571),
            .I(N__29353));
    InMux I__6712 (
            .O(N__29570),
            .I(N__29353));
    Span4Mux_v I__6711 (
            .O(N__29567),
            .I(N__29332));
    LocalMux I__6710 (
            .O(N__29560),
            .I(N__29332));
    LocalMux I__6709 (
            .O(N__29551),
            .I(N__29332));
    LocalMux I__6708 (
            .O(N__29536),
            .I(N__29332));
    Span4Mux_v I__6707 (
            .O(N__29531),
            .I(N__29332));
    LocalMux I__6706 (
            .O(N__29528),
            .I(N__29332));
    Span4Mux_v I__6705 (
            .O(N__29521),
            .I(N__29332));
    Span4Mux_h I__6704 (
            .O(N__29508),
            .I(N__29332));
    LocalMux I__6703 (
            .O(N__29503),
            .I(N__29332));
    Span4Mux_v I__6702 (
            .O(N__29498),
            .I(N__29332));
    InMux I__6701 (
            .O(N__29497),
            .I(N__29325));
    InMux I__6700 (
            .O(N__29494),
            .I(N__29325));
    InMux I__6699 (
            .O(N__29493),
            .I(N__29325));
    InMux I__6698 (
            .O(N__29492),
            .I(N__29322));
    InMux I__6697 (
            .O(N__29489),
            .I(N__29311));
    InMux I__6696 (
            .O(N__29488),
            .I(N__29311));
    InMux I__6695 (
            .O(N__29487),
            .I(N__29311));
    InMux I__6694 (
            .O(N__29486),
            .I(N__29311));
    InMux I__6693 (
            .O(N__29485),
            .I(N__29311));
    LocalMux I__6692 (
            .O(N__29482),
            .I(N__29288));
    LocalMux I__6691 (
            .O(N__29477),
            .I(N__29288));
    Span4Mux_v I__6690 (
            .O(N__29472),
            .I(N__29288));
    Span4Mux_v I__6689 (
            .O(N__29467),
            .I(N__29288));
    Span4Mux_v I__6688 (
            .O(N__29464),
            .I(N__29288));
    Span4Mux_h I__6687 (
            .O(N__29461),
            .I(N__29288));
    LocalMux I__6686 (
            .O(N__29452),
            .I(N__29288));
    LocalMux I__6685 (
            .O(N__29447),
            .I(N__29288));
    LocalMux I__6684 (
            .O(N__29444),
            .I(N__29288));
    LocalMux I__6683 (
            .O(N__29437),
            .I(N__29288));
    LocalMux I__6682 (
            .O(N__29428),
            .I(N__29288));
    LocalMux I__6681 (
            .O(N__29425),
            .I(N__29279));
    LocalMux I__6680 (
            .O(N__29414),
            .I(N__29279));
    LocalMux I__6679 (
            .O(N__29409),
            .I(N__29279));
    LocalMux I__6678 (
            .O(N__29400),
            .I(N__29279));
    LocalMux I__6677 (
            .O(N__29397),
            .I(N__29276));
    InMux I__6676 (
            .O(N__29396),
            .I(N__29273));
    InMux I__6675 (
            .O(N__29395),
            .I(N__29270));
    InMux I__6674 (
            .O(N__29394),
            .I(N__29267));
    InMux I__6673 (
            .O(N__29393),
            .I(N__29258));
    InMux I__6672 (
            .O(N__29390),
            .I(N__29258));
    InMux I__6671 (
            .O(N__29389),
            .I(N__29258));
    InMux I__6670 (
            .O(N__29388),
            .I(N__29258));
    InMux I__6669 (
            .O(N__29387),
            .I(N__29255));
    Span4Mux_v I__6668 (
            .O(N__29384),
            .I(N__29251));
    Span4Mux_v I__6667 (
            .O(N__29381),
            .I(N__29248));
    InMux I__6666 (
            .O(N__29380),
            .I(N__29245));
    LocalMux I__6665 (
            .O(N__29375),
            .I(N__29238));
    LocalMux I__6664 (
            .O(N__29372),
            .I(N__29238));
    Span4Mux_h I__6663 (
            .O(N__29359),
            .I(N__29238));
    InMux I__6662 (
            .O(N__29358),
            .I(N__29235));
    LocalMux I__6661 (
            .O(N__29353),
            .I(N__29230));
    Sp12to4 I__6660 (
            .O(N__29332),
            .I(N__29230));
    LocalMux I__6659 (
            .O(N__29325),
            .I(N__29219));
    LocalMux I__6658 (
            .O(N__29322),
            .I(N__29219));
    LocalMux I__6657 (
            .O(N__29311),
            .I(N__29219));
    Span4Mux_h I__6656 (
            .O(N__29288),
            .I(N__29219));
    Span4Mux_s2_h I__6655 (
            .O(N__29279),
            .I(N__29219));
    Span4Mux_v I__6654 (
            .O(N__29276),
            .I(N__29216));
    LocalMux I__6653 (
            .O(N__29273),
            .I(N__29213));
    LocalMux I__6652 (
            .O(N__29270),
            .I(N__29206));
    LocalMux I__6651 (
            .O(N__29267),
            .I(N__29206));
    LocalMux I__6650 (
            .O(N__29258),
            .I(N__29206));
    LocalMux I__6649 (
            .O(N__29255),
            .I(N__29203));
    InMux I__6648 (
            .O(N__29254),
            .I(N__29200));
    Span4Mux_s0_v I__6647 (
            .O(N__29251),
            .I(N__29195));
    Span4Mux_v I__6646 (
            .O(N__29248),
            .I(N__29195));
    LocalMux I__6645 (
            .O(N__29245),
            .I(N__29184));
    Sp12to4 I__6644 (
            .O(N__29238),
            .I(N__29184));
    LocalMux I__6643 (
            .O(N__29235),
            .I(N__29184));
    Span12Mux_s2_h I__6642 (
            .O(N__29230),
            .I(N__29184));
    Sp12to4 I__6641 (
            .O(N__29219),
            .I(N__29184));
    Span4Mux_v I__6640 (
            .O(N__29216),
            .I(N__29179));
    Span4Mux_s3_h I__6639 (
            .O(N__29213),
            .I(N__29179));
    Span12Mux_v I__6638 (
            .O(N__29206),
            .I(N__29176));
    Span12Mux_v I__6637 (
            .O(N__29203),
            .I(N__29173));
    LocalMux I__6636 (
            .O(N__29200),
            .I(N__29166));
    Sp12to4 I__6635 (
            .O(N__29195),
            .I(N__29166));
    Span12Mux_v I__6634 (
            .O(N__29184),
            .I(N__29166));
    Odrv4 I__6633 (
            .O(N__29179),
            .I(rx_data_ready));
    Odrv12 I__6632 (
            .O(N__29176),
            .I(rx_data_ready));
    Odrv12 I__6631 (
            .O(N__29173),
            .I(rx_data_ready));
    Odrv12 I__6630 (
            .O(N__29166),
            .I(rx_data_ready));
    InMux I__6629 (
            .O(N__29157),
            .I(N__29154));
    LocalMux I__6628 (
            .O(N__29154),
            .I(N__29151));
    Span4Mux_h I__6627 (
            .O(N__29151),
            .I(N__29148));
    Span4Mux_v I__6626 (
            .O(N__29148),
            .I(N__29144));
    InMux I__6625 (
            .O(N__29147),
            .I(N__29141));
    Odrv4 I__6624 (
            .O(N__29144),
            .I(data_in_19_0));
    LocalMux I__6623 (
            .O(N__29141),
            .I(data_in_19_0));
    InMux I__6622 (
            .O(N__29136),
            .I(N__29133));
    LocalMux I__6621 (
            .O(N__29133),
            .I(N__29130));
    Span4Mux_h I__6620 (
            .O(N__29130),
            .I(N__29127));
    Span4Mux_h I__6619 (
            .O(N__29127),
            .I(N__29123));
    InMux I__6618 (
            .O(N__29126),
            .I(N__29120));
    Odrv4 I__6617 (
            .O(N__29123),
            .I(data_in_18_0));
    LocalMux I__6616 (
            .O(N__29120),
            .I(data_in_18_0));
    InMux I__6615 (
            .O(N__29115),
            .I(N__29112));
    LocalMux I__6614 (
            .O(N__29112),
            .I(N__29109));
    Span4Mux_v I__6613 (
            .O(N__29109),
            .I(N__29104));
    InMux I__6612 (
            .O(N__29108),
            .I(N__29101));
    InMux I__6611 (
            .O(N__29107),
            .I(N__29098));
    Span4Mux_h I__6610 (
            .O(N__29104),
            .I(N__29093));
    LocalMux I__6609 (
            .O(N__29101),
            .I(N__29088));
    LocalMux I__6608 (
            .O(N__29098),
            .I(N__29088));
    InMux I__6607 (
            .O(N__29097),
            .I(N__29085));
    InMux I__6606 (
            .O(N__29096),
            .I(N__29082));
    Odrv4 I__6605 (
            .O(N__29093),
            .I(rand_data_12));
    Odrv4 I__6604 (
            .O(N__29088),
            .I(rand_data_12));
    LocalMux I__6603 (
            .O(N__29085),
            .I(rand_data_12));
    LocalMux I__6602 (
            .O(N__29082),
            .I(rand_data_12));
    CEMux I__6601 (
            .O(N__29073),
            .I(N__29059));
    CEMux I__6600 (
            .O(N__29072),
            .I(N__29049));
    CascadeMux I__6599 (
            .O(N__29071),
            .I(N__29043));
    InMux I__6598 (
            .O(N__29070),
            .I(N__29039));
    CascadeMux I__6597 (
            .O(N__29069),
            .I(N__29036));
    CascadeMux I__6596 (
            .O(N__29068),
            .I(N__29033));
    CEMux I__6595 (
            .O(N__29067),
            .I(N__29027));
    CEMux I__6594 (
            .O(N__29066),
            .I(N__29022));
    CascadeMux I__6593 (
            .O(N__29065),
            .I(N__29016));
    InMux I__6592 (
            .O(N__29064),
            .I(N__29000));
    CascadeMux I__6591 (
            .O(N__29063),
            .I(N__28993));
    CascadeMux I__6590 (
            .O(N__29062),
            .I(N__28987));
    LocalMux I__6589 (
            .O(N__29059),
            .I(N__28981));
    InMux I__6588 (
            .O(N__29058),
            .I(N__28976));
    InMux I__6587 (
            .O(N__29057),
            .I(N__28976));
    InMux I__6586 (
            .O(N__29056),
            .I(N__28973));
    CascadeMux I__6585 (
            .O(N__29055),
            .I(N__28969));
    CascadeMux I__6584 (
            .O(N__29054),
            .I(N__28963));
    CascadeMux I__6583 (
            .O(N__29053),
            .I(N__28958));
    CascadeMux I__6582 (
            .O(N__29052),
            .I(N__28954));
    LocalMux I__6581 (
            .O(N__29049),
            .I(N__28950));
    CEMux I__6580 (
            .O(N__29048),
            .I(N__28947));
    CEMux I__6579 (
            .O(N__29047),
            .I(N__28944));
    InMux I__6578 (
            .O(N__29046),
            .I(N__28937));
    InMux I__6577 (
            .O(N__29043),
            .I(N__28937));
    InMux I__6576 (
            .O(N__29042),
            .I(N__28937));
    LocalMux I__6575 (
            .O(N__29039),
            .I(N__28934));
    InMux I__6574 (
            .O(N__29036),
            .I(N__28925));
    InMux I__6573 (
            .O(N__29033),
            .I(N__28925));
    InMux I__6572 (
            .O(N__29032),
            .I(N__28925));
    InMux I__6571 (
            .O(N__29031),
            .I(N__28925));
    CEMux I__6570 (
            .O(N__29030),
            .I(N__28921));
    LocalMux I__6569 (
            .O(N__29027),
            .I(N__28918));
    CEMux I__6568 (
            .O(N__29026),
            .I(N__28915));
    CEMux I__6567 (
            .O(N__29025),
            .I(N__28912));
    LocalMux I__6566 (
            .O(N__29022),
            .I(N__28909));
    CEMux I__6565 (
            .O(N__29021),
            .I(N__28906));
    InMux I__6564 (
            .O(N__29020),
            .I(N__28897));
    InMux I__6563 (
            .O(N__29019),
            .I(N__28897));
    InMux I__6562 (
            .O(N__29016),
            .I(N__28897));
    InMux I__6561 (
            .O(N__29015),
            .I(N__28897));
    CascadeMux I__6560 (
            .O(N__29014),
            .I(N__28893));
    CascadeMux I__6559 (
            .O(N__29013),
            .I(N__28889));
    InMux I__6558 (
            .O(N__29012),
            .I(N__28886));
    CascadeMux I__6557 (
            .O(N__29011),
            .I(N__28882));
    CascadeMux I__6556 (
            .O(N__29010),
            .I(N__28878));
    CEMux I__6555 (
            .O(N__29009),
            .I(N__28874));
    CascadeMux I__6554 (
            .O(N__29008),
            .I(N__28870));
    CascadeMux I__6553 (
            .O(N__29007),
            .I(N__28864));
    CascadeMux I__6552 (
            .O(N__29006),
            .I(N__28860));
    CascadeMux I__6551 (
            .O(N__29005),
            .I(N__28857));
    CEMux I__6550 (
            .O(N__29004),
            .I(N__28845));
    CEMux I__6549 (
            .O(N__29003),
            .I(N__28842));
    LocalMux I__6548 (
            .O(N__29000),
            .I(N__28839));
    InMux I__6547 (
            .O(N__28999),
            .I(N__28834));
    InMux I__6546 (
            .O(N__28998),
            .I(N__28834));
    CEMux I__6545 (
            .O(N__28997),
            .I(N__28831));
    CEMux I__6544 (
            .O(N__28996),
            .I(N__28828));
    InMux I__6543 (
            .O(N__28993),
            .I(N__28823));
    InMux I__6542 (
            .O(N__28992),
            .I(N__28823));
    InMux I__6541 (
            .O(N__28991),
            .I(N__28814));
    InMux I__6540 (
            .O(N__28990),
            .I(N__28814));
    InMux I__6539 (
            .O(N__28987),
            .I(N__28814));
    InMux I__6538 (
            .O(N__28986),
            .I(N__28814));
    InMux I__6537 (
            .O(N__28985),
            .I(N__28809));
    InMux I__6536 (
            .O(N__28984),
            .I(N__28809));
    Span4Mux_h I__6535 (
            .O(N__28981),
            .I(N__28802));
    LocalMux I__6534 (
            .O(N__28976),
            .I(N__28802));
    LocalMux I__6533 (
            .O(N__28973),
            .I(N__28802));
    InMux I__6532 (
            .O(N__28972),
            .I(N__28799));
    InMux I__6531 (
            .O(N__28969),
            .I(N__28794));
    InMux I__6530 (
            .O(N__28968),
            .I(N__28794));
    InMux I__6529 (
            .O(N__28967),
            .I(N__28791));
    InMux I__6528 (
            .O(N__28966),
            .I(N__28784));
    InMux I__6527 (
            .O(N__28963),
            .I(N__28784));
    InMux I__6526 (
            .O(N__28962),
            .I(N__28784));
    InMux I__6525 (
            .O(N__28961),
            .I(N__28773));
    InMux I__6524 (
            .O(N__28958),
            .I(N__28773));
    InMux I__6523 (
            .O(N__28957),
            .I(N__28773));
    InMux I__6522 (
            .O(N__28954),
            .I(N__28773));
    InMux I__6521 (
            .O(N__28953),
            .I(N__28773));
    Span4Mux_s1_v I__6520 (
            .O(N__28950),
            .I(N__28769));
    LocalMux I__6519 (
            .O(N__28947),
            .I(N__28764));
    LocalMux I__6518 (
            .O(N__28944),
            .I(N__28764));
    LocalMux I__6517 (
            .O(N__28937),
            .I(N__28761));
    Span4Mux_v I__6516 (
            .O(N__28934),
            .I(N__28756));
    LocalMux I__6515 (
            .O(N__28925),
            .I(N__28756));
    InMux I__6514 (
            .O(N__28924),
            .I(N__28753));
    LocalMux I__6513 (
            .O(N__28921),
            .I(N__28739));
    Span4Mux_s1_h I__6512 (
            .O(N__28918),
            .I(N__28734));
    LocalMux I__6511 (
            .O(N__28915),
            .I(N__28734));
    LocalMux I__6510 (
            .O(N__28912),
            .I(N__28731));
    Span4Mux_s1_h I__6509 (
            .O(N__28909),
            .I(N__28728));
    LocalMux I__6508 (
            .O(N__28906),
            .I(N__28723));
    LocalMux I__6507 (
            .O(N__28897),
            .I(N__28723));
    InMux I__6506 (
            .O(N__28896),
            .I(N__28714));
    InMux I__6505 (
            .O(N__28893),
            .I(N__28714));
    InMux I__6504 (
            .O(N__28892),
            .I(N__28714));
    InMux I__6503 (
            .O(N__28889),
            .I(N__28714));
    LocalMux I__6502 (
            .O(N__28886),
            .I(N__28711));
    InMux I__6501 (
            .O(N__28885),
            .I(N__28700));
    InMux I__6500 (
            .O(N__28882),
            .I(N__28700));
    InMux I__6499 (
            .O(N__28881),
            .I(N__28700));
    InMux I__6498 (
            .O(N__28878),
            .I(N__28700));
    InMux I__6497 (
            .O(N__28877),
            .I(N__28700));
    LocalMux I__6496 (
            .O(N__28874),
            .I(N__28697));
    InMux I__6495 (
            .O(N__28873),
            .I(N__28690));
    InMux I__6494 (
            .O(N__28870),
            .I(N__28690));
    InMux I__6493 (
            .O(N__28869),
            .I(N__28690));
    InMux I__6492 (
            .O(N__28868),
            .I(N__28685));
    InMux I__6491 (
            .O(N__28867),
            .I(N__28685));
    InMux I__6490 (
            .O(N__28864),
            .I(N__28674));
    InMux I__6489 (
            .O(N__28863),
            .I(N__28674));
    InMux I__6488 (
            .O(N__28860),
            .I(N__28674));
    InMux I__6487 (
            .O(N__28857),
            .I(N__28674));
    InMux I__6486 (
            .O(N__28856),
            .I(N__28674));
    CascadeMux I__6485 (
            .O(N__28855),
            .I(N__28669));
    CascadeMux I__6484 (
            .O(N__28854),
            .I(N__28666));
    CascadeMux I__6483 (
            .O(N__28853),
            .I(N__28662));
    CascadeMux I__6482 (
            .O(N__28852),
            .I(N__28659));
    CascadeMux I__6481 (
            .O(N__28851),
            .I(N__28655));
    CascadeMux I__6480 (
            .O(N__28850),
            .I(N__28651));
    CascadeMux I__6479 (
            .O(N__28849),
            .I(N__28648));
    CascadeMux I__6478 (
            .O(N__28848),
            .I(N__28644));
    LocalMux I__6477 (
            .O(N__28845),
            .I(N__28639));
    LocalMux I__6476 (
            .O(N__28842),
            .I(N__28636));
    Span4Mux_s3_h I__6475 (
            .O(N__28839),
            .I(N__28633));
    LocalMux I__6474 (
            .O(N__28834),
            .I(N__28630));
    LocalMux I__6473 (
            .O(N__28831),
            .I(N__28613));
    LocalMux I__6472 (
            .O(N__28828),
            .I(N__28613));
    LocalMux I__6471 (
            .O(N__28823),
            .I(N__28613));
    LocalMux I__6470 (
            .O(N__28814),
            .I(N__28613));
    LocalMux I__6469 (
            .O(N__28809),
            .I(N__28613));
    Span4Mux_h I__6468 (
            .O(N__28802),
            .I(N__28613));
    LocalMux I__6467 (
            .O(N__28799),
            .I(N__28613));
    LocalMux I__6466 (
            .O(N__28794),
            .I(N__28613));
    LocalMux I__6465 (
            .O(N__28791),
            .I(N__28606));
    LocalMux I__6464 (
            .O(N__28784),
            .I(N__28606));
    LocalMux I__6463 (
            .O(N__28773),
            .I(N__28606));
    InMux I__6462 (
            .O(N__28772),
            .I(N__28603));
    Span4Mux_v I__6461 (
            .O(N__28769),
            .I(N__28592));
    Span4Mux_v I__6460 (
            .O(N__28764),
            .I(N__28592));
    Span4Mux_v I__6459 (
            .O(N__28761),
            .I(N__28592));
    Span4Mux_h I__6458 (
            .O(N__28756),
            .I(N__28592));
    LocalMux I__6457 (
            .O(N__28753),
            .I(N__28592));
    InMux I__6456 (
            .O(N__28752),
            .I(N__28589));
    CascadeMux I__6455 (
            .O(N__28751),
            .I(N__28586));
    CascadeMux I__6454 (
            .O(N__28750),
            .I(N__28582));
    CascadeMux I__6453 (
            .O(N__28749),
            .I(N__28579));
    CascadeMux I__6452 (
            .O(N__28748),
            .I(N__28574));
    CascadeMux I__6451 (
            .O(N__28747),
            .I(N__28571));
    CascadeMux I__6450 (
            .O(N__28746),
            .I(N__28568));
    CascadeMux I__6449 (
            .O(N__28745),
            .I(N__28564));
    CascadeMux I__6448 (
            .O(N__28744),
            .I(N__28560));
    CascadeMux I__6447 (
            .O(N__28743),
            .I(N__28554));
    CascadeMux I__6446 (
            .O(N__28742),
            .I(N__28551));
    Span4Mux_h I__6445 (
            .O(N__28739),
            .I(N__28547));
    Span4Mux_h I__6444 (
            .O(N__28734),
            .I(N__28542));
    Span4Mux_h I__6443 (
            .O(N__28731),
            .I(N__28542));
    Span4Mux_h I__6442 (
            .O(N__28728),
            .I(N__28531));
    Span4Mux_s3_v I__6441 (
            .O(N__28723),
            .I(N__28531));
    LocalMux I__6440 (
            .O(N__28714),
            .I(N__28531));
    Span4Mux_v I__6439 (
            .O(N__28711),
            .I(N__28531));
    LocalMux I__6438 (
            .O(N__28700),
            .I(N__28531));
    Span4Mux_h I__6437 (
            .O(N__28697),
            .I(N__28526));
    LocalMux I__6436 (
            .O(N__28690),
            .I(N__28526));
    LocalMux I__6435 (
            .O(N__28685),
            .I(N__28521));
    LocalMux I__6434 (
            .O(N__28674),
            .I(N__28521));
    InMux I__6433 (
            .O(N__28673),
            .I(N__28518));
    InMux I__6432 (
            .O(N__28672),
            .I(N__28503));
    InMux I__6431 (
            .O(N__28669),
            .I(N__28503));
    InMux I__6430 (
            .O(N__28666),
            .I(N__28503));
    InMux I__6429 (
            .O(N__28665),
            .I(N__28503));
    InMux I__6428 (
            .O(N__28662),
            .I(N__28503));
    InMux I__6427 (
            .O(N__28659),
            .I(N__28503));
    InMux I__6426 (
            .O(N__28658),
            .I(N__28503));
    InMux I__6425 (
            .O(N__28655),
            .I(N__28486));
    InMux I__6424 (
            .O(N__28654),
            .I(N__28486));
    InMux I__6423 (
            .O(N__28651),
            .I(N__28486));
    InMux I__6422 (
            .O(N__28648),
            .I(N__28486));
    InMux I__6421 (
            .O(N__28647),
            .I(N__28486));
    InMux I__6420 (
            .O(N__28644),
            .I(N__28486));
    InMux I__6419 (
            .O(N__28643),
            .I(N__28486));
    InMux I__6418 (
            .O(N__28642),
            .I(N__28486));
    Span4Mux_s3_h I__6417 (
            .O(N__28639),
            .I(N__28471));
    Span4Mux_s3_h I__6416 (
            .O(N__28636),
            .I(N__28471));
    Span4Mux_v I__6415 (
            .O(N__28633),
            .I(N__28471));
    Span4Mux_v I__6414 (
            .O(N__28630),
            .I(N__28471));
    Span4Mux_v I__6413 (
            .O(N__28613),
            .I(N__28471));
    Span4Mux_h I__6412 (
            .O(N__28606),
            .I(N__28471));
    LocalMux I__6411 (
            .O(N__28603),
            .I(N__28471));
    Span4Mux_h I__6410 (
            .O(N__28592),
            .I(N__28466));
    LocalMux I__6409 (
            .O(N__28589),
            .I(N__28466));
    InMux I__6408 (
            .O(N__28586),
            .I(N__28455));
    InMux I__6407 (
            .O(N__28585),
            .I(N__28455));
    InMux I__6406 (
            .O(N__28582),
            .I(N__28455));
    InMux I__6405 (
            .O(N__28579),
            .I(N__28455));
    InMux I__6404 (
            .O(N__28578),
            .I(N__28455));
    InMux I__6403 (
            .O(N__28577),
            .I(N__28440));
    InMux I__6402 (
            .O(N__28574),
            .I(N__28440));
    InMux I__6401 (
            .O(N__28571),
            .I(N__28440));
    InMux I__6400 (
            .O(N__28568),
            .I(N__28440));
    InMux I__6399 (
            .O(N__28567),
            .I(N__28440));
    InMux I__6398 (
            .O(N__28564),
            .I(N__28440));
    InMux I__6397 (
            .O(N__28563),
            .I(N__28440));
    InMux I__6396 (
            .O(N__28560),
            .I(N__28425));
    InMux I__6395 (
            .O(N__28559),
            .I(N__28425));
    InMux I__6394 (
            .O(N__28558),
            .I(N__28425));
    InMux I__6393 (
            .O(N__28557),
            .I(N__28425));
    InMux I__6392 (
            .O(N__28554),
            .I(N__28425));
    InMux I__6391 (
            .O(N__28551),
            .I(N__28425));
    InMux I__6390 (
            .O(N__28550),
            .I(N__28425));
    Odrv4 I__6389 (
            .O(N__28547),
            .I(n4806));
    Odrv4 I__6388 (
            .O(N__28542),
            .I(n4806));
    Odrv4 I__6387 (
            .O(N__28531),
            .I(n4806));
    Odrv4 I__6386 (
            .O(N__28526),
            .I(n4806));
    Odrv4 I__6385 (
            .O(N__28521),
            .I(n4806));
    LocalMux I__6384 (
            .O(N__28518),
            .I(n4806));
    LocalMux I__6383 (
            .O(N__28503),
            .I(n4806));
    LocalMux I__6382 (
            .O(N__28486),
            .I(n4806));
    Odrv4 I__6381 (
            .O(N__28471),
            .I(n4806));
    Odrv4 I__6380 (
            .O(N__28466),
            .I(n4806));
    LocalMux I__6379 (
            .O(N__28455),
            .I(n4806));
    LocalMux I__6378 (
            .O(N__28440),
            .I(n4806));
    LocalMux I__6377 (
            .O(N__28425),
            .I(n4806));
    InMux I__6376 (
            .O(N__28398),
            .I(N__28392));
    InMux I__6375 (
            .O(N__28397),
            .I(N__28389));
    InMux I__6374 (
            .O(N__28396),
            .I(N__28385));
    InMux I__6373 (
            .O(N__28395),
            .I(N__28382));
    LocalMux I__6372 (
            .O(N__28392),
            .I(N__28378));
    LocalMux I__6371 (
            .O(N__28389),
            .I(N__28375));
    InMux I__6370 (
            .O(N__28388),
            .I(N__28372));
    LocalMux I__6369 (
            .O(N__28385),
            .I(N__28367));
    LocalMux I__6368 (
            .O(N__28382),
            .I(N__28367));
    InMux I__6367 (
            .O(N__28381),
            .I(N__28364));
    Span4Mux_h I__6366 (
            .O(N__28378),
            .I(N__28361));
    Span12Mux_s6_v I__6365 (
            .O(N__28375),
            .I(N__28358));
    LocalMux I__6364 (
            .O(N__28372),
            .I(N__28353));
    Span4Mux_v I__6363 (
            .O(N__28367),
            .I(N__28353));
    LocalMux I__6362 (
            .O(N__28364),
            .I(data_in_field_88));
    Odrv4 I__6361 (
            .O(N__28361),
            .I(data_in_field_88));
    Odrv12 I__6360 (
            .O(N__28358),
            .I(data_in_field_88));
    Odrv4 I__6359 (
            .O(N__28353),
            .I(data_in_field_88));
    InMux I__6358 (
            .O(N__28344),
            .I(N__28340));
    InMux I__6357 (
            .O(N__28343),
            .I(N__28337));
    LocalMux I__6356 (
            .O(N__28340),
            .I(N__28334));
    LocalMux I__6355 (
            .O(N__28337),
            .I(N__28331));
    Span12Mux_s10_h I__6354 (
            .O(N__28334),
            .I(N__28328));
    Span4Mux_h I__6353 (
            .O(N__28331),
            .I(N__28325));
    Odrv12 I__6352 (
            .O(N__28328),
            .I(\c0.n4292 ));
    Odrv4 I__6351 (
            .O(N__28325),
            .I(\c0.n4292 ));
    InMux I__6350 (
            .O(N__28320),
            .I(N__28316));
    InMux I__6349 (
            .O(N__28319),
            .I(N__28313));
    LocalMux I__6348 (
            .O(N__28316),
            .I(N__28310));
    LocalMux I__6347 (
            .O(N__28313),
            .I(\c0.n8957 ));
    Odrv4 I__6346 (
            .O(N__28310),
            .I(\c0.n8957 ));
    CascadeMux I__6345 (
            .O(N__28305),
            .I(N__28302));
    InMux I__6344 (
            .O(N__28302),
            .I(N__28296));
    InMux I__6343 (
            .O(N__28301),
            .I(N__28293));
    CascadeMux I__6342 (
            .O(N__28300),
            .I(N__28289));
    CascadeMux I__6341 (
            .O(N__28299),
            .I(N__28286));
    LocalMux I__6340 (
            .O(N__28296),
            .I(N__28283));
    LocalMux I__6339 (
            .O(N__28293),
            .I(N__28280));
    InMux I__6338 (
            .O(N__28292),
            .I(N__28277));
    InMux I__6337 (
            .O(N__28289),
            .I(N__28274));
    InMux I__6336 (
            .O(N__28286),
            .I(N__28271));
    Span4Mux_s3_h I__6335 (
            .O(N__28283),
            .I(N__28268));
    Span12Mux_h I__6334 (
            .O(N__28280),
            .I(N__28265));
    LocalMux I__6333 (
            .O(N__28277),
            .I(N__28262));
    LocalMux I__6332 (
            .O(N__28274),
            .I(N__28259));
    LocalMux I__6331 (
            .O(N__28271),
            .I(\c0.data_in_field_27 ));
    Odrv4 I__6330 (
            .O(N__28268),
            .I(\c0.data_in_field_27 ));
    Odrv12 I__6329 (
            .O(N__28265),
            .I(\c0.data_in_field_27 ));
    Odrv4 I__6328 (
            .O(N__28262),
            .I(\c0.data_in_field_27 ));
    Odrv4 I__6327 (
            .O(N__28259),
            .I(\c0.data_in_field_27 ));
    InMux I__6326 (
            .O(N__28248),
            .I(N__28245));
    LocalMux I__6325 (
            .O(N__28245),
            .I(N__28241));
    CascadeMux I__6324 (
            .O(N__28244),
            .I(N__28237));
    Span4Mux_v I__6323 (
            .O(N__28241),
            .I(N__28234));
    InMux I__6322 (
            .O(N__28240),
            .I(N__28231));
    InMux I__6321 (
            .O(N__28237),
            .I(N__28226));
    Span4Mux_h I__6320 (
            .O(N__28234),
            .I(N__28223));
    LocalMux I__6319 (
            .O(N__28231),
            .I(N__28220));
    InMux I__6318 (
            .O(N__28230),
            .I(N__28215));
    InMux I__6317 (
            .O(N__28229),
            .I(N__28215));
    LocalMux I__6316 (
            .O(N__28226),
            .I(\c0.data_in_field_25 ));
    Odrv4 I__6315 (
            .O(N__28223),
            .I(\c0.data_in_field_25 ));
    Odrv4 I__6314 (
            .O(N__28220),
            .I(\c0.data_in_field_25 ));
    LocalMux I__6313 (
            .O(N__28215),
            .I(\c0.data_in_field_25 ));
    InMux I__6312 (
            .O(N__28206),
            .I(N__28203));
    LocalMux I__6311 (
            .O(N__28203),
            .I(N__28200));
    Sp12to4 I__6310 (
            .O(N__28200),
            .I(N__28197));
    Span12Mux_s8_h I__6309 (
            .O(N__28197),
            .I(N__28194));
    Odrv12 I__6308 (
            .O(N__28194),
            .I(\c0.n8871 ));
    InMux I__6307 (
            .O(N__28191),
            .I(N__28188));
    LocalMux I__6306 (
            .O(N__28188),
            .I(n26));
    InMux I__6305 (
            .O(N__28185),
            .I(bfn_11_27_0_));
    InMux I__6304 (
            .O(N__28182),
            .I(N__28179));
    LocalMux I__6303 (
            .O(N__28179),
            .I(n25_adj_1722));
    InMux I__6302 (
            .O(N__28176),
            .I(n8130));
    InMux I__6301 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__6300 (
            .O(N__28170),
            .I(n1));
    InMux I__6299 (
            .O(N__28167),
            .I(N__28160));
    CascadeMux I__6298 (
            .O(N__28166),
            .I(N__28153));
    InMux I__6297 (
            .O(N__28165),
            .I(N__28146));
    InMux I__6296 (
            .O(N__28164),
            .I(N__28146));
    InMux I__6295 (
            .O(N__28163),
            .I(N__28143));
    LocalMux I__6294 (
            .O(N__28160),
            .I(N__28140));
    InMux I__6293 (
            .O(N__28159),
            .I(N__28133));
    InMux I__6292 (
            .O(N__28158),
            .I(N__28133));
    InMux I__6291 (
            .O(N__28157),
            .I(N__28133));
    InMux I__6290 (
            .O(N__28156),
            .I(N__28124));
    InMux I__6289 (
            .O(N__28153),
            .I(N__28124));
    InMux I__6288 (
            .O(N__28152),
            .I(N__28124));
    InMux I__6287 (
            .O(N__28151),
            .I(N__28124));
    LocalMux I__6286 (
            .O(N__28146),
            .I(N__28121));
    LocalMux I__6285 (
            .O(N__28143),
            .I(N__28118));
    Sp12to4 I__6284 (
            .O(N__28140),
            .I(N__28111));
    LocalMux I__6283 (
            .O(N__28133),
            .I(N__28111));
    LocalMux I__6282 (
            .O(N__28124),
            .I(N__28111));
    Span4Mux_h I__6281 (
            .O(N__28121),
            .I(N__28108));
    Span4Mux_h I__6280 (
            .O(N__28118),
            .I(N__28105));
    Odrv12 I__6279 (
            .O(N__28111),
            .I(r_Rx_Data));
    Odrv4 I__6278 (
            .O(N__28108),
            .I(r_Rx_Data));
    Odrv4 I__6277 (
            .O(N__28105),
            .I(r_Rx_Data));
    InMux I__6276 (
            .O(N__28098),
            .I(N__28092));
    InMux I__6275 (
            .O(N__28097),
            .I(N__28092));
    LocalMux I__6274 (
            .O(N__28092),
            .I(\c0.rx.r_SM_Main_2_N_1543_0 ));
    InMux I__6273 (
            .O(N__28089),
            .I(N__28086));
    LocalMux I__6272 (
            .O(N__28086),
            .I(n9300));
    InMux I__6271 (
            .O(N__28083),
            .I(N__28080));
    LocalMux I__6270 (
            .O(N__28080),
            .I(N__28076));
    CascadeMux I__6269 (
            .O(N__28079),
            .I(N__28073));
    Span4Mux_h I__6268 (
            .O(N__28076),
            .I(N__28070));
    InMux I__6267 (
            .O(N__28073),
            .I(N__28066));
    Span4Mux_h I__6266 (
            .O(N__28070),
            .I(N__28063));
    InMux I__6265 (
            .O(N__28069),
            .I(N__28060));
    LocalMux I__6264 (
            .O(N__28066),
            .I(\c0.data_in_field_24 ));
    Odrv4 I__6263 (
            .O(N__28063),
            .I(\c0.data_in_field_24 ));
    LocalMux I__6262 (
            .O(N__28060),
            .I(\c0.data_in_field_24 ));
    InMux I__6261 (
            .O(N__28053),
            .I(N__28050));
    LocalMux I__6260 (
            .O(N__28050),
            .I(N__28047));
    Span4Mux_h I__6259 (
            .O(N__28047),
            .I(N__28044));
    Span4Mux_h I__6258 (
            .O(N__28044),
            .I(N__28038));
    InMux I__6257 (
            .O(N__28043),
            .I(N__28033));
    InMux I__6256 (
            .O(N__28042),
            .I(N__28033));
    InMux I__6255 (
            .O(N__28041),
            .I(N__28030));
    Odrv4 I__6254 (
            .O(N__28038),
            .I(\c0.data_in_field_16 ));
    LocalMux I__6253 (
            .O(N__28033),
            .I(\c0.data_in_field_16 ));
    LocalMux I__6252 (
            .O(N__28030),
            .I(\c0.data_in_field_16 ));
    InMux I__6251 (
            .O(N__28023),
            .I(N__28020));
    LocalMux I__6250 (
            .O(N__28020),
            .I(N__28016));
    CascadeMux I__6249 (
            .O(N__28019),
            .I(N__28013));
    Span4Mux_h I__6248 (
            .O(N__28016),
            .I(N__28010));
    InMux I__6247 (
            .O(N__28013),
            .I(N__28006));
    Span4Mux_h I__6246 (
            .O(N__28010),
            .I(N__28003));
    InMux I__6245 (
            .O(N__28009),
            .I(N__28000));
    LocalMux I__6244 (
            .O(N__28006),
            .I(\c0.data_in_field_8 ));
    Odrv4 I__6243 (
            .O(N__28003),
            .I(\c0.data_in_field_8 ));
    LocalMux I__6242 (
            .O(N__28000),
            .I(\c0.data_in_field_8 ));
    InMux I__6241 (
            .O(N__27993),
            .I(N__27990));
    LocalMux I__6240 (
            .O(N__27990),
            .I(N__27986));
    InMux I__6239 (
            .O(N__27989),
            .I(N__27983));
    Span4Mux_h I__6238 (
            .O(N__27986),
            .I(N__27979));
    LocalMux I__6237 (
            .O(N__27983),
            .I(N__27976));
    InMux I__6236 (
            .O(N__27982),
            .I(N__27972));
    Span4Mux_h I__6235 (
            .O(N__27979),
            .I(N__27967));
    Span4Mux_v I__6234 (
            .O(N__27976),
            .I(N__27967));
    InMux I__6233 (
            .O(N__27975),
            .I(N__27964));
    LocalMux I__6232 (
            .O(N__27972),
            .I(\c0.data_in_field_0 ));
    Odrv4 I__6231 (
            .O(N__27967),
            .I(\c0.data_in_field_0 ));
    LocalMux I__6230 (
            .O(N__27964),
            .I(\c0.data_in_field_0 ));
    CascadeMux I__6229 (
            .O(N__27957),
            .I(\c0.n9446_cascade_ ));
    InMux I__6228 (
            .O(N__27954),
            .I(N__27951));
    LocalMux I__6227 (
            .O(N__27951),
            .I(N__27948));
    Span4Mux_h I__6226 (
            .O(N__27948),
            .I(N__27945));
    Span4Mux_h I__6225 (
            .O(N__27945),
            .I(N__27942));
    Odrv4 I__6224 (
            .O(N__27942),
            .I(\c0.n9228 ));
    CascadeMux I__6223 (
            .O(N__27939),
            .I(\c0.n9449_cascade_ ));
    InMux I__6222 (
            .O(N__27936),
            .I(N__27933));
    LocalMux I__6221 (
            .O(N__27933),
            .I(N__27927));
    InMux I__6220 (
            .O(N__27932),
            .I(N__27923));
    InMux I__6219 (
            .O(N__27931),
            .I(N__27920));
    InMux I__6218 (
            .O(N__27930),
            .I(N__27917));
    Span4Mux_v I__6217 (
            .O(N__27927),
            .I(N__27914));
    InMux I__6216 (
            .O(N__27926),
            .I(N__27911));
    LocalMux I__6215 (
            .O(N__27923),
            .I(N__27906));
    LocalMux I__6214 (
            .O(N__27920),
            .I(N__27906));
    LocalMux I__6213 (
            .O(N__27917),
            .I(data_in_field_80));
    Odrv4 I__6212 (
            .O(N__27914),
            .I(data_in_field_80));
    LocalMux I__6211 (
            .O(N__27911),
            .I(data_in_field_80));
    Odrv12 I__6210 (
            .O(N__27906),
            .I(data_in_field_80));
    InMux I__6209 (
            .O(N__27897),
            .I(N__27893));
    InMux I__6208 (
            .O(N__27896),
            .I(N__27890));
    LocalMux I__6207 (
            .O(N__27893),
            .I(N__27887));
    LocalMux I__6206 (
            .O(N__27890),
            .I(N__27883));
    Span4Mux_h I__6205 (
            .O(N__27887),
            .I(N__27880));
    InMux I__6204 (
            .O(N__27886),
            .I(N__27876));
    Span4Mux_h I__6203 (
            .O(N__27883),
            .I(N__27873));
    Span4Mux_h I__6202 (
            .O(N__27880),
            .I(N__27870));
    InMux I__6201 (
            .O(N__27879),
            .I(N__27867));
    LocalMux I__6200 (
            .O(N__27876),
            .I(data_in_field_72));
    Odrv4 I__6199 (
            .O(N__27873),
            .I(data_in_field_72));
    Odrv4 I__6198 (
            .O(N__27870),
            .I(data_in_field_72));
    LocalMux I__6197 (
            .O(N__27867),
            .I(data_in_field_72));
    CascadeMux I__6196 (
            .O(N__27858),
            .I(\c0.n9740_cascade_ ));
    InMux I__6195 (
            .O(N__27855),
            .I(N__27850));
    InMux I__6194 (
            .O(N__27854),
            .I(N__27847));
    InMux I__6193 (
            .O(N__27853),
            .I(N__27844));
    LocalMux I__6192 (
            .O(N__27850),
            .I(N__27840));
    LocalMux I__6191 (
            .O(N__27847),
            .I(N__27835));
    LocalMux I__6190 (
            .O(N__27844),
            .I(N__27835));
    InMux I__6189 (
            .O(N__27843),
            .I(N__27832));
    Span4Mux_h I__6188 (
            .O(N__27840),
            .I(N__27827));
    Span4Mux_v I__6187 (
            .O(N__27835),
            .I(N__27827));
    LocalMux I__6186 (
            .O(N__27832),
            .I(data_in_field_64));
    Odrv4 I__6185 (
            .O(N__27827),
            .I(data_in_field_64));
    InMux I__6184 (
            .O(N__27822),
            .I(N__27819));
    LocalMux I__6183 (
            .O(N__27819),
            .I(N__27816));
    Span4Mux_v I__6182 (
            .O(N__27816),
            .I(N__27813));
    Span4Mux_h I__6181 (
            .O(N__27813),
            .I(N__27810));
    Odrv4 I__6180 (
            .O(N__27810),
            .I(\c0.n9234 ));
    CascadeMux I__6179 (
            .O(N__27807),
            .I(\c0.n9231_cascade_ ));
    InMux I__6178 (
            .O(N__27804),
            .I(N__27801));
    LocalMux I__6177 (
            .O(N__27801),
            .I(\c0.n9728 ));
    CascadeMux I__6176 (
            .O(N__27798),
            .I(n6_adj_1751_cascade_));
    CascadeMux I__6175 (
            .O(N__27795),
            .I(n30_cascade_));
    InMux I__6174 (
            .O(N__27792),
            .I(N__27788));
    InMux I__6173 (
            .O(N__27791),
            .I(N__27781));
    LocalMux I__6172 (
            .O(N__27788),
            .I(N__27778));
    InMux I__6171 (
            .O(N__27787),
            .I(N__27775));
    InMux I__6170 (
            .O(N__27786),
            .I(N__27772));
    InMux I__6169 (
            .O(N__27785),
            .I(N__27767));
    InMux I__6168 (
            .O(N__27784),
            .I(N__27767));
    LocalMux I__6167 (
            .O(N__27781),
            .I(N__27764));
    Span4Mux_v I__6166 (
            .O(N__27778),
            .I(N__27760));
    LocalMux I__6165 (
            .O(N__27775),
            .I(N__27757));
    LocalMux I__6164 (
            .O(N__27772),
            .I(N__27754));
    LocalMux I__6163 (
            .O(N__27767),
            .I(N__27749));
    Span4Mux_s2_h I__6162 (
            .O(N__27764),
            .I(N__27749));
    InMux I__6161 (
            .O(N__27763),
            .I(N__27746));
    Span4Mux_h I__6160 (
            .O(N__27760),
            .I(N__27739));
    Span4Mux_v I__6159 (
            .O(N__27757),
            .I(N__27739));
    Span4Mux_v I__6158 (
            .O(N__27754),
            .I(N__27739));
    Span4Mux_h I__6157 (
            .O(N__27749),
            .I(N__27736));
    LocalMux I__6156 (
            .O(N__27746),
            .I(data_in_field_97));
    Odrv4 I__6155 (
            .O(N__27739),
            .I(data_in_field_97));
    Odrv4 I__6154 (
            .O(N__27736),
            .I(data_in_field_97));
    InMux I__6153 (
            .O(N__27729),
            .I(N__27724));
    InMux I__6152 (
            .O(N__27728),
            .I(N__27721));
    InMux I__6151 (
            .O(N__27727),
            .I(N__27717));
    LocalMux I__6150 (
            .O(N__27724),
            .I(N__27714));
    LocalMux I__6149 (
            .O(N__27721),
            .I(N__27711));
    InMux I__6148 (
            .O(N__27720),
            .I(N__27708));
    LocalMux I__6147 (
            .O(N__27717),
            .I(N__27705));
    Span4Mux_s3_h I__6146 (
            .O(N__27714),
            .I(N__27698));
    Span4Mux_s2_v I__6145 (
            .O(N__27711),
            .I(N__27698));
    LocalMux I__6144 (
            .O(N__27708),
            .I(N__27693));
    Span4Mux_s2_v I__6143 (
            .O(N__27705),
            .I(N__27693));
    InMux I__6142 (
            .O(N__27704),
            .I(N__27690));
    InMux I__6141 (
            .O(N__27703),
            .I(N__27687));
    Span4Mux_v I__6140 (
            .O(N__27698),
            .I(N__27684));
    Span4Mux_v I__6139 (
            .O(N__27693),
            .I(N__27679));
    LocalMux I__6138 (
            .O(N__27690),
            .I(N__27679));
    LocalMux I__6137 (
            .O(N__27687),
            .I(data_in_field_95));
    Odrv4 I__6136 (
            .O(N__27684),
            .I(data_in_field_95));
    Odrv4 I__6135 (
            .O(N__27679),
            .I(data_in_field_95));
    InMux I__6134 (
            .O(N__27672),
            .I(N__27668));
    InMux I__6133 (
            .O(N__27671),
            .I(N__27663));
    LocalMux I__6132 (
            .O(N__27668),
            .I(N__27660));
    InMux I__6131 (
            .O(N__27667),
            .I(N__27654));
    InMux I__6130 (
            .O(N__27666),
            .I(N__27654));
    LocalMux I__6129 (
            .O(N__27663),
            .I(N__27651));
    Span4Mux_s3_v I__6128 (
            .O(N__27660),
            .I(N__27648));
    InMux I__6127 (
            .O(N__27659),
            .I(N__27643));
    LocalMux I__6126 (
            .O(N__27654),
            .I(N__27640));
    Span4Mux_s3_v I__6125 (
            .O(N__27651),
            .I(N__27635));
    Span4Mux_h I__6124 (
            .O(N__27648),
            .I(N__27635));
    InMux I__6123 (
            .O(N__27647),
            .I(N__27630));
    InMux I__6122 (
            .O(N__27646),
            .I(N__27630));
    LocalMux I__6121 (
            .O(N__27643),
            .I(data_in_field_96));
    Odrv12 I__6120 (
            .O(N__27640),
            .I(data_in_field_96));
    Odrv4 I__6119 (
            .O(N__27635),
            .I(data_in_field_96));
    LocalMux I__6118 (
            .O(N__27630),
            .I(data_in_field_96));
    CascadeMux I__6117 (
            .O(N__27621),
            .I(N__27618));
    InMux I__6116 (
            .O(N__27618),
            .I(N__27615));
    LocalMux I__6115 (
            .O(N__27615),
            .I(N__27611));
    InMux I__6114 (
            .O(N__27614),
            .I(N__27608));
    Span4Mux_h I__6113 (
            .O(N__27611),
            .I(N__27605));
    LocalMux I__6112 (
            .O(N__27608),
            .I(N__27602));
    Span4Mux_v I__6111 (
            .O(N__27605),
            .I(N__27599));
    Odrv4 I__6110 (
            .O(N__27602),
            .I(\c0.n4296 ));
    Odrv4 I__6109 (
            .O(N__27599),
            .I(\c0.n4296 ));
    CascadeMux I__6108 (
            .O(N__27594),
            .I(N__27591));
    InMux I__6107 (
            .O(N__27591),
            .I(N__27588));
    LocalMux I__6106 (
            .O(N__27588),
            .I(\c0.rx.n12 ));
    IoInMux I__6105 (
            .O(N__27585),
            .I(N__27582));
    LocalMux I__6104 (
            .O(N__27582),
            .I(N__27579));
    Span4Mux_s0_v I__6103 (
            .O(N__27579),
            .I(N__27576));
    Span4Mux_h I__6102 (
            .O(N__27576),
            .I(N__27573));
    Odrv4 I__6101 (
            .O(N__27573),
            .I(tx_enable));
    CascadeMux I__6100 (
            .O(N__27570),
            .I(N__27565));
    InMux I__6099 (
            .O(N__27569),
            .I(N__27562));
    InMux I__6098 (
            .O(N__27568),
            .I(N__27557));
    InMux I__6097 (
            .O(N__27565),
            .I(N__27557));
    LocalMux I__6096 (
            .O(N__27562),
            .I(n2185));
    LocalMux I__6095 (
            .O(N__27557),
            .I(n2185));
    InMux I__6094 (
            .O(N__27552),
            .I(N__27548));
    InMux I__6093 (
            .O(N__27551),
            .I(N__27545));
    LocalMux I__6092 (
            .O(N__27548),
            .I(N__27539));
    LocalMux I__6091 (
            .O(N__27545),
            .I(N__27539));
    InMux I__6090 (
            .O(N__27544),
            .I(N__27536));
    Span4Mux_h I__6089 (
            .O(N__27539),
            .I(N__27530));
    LocalMux I__6088 (
            .O(N__27536),
            .I(N__27530));
    CascadeMux I__6087 (
            .O(N__27535),
            .I(N__27526));
    Span4Mux_v I__6086 (
            .O(N__27530),
            .I(N__27523));
    InMux I__6085 (
            .O(N__27529),
            .I(N__27520));
    InMux I__6084 (
            .O(N__27526),
            .I(N__27515));
    Span4Mux_v I__6083 (
            .O(N__27523),
            .I(N__27512));
    LocalMux I__6082 (
            .O(N__27520),
            .I(N__27509));
    InMux I__6081 (
            .O(N__27519),
            .I(N__27504));
    InMux I__6080 (
            .O(N__27518),
            .I(N__27504));
    LocalMux I__6079 (
            .O(N__27515),
            .I(r_Bit_Index_2_adj_1731));
    Odrv4 I__6078 (
            .O(N__27512),
            .I(r_Bit_Index_2_adj_1731));
    Odrv12 I__6077 (
            .O(N__27509),
            .I(r_Bit_Index_2_adj_1731));
    LocalMux I__6076 (
            .O(N__27504),
            .I(r_Bit_Index_2_adj_1731));
    CascadeMux I__6075 (
            .O(N__27495),
            .I(n7415_cascade_));
    CascadeMux I__6074 (
            .O(N__27492),
            .I(n9301_cascade_));
    InMux I__6073 (
            .O(N__27489),
            .I(N__27486));
    LocalMux I__6072 (
            .O(N__27486),
            .I(N__27483));
    Odrv12 I__6071 (
            .O(N__27483),
            .I(\c0.n20_adj_1642 ));
    CascadeMux I__6070 (
            .O(N__27480),
            .I(n12_adj_1753_cascade_));
    CascadeMux I__6069 (
            .O(N__27477),
            .I(r_SM_Main_2_N_1537_2_cascade_));
    InMux I__6068 (
            .O(N__27474),
            .I(N__27470));
    InMux I__6067 (
            .O(N__27473),
            .I(N__27467));
    LocalMux I__6066 (
            .O(N__27470),
            .I(N__27464));
    LocalMux I__6065 (
            .O(N__27467),
            .I(N__27461));
    Span4Mux_h I__6064 (
            .O(N__27464),
            .I(N__27458));
    Span12Mux_s9_h I__6063 (
            .O(N__27461),
            .I(N__27455));
    Span4Mux_v I__6062 (
            .O(N__27458),
            .I(N__27452));
    Odrv12 I__6061 (
            .O(N__27455),
            .I(\c0.rx.n4090 ));
    Odrv4 I__6060 (
            .O(N__27452),
            .I(\c0.rx.n4090 ));
    InMux I__6059 (
            .O(N__27447),
            .I(N__27444));
    LocalMux I__6058 (
            .O(N__27444),
            .I(N__27441));
    Span4Mux_h I__6057 (
            .O(N__27441),
            .I(N__27437));
    InMux I__6056 (
            .O(N__27440),
            .I(N__27434));
    Odrv4 I__6055 (
            .O(N__27437),
            .I(\c0.rx.n7393 ));
    LocalMux I__6054 (
            .O(N__27434),
            .I(\c0.rx.n7393 ));
    InMux I__6053 (
            .O(N__27429),
            .I(N__27426));
    LocalMux I__6052 (
            .O(N__27426),
            .I(N__27422));
    InMux I__6051 (
            .O(N__27425),
            .I(N__27419));
    Span4Mux_s3_v I__6050 (
            .O(N__27422),
            .I(N__27416));
    LocalMux I__6049 (
            .O(N__27419),
            .I(N__27413));
    Span4Mux_h I__6048 (
            .O(N__27416),
            .I(N__27405));
    Span4Mux_s3_v I__6047 (
            .O(N__27413),
            .I(N__27405));
    InMux I__6046 (
            .O(N__27412),
            .I(N__27400));
    InMux I__6045 (
            .O(N__27411),
            .I(N__27400));
    InMux I__6044 (
            .O(N__27410),
            .I(N__27397));
    Odrv4 I__6043 (
            .O(N__27405),
            .I(data_in_field_122));
    LocalMux I__6042 (
            .O(N__27400),
            .I(data_in_field_122));
    LocalMux I__6041 (
            .O(N__27397),
            .I(data_in_field_122));
    InMux I__6040 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__6039 (
            .O(N__27387),
            .I(N__27384));
    Span4Mux_h I__6038 (
            .O(N__27384),
            .I(N__27381));
    Span4Mux_v I__6037 (
            .O(N__27381),
            .I(N__27378));
    Odrv4 I__6036 (
            .O(N__27378),
            .I(\c0.n4537 ));
    CascadeMux I__6035 (
            .O(N__27375),
            .I(\c0.rx.r_SM_Main_2_N_1543_0_cascade_ ));
    InMux I__6034 (
            .O(N__27372),
            .I(N__27368));
    InMux I__6033 (
            .O(N__27371),
            .I(N__27365));
    LocalMux I__6032 (
            .O(N__27368),
            .I(N__27362));
    LocalMux I__6031 (
            .O(N__27365),
            .I(N__27359));
    Span4Mux_v I__6030 (
            .O(N__27362),
            .I(N__27356));
    Span4Mux_h I__6029 (
            .O(N__27359),
            .I(N__27353));
    Span4Mux_h I__6028 (
            .O(N__27356),
            .I(N__27350));
    Odrv4 I__6027 (
            .O(N__27353),
            .I(\c0.n8782 ));
    Odrv4 I__6026 (
            .O(N__27350),
            .I(\c0.n8782 ));
    CascadeMux I__6025 (
            .O(N__27345),
            .I(N__27342));
    InMux I__6024 (
            .O(N__27342),
            .I(N__27339));
    LocalMux I__6023 (
            .O(N__27339),
            .I(N__27336));
    Span12Mux_v I__6022 (
            .O(N__27336),
            .I(N__27333));
    Odrv12 I__6021 (
            .O(N__27333),
            .I(\c0.n8807 ));
    CascadeMux I__6020 (
            .O(N__27330),
            .I(N__27324));
    InMux I__6019 (
            .O(N__27329),
            .I(N__27321));
    InMux I__6018 (
            .O(N__27328),
            .I(N__27318));
    InMux I__6017 (
            .O(N__27327),
            .I(N__27315));
    InMux I__6016 (
            .O(N__27324),
            .I(N__27312));
    LocalMux I__6015 (
            .O(N__27321),
            .I(N__27309));
    LocalMux I__6014 (
            .O(N__27318),
            .I(N__27304));
    LocalMux I__6013 (
            .O(N__27315),
            .I(N__27301));
    LocalMux I__6012 (
            .O(N__27312),
            .I(N__27298));
    Span4Mux_v I__6011 (
            .O(N__27309),
            .I(N__27295));
    InMux I__6010 (
            .O(N__27308),
            .I(N__27290));
    InMux I__6009 (
            .O(N__27307),
            .I(N__27290));
    Span4Mux_s2_v I__6008 (
            .O(N__27304),
            .I(N__27285));
    Span4Mux_s2_v I__6007 (
            .O(N__27301),
            .I(N__27285));
    Odrv12 I__6006 (
            .O(N__27298),
            .I(data_in_field_110));
    Odrv4 I__6005 (
            .O(N__27295),
            .I(data_in_field_110));
    LocalMux I__6004 (
            .O(N__27290),
            .I(data_in_field_110));
    Odrv4 I__6003 (
            .O(N__27285),
            .I(data_in_field_110));
    InMux I__6002 (
            .O(N__27276),
            .I(N__27273));
    LocalMux I__6001 (
            .O(N__27273),
            .I(\c0.n8819 ));
    CascadeMux I__6000 (
            .O(N__27270),
            .I(N__27266));
    InMux I__5999 (
            .O(N__27269),
            .I(N__27263));
    InMux I__5998 (
            .O(N__27266),
            .I(N__27260));
    LocalMux I__5997 (
            .O(N__27263),
            .I(N__27257));
    LocalMux I__5996 (
            .O(N__27260),
            .I(N__27254));
    Span4Mux_v I__5995 (
            .O(N__27257),
            .I(N__27251));
    Span4Mux_v I__5994 (
            .O(N__27254),
            .I(N__27248));
    Span4Mux_s3_h I__5993 (
            .O(N__27251),
            .I(N__27245));
    Odrv4 I__5992 (
            .O(N__27248),
            .I(\c0.n8893 ));
    Odrv4 I__5991 (
            .O(N__27245),
            .I(\c0.n8893 ));
    InMux I__5990 (
            .O(N__27240),
            .I(N__27237));
    LocalMux I__5989 (
            .O(N__27237),
            .I(N__27234));
    Span12Mux_s7_v I__5988 (
            .O(N__27234),
            .I(N__27230));
    InMux I__5987 (
            .O(N__27233),
            .I(N__27227));
    Odrv12 I__5986 (
            .O(N__27230),
            .I(\c0.n8427 ));
    LocalMux I__5985 (
            .O(N__27227),
            .I(\c0.n8427 ));
    InMux I__5984 (
            .O(N__27222),
            .I(N__27219));
    LocalMux I__5983 (
            .O(N__27219),
            .I(N__27216));
    Odrv12 I__5982 (
            .O(N__27216),
            .I(\c0.n28_adj_1612 ));
    InMux I__5981 (
            .O(N__27213),
            .I(N__27210));
    LocalMux I__5980 (
            .O(N__27210),
            .I(\c0.n26_adj_1613 ));
    CascadeMux I__5979 (
            .O(N__27207),
            .I(\c0.n27_cascade_ ));
    InMux I__5978 (
            .O(N__27204),
            .I(N__27201));
    LocalMux I__5977 (
            .O(N__27201),
            .I(N__27198));
    Odrv4 I__5976 (
            .O(N__27198),
            .I(\c0.n25_adj_1614 ));
    InMux I__5975 (
            .O(N__27195),
            .I(N__27192));
    LocalMux I__5974 (
            .O(N__27192),
            .I(N__27189));
    Odrv12 I__5973 (
            .O(N__27189),
            .I(\c0.data_in_frame_20_0 ));
    InMux I__5972 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__5971 (
            .O(N__27183),
            .I(N__27180));
    Span4Mux_v I__5970 (
            .O(N__27180),
            .I(N__27177));
    Span4Mux_h I__5969 (
            .O(N__27177),
            .I(N__27173));
    InMux I__5968 (
            .O(N__27176),
            .I(N__27170));
    Span4Mux_h I__5967 (
            .O(N__27173),
            .I(N__27167));
    LocalMux I__5966 (
            .O(N__27170),
            .I(\c0.n8995 ));
    Odrv4 I__5965 (
            .O(N__27167),
            .I(\c0.n8995 ));
    InMux I__5964 (
            .O(N__27162),
            .I(N__27156));
    InMux I__5963 (
            .O(N__27161),
            .I(N__27156));
    LocalMux I__5962 (
            .O(N__27156),
            .I(N__27153));
    Span4Mux_h I__5961 (
            .O(N__27153),
            .I(N__27150));
    Odrv4 I__5960 (
            .O(N__27150),
            .I(\c0.n8834 ));
    CascadeMux I__5959 (
            .O(N__27147),
            .I(N__27144));
    InMux I__5958 (
            .O(N__27144),
            .I(N__27141));
    LocalMux I__5957 (
            .O(N__27141),
            .I(N__27138));
    Span4Mux_h I__5956 (
            .O(N__27138),
            .I(N__27134));
    InMux I__5955 (
            .O(N__27137),
            .I(N__27131));
    Span4Mux_h I__5954 (
            .O(N__27134),
            .I(N__27128));
    LocalMux I__5953 (
            .O(N__27131),
            .I(\c0.n8924 ));
    Odrv4 I__5952 (
            .O(N__27128),
            .I(\c0.n8924 ));
    InMux I__5951 (
            .O(N__27123),
            .I(N__27120));
    LocalMux I__5950 (
            .O(N__27120),
            .I(N__27116));
    InMux I__5949 (
            .O(N__27119),
            .I(N__27113));
    Span12Mux_s10_v I__5948 (
            .O(N__27116),
            .I(N__27110));
    LocalMux I__5947 (
            .O(N__27113),
            .I(N__27107));
    Odrv12 I__5946 (
            .O(N__27110),
            .I(\c0.n8852 ));
    Odrv4 I__5945 (
            .O(N__27107),
            .I(\c0.n8852 ));
    InMux I__5944 (
            .O(N__27102),
            .I(N__27099));
    LocalMux I__5943 (
            .O(N__27099),
            .I(N__27095));
    InMux I__5942 (
            .O(N__27098),
            .I(N__27092));
    Span4Mux_h I__5941 (
            .O(N__27095),
            .I(N__27089));
    LocalMux I__5940 (
            .O(N__27092),
            .I(N__27086));
    Odrv4 I__5939 (
            .O(N__27089),
            .I(\c0.n9013 ));
    Odrv4 I__5938 (
            .O(N__27086),
            .I(\c0.n9013 ));
    InMux I__5937 (
            .O(N__27081),
            .I(N__27078));
    LocalMux I__5936 (
            .O(N__27078),
            .I(N__27074));
    InMux I__5935 (
            .O(N__27077),
            .I(N__27071));
    Span4Mux_s2_v I__5934 (
            .O(N__27074),
            .I(N__27068));
    LocalMux I__5933 (
            .O(N__27071),
            .I(N__27063));
    Span4Mux_v I__5932 (
            .O(N__27068),
            .I(N__27060));
    InMux I__5931 (
            .O(N__27067),
            .I(N__27055));
    InMux I__5930 (
            .O(N__27066),
            .I(N__27055));
    Odrv4 I__5929 (
            .O(N__27063),
            .I(data_in_field_70));
    Odrv4 I__5928 (
            .O(N__27060),
            .I(data_in_field_70));
    LocalMux I__5927 (
            .O(N__27055),
            .I(data_in_field_70));
    CascadeMux I__5926 (
            .O(N__27048),
            .I(\c0.n12_cascade_ ));
    InMux I__5925 (
            .O(N__27045),
            .I(N__27042));
    LocalMux I__5924 (
            .O(N__27042),
            .I(N__27038));
    InMux I__5923 (
            .O(N__27041),
            .I(N__27035));
    Span4Mux_v I__5922 (
            .O(N__27038),
            .I(N__27030));
    LocalMux I__5921 (
            .O(N__27035),
            .I(N__27027));
    InMux I__5920 (
            .O(N__27034),
            .I(N__27024));
    InMux I__5919 (
            .O(N__27033),
            .I(N__27021));
    Span4Mux_h I__5918 (
            .O(N__27030),
            .I(N__27016));
    Span4Mux_h I__5917 (
            .O(N__27027),
            .I(N__27016));
    LocalMux I__5916 (
            .O(N__27024),
            .I(data_in_field_112));
    LocalMux I__5915 (
            .O(N__27021),
            .I(data_in_field_112));
    Odrv4 I__5914 (
            .O(N__27016),
            .I(data_in_field_112));
    InMux I__5913 (
            .O(N__27009),
            .I(N__27006));
    LocalMux I__5912 (
            .O(N__27006),
            .I(\c0.data_in_frame_20_2 ));
    InMux I__5911 (
            .O(N__27003),
            .I(N__27000));
    LocalMux I__5910 (
            .O(N__27000),
            .I(N__26997));
    Span4Mux_v I__5909 (
            .O(N__26997),
            .I(N__26992));
    InMux I__5908 (
            .O(N__26996),
            .I(N__26987));
    InMux I__5907 (
            .O(N__26995),
            .I(N__26987));
    Odrv4 I__5906 (
            .O(N__26992),
            .I(data_in_5_2));
    LocalMux I__5905 (
            .O(N__26987),
            .I(data_in_5_2));
    InMux I__5904 (
            .O(N__26982),
            .I(N__26979));
    LocalMux I__5903 (
            .O(N__26979),
            .I(N__26975));
    InMux I__5902 (
            .O(N__26978),
            .I(N__26972));
    Span4Mux_s3_h I__5901 (
            .O(N__26975),
            .I(N__26969));
    LocalMux I__5900 (
            .O(N__26972),
            .I(N__26966));
    Span4Mux_v I__5899 (
            .O(N__26969),
            .I(N__26963));
    Span4Mux_h I__5898 (
            .O(N__26966),
            .I(N__26960));
    Span4Mux_h I__5897 (
            .O(N__26963),
            .I(N__26956));
    Span4Mux_v I__5896 (
            .O(N__26960),
            .I(N__26953));
    InMux I__5895 (
            .O(N__26959),
            .I(N__26950));
    Odrv4 I__5894 (
            .O(N__26956),
            .I(data_in_4_2));
    Odrv4 I__5893 (
            .O(N__26953),
            .I(data_in_4_2));
    LocalMux I__5892 (
            .O(N__26950),
            .I(data_in_4_2));
    InMux I__5891 (
            .O(N__26943),
            .I(N__26939));
    InMux I__5890 (
            .O(N__26942),
            .I(N__26935));
    LocalMux I__5889 (
            .O(N__26939),
            .I(N__26931));
    InMux I__5888 (
            .O(N__26938),
            .I(N__26928));
    LocalMux I__5887 (
            .O(N__26935),
            .I(N__26925));
    CascadeMux I__5886 (
            .O(N__26934),
            .I(N__26922));
    Span4Mux_h I__5885 (
            .O(N__26931),
            .I(N__26914));
    LocalMux I__5884 (
            .O(N__26928),
            .I(N__26911));
    Span12Mux_h I__5883 (
            .O(N__26925),
            .I(N__26908));
    InMux I__5882 (
            .O(N__26922),
            .I(N__26905));
    InMux I__5881 (
            .O(N__26921),
            .I(N__26898));
    InMux I__5880 (
            .O(N__26920),
            .I(N__26898));
    InMux I__5879 (
            .O(N__26919),
            .I(N__26898));
    InMux I__5878 (
            .O(N__26918),
            .I(N__26893));
    InMux I__5877 (
            .O(N__26917),
            .I(N__26893));
    Odrv4 I__5876 (
            .O(N__26914),
            .I(r_SM_Main_2_adj_1738));
    Odrv4 I__5875 (
            .O(N__26911),
            .I(r_SM_Main_2_adj_1738));
    Odrv12 I__5874 (
            .O(N__26908),
            .I(r_SM_Main_2_adj_1738));
    LocalMux I__5873 (
            .O(N__26905),
            .I(r_SM_Main_2_adj_1738));
    LocalMux I__5872 (
            .O(N__26898),
            .I(r_SM_Main_2_adj_1738));
    LocalMux I__5871 (
            .O(N__26893),
            .I(r_SM_Main_2_adj_1738));
    CEMux I__5870 (
            .O(N__26880),
            .I(N__26877));
    LocalMux I__5869 (
            .O(N__26877),
            .I(N__26873));
    CEMux I__5868 (
            .O(N__26876),
            .I(N__26870));
    Span4Mux_s1_v I__5867 (
            .O(N__26873),
            .I(N__26865));
    LocalMux I__5866 (
            .O(N__26870),
            .I(N__26865));
    Span4Mux_s1_h I__5865 (
            .O(N__26865),
            .I(N__26862));
    Span4Mux_h I__5864 (
            .O(N__26862),
            .I(N__26859));
    Span4Mux_h I__5863 (
            .O(N__26859),
            .I(N__26856));
    Odrv4 I__5862 (
            .O(N__26856),
            .I(\c0.tx2.n4880 ));
    InMux I__5861 (
            .O(N__26853),
            .I(N__26850));
    LocalMux I__5860 (
            .O(N__26850),
            .I(N__26847));
    Span4Mux_v I__5859 (
            .O(N__26847),
            .I(N__26844));
    Span4Mux_h I__5858 (
            .O(N__26844),
            .I(N__26841));
    Odrv4 I__5857 (
            .O(N__26841),
            .I(\c0.n4525 ));
    CascadeMux I__5856 (
            .O(N__26838),
            .I(N__26835));
    InMux I__5855 (
            .O(N__26835),
            .I(N__26832));
    LocalMux I__5854 (
            .O(N__26832),
            .I(N__26829));
    Span4Mux_v I__5853 (
            .O(N__26829),
            .I(N__26826));
    Odrv4 I__5852 (
            .O(N__26826),
            .I(\c0.n4244 ));
    InMux I__5851 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__5850 (
            .O(N__26820),
            .I(N__26817));
    Span4Mux_v I__5849 (
            .O(N__26817),
            .I(N__26810));
    InMux I__5848 (
            .O(N__26816),
            .I(N__26805));
    InMux I__5847 (
            .O(N__26815),
            .I(N__26805));
    InMux I__5846 (
            .O(N__26814),
            .I(N__26802));
    InMux I__5845 (
            .O(N__26813),
            .I(N__26799));
    Span4Mux_h I__5844 (
            .O(N__26810),
            .I(N__26794));
    LocalMux I__5843 (
            .O(N__26805),
            .I(N__26794));
    LocalMux I__5842 (
            .O(N__26802),
            .I(data_in_field_50));
    LocalMux I__5841 (
            .O(N__26799),
            .I(data_in_field_50));
    Odrv4 I__5840 (
            .O(N__26794),
            .I(data_in_field_50));
    InMux I__5839 (
            .O(N__26787),
            .I(N__26784));
    LocalMux I__5838 (
            .O(N__26784),
            .I(N__26780));
    InMux I__5837 (
            .O(N__26783),
            .I(N__26777));
    Odrv12 I__5836 (
            .O(N__26780),
            .I(\c0.n8918 ));
    LocalMux I__5835 (
            .O(N__26777),
            .I(\c0.n8918 ));
    CascadeMux I__5834 (
            .O(N__26772),
            .I(\c0.n8840_cascade_ ));
    InMux I__5833 (
            .O(N__26769),
            .I(N__26765));
    InMux I__5832 (
            .O(N__26768),
            .I(N__26762));
    LocalMux I__5831 (
            .O(N__26765),
            .I(\c0.n4511 ));
    LocalMux I__5830 (
            .O(N__26762),
            .I(\c0.n4511 ));
    InMux I__5829 (
            .O(N__26757),
            .I(N__26754));
    LocalMux I__5828 (
            .O(N__26754),
            .I(N__26751));
    Span12Mux_s7_h I__5827 (
            .O(N__26751),
            .I(N__26747));
    InMux I__5826 (
            .O(N__26750),
            .I(N__26744));
    Odrv12 I__5825 (
            .O(N__26747),
            .I(\c0.n4309 ));
    LocalMux I__5824 (
            .O(N__26744),
            .I(\c0.n4309 ));
    InMux I__5823 (
            .O(N__26739),
            .I(N__26735));
    InMux I__5822 (
            .O(N__26738),
            .I(N__26732));
    LocalMux I__5821 (
            .O(N__26735),
            .I(N__26729));
    LocalMux I__5820 (
            .O(N__26732),
            .I(N__26725));
    Span4Mux_h I__5819 (
            .O(N__26729),
            .I(N__26722));
    InMux I__5818 (
            .O(N__26728),
            .I(N__26718));
    Span4Mux_v I__5817 (
            .O(N__26725),
            .I(N__26714));
    Sp12to4 I__5816 (
            .O(N__26722),
            .I(N__26711));
    InMux I__5815 (
            .O(N__26721),
            .I(N__26708));
    LocalMux I__5814 (
            .O(N__26718),
            .I(N__26705));
    InMux I__5813 (
            .O(N__26717),
            .I(N__26702));
    Odrv4 I__5812 (
            .O(N__26714),
            .I(rand_data_11));
    Odrv12 I__5811 (
            .O(N__26711),
            .I(rand_data_11));
    LocalMux I__5810 (
            .O(N__26708),
            .I(rand_data_11));
    Odrv12 I__5809 (
            .O(N__26705),
            .I(rand_data_11));
    LocalMux I__5808 (
            .O(N__26702),
            .I(rand_data_11));
    CascadeMux I__5807 (
            .O(N__26691),
            .I(N__26686));
    InMux I__5806 (
            .O(N__26690),
            .I(N__26680));
    InMux I__5805 (
            .O(N__26689),
            .I(N__26680));
    InMux I__5804 (
            .O(N__26686),
            .I(N__26677));
    InMux I__5803 (
            .O(N__26685),
            .I(N__26674));
    LocalMux I__5802 (
            .O(N__26680),
            .I(N__26671));
    LocalMux I__5801 (
            .O(N__26677),
            .I(N__26668));
    LocalMux I__5800 (
            .O(N__26674),
            .I(N__26665));
    Span4Mux_v I__5799 (
            .O(N__26671),
            .I(N__26660));
    Span4Mux_s3_h I__5798 (
            .O(N__26668),
            .I(N__26660));
    Span4Mux_v I__5797 (
            .O(N__26665),
            .I(N__26656));
    Span4Mux_h I__5796 (
            .O(N__26660),
            .I(N__26651));
    InMux I__5795 (
            .O(N__26659),
            .I(N__26648));
    Sp12to4 I__5794 (
            .O(N__26656),
            .I(N__26645));
    InMux I__5793 (
            .O(N__26655),
            .I(N__26640));
    InMux I__5792 (
            .O(N__26654),
            .I(N__26640));
    Span4Mux_v I__5791 (
            .O(N__26651),
            .I(N__26637));
    LocalMux I__5790 (
            .O(N__26648),
            .I(data_in_field_123));
    Odrv12 I__5789 (
            .O(N__26645),
            .I(data_in_field_123));
    LocalMux I__5788 (
            .O(N__26640),
            .I(data_in_field_123));
    Odrv4 I__5787 (
            .O(N__26637),
            .I(data_in_field_123));
    InMux I__5786 (
            .O(N__26628),
            .I(N__26624));
    CascadeMux I__5785 (
            .O(N__26627),
            .I(N__26620));
    LocalMux I__5784 (
            .O(N__26624),
            .I(N__26616));
    InMux I__5783 (
            .O(N__26623),
            .I(N__26613));
    InMux I__5782 (
            .O(N__26620),
            .I(N__26607));
    InMux I__5781 (
            .O(N__26619),
            .I(N__26607));
    Span4Mux_h I__5780 (
            .O(N__26616),
            .I(N__26602));
    LocalMux I__5779 (
            .O(N__26613),
            .I(N__26599));
    InMux I__5778 (
            .O(N__26612),
            .I(N__26596));
    LocalMux I__5777 (
            .O(N__26607),
            .I(N__26593));
    InMux I__5776 (
            .O(N__26606),
            .I(N__26588));
    InMux I__5775 (
            .O(N__26605),
            .I(N__26585));
    Span4Mux_v I__5774 (
            .O(N__26602),
            .I(N__26578));
    Span4Mux_h I__5773 (
            .O(N__26599),
            .I(N__26578));
    LocalMux I__5772 (
            .O(N__26596),
            .I(N__26578));
    Span12Mux_s8_h I__5771 (
            .O(N__26593),
            .I(N__26575));
    InMux I__5770 (
            .O(N__26592),
            .I(N__26572));
    InMux I__5769 (
            .O(N__26591),
            .I(N__26569));
    LocalMux I__5768 (
            .O(N__26588),
            .I(data_in_field_146));
    LocalMux I__5767 (
            .O(N__26585),
            .I(data_in_field_146));
    Odrv4 I__5766 (
            .O(N__26578),
            .I(data_in_field_146));
    Odrv12 I__5765 (
            .O(N__26575),
            .I(data_in_field_146));
    LocalMux I__5764 (
            .O(N__26572),
            .I(data_in_field_146));
    LocalMux I__5763 (
            .O(N__26569),
            .I(data_in_field_146));
    InMux I__5762 (
            .O(N__26556),
            .I(N__26551));
    InMux I__5761 (
            .O(N__26555),
            .I(N__26548));
    InMux I__5760 (
            .O(N__26554),
            .I(N__26545));
    LocalMux I__5759 (
            .O(N__26551),
            .I(N__26542));
    LocalMux I__5758 (
            .O(N__26548),
            .I(N__26536));
    LocalMux I__5757 (
            .O(N__26545),
            .I(N__26536));
    Span4Mux_h I__5756 (
            .O(N__26542),
            .I(N__26533));
    CascadeMux I__5755 (
            .O(N__26541),
            .I(N__26529));
    Span4Mux_v I__5754 (
            .O(N__26536),
            .I(N__26526));
    Span4Mux_v I__5753 (
            .O(N__26533),
            .I(N__26523));
    InMux I__5752 (
            .O(N__26532),
            .I(N__26518));
    InMux I__5751 (
            .O(N__26529),
            .I(N__26518));
    Span4Mux_h I__5750 (
            .O(N__26526),
            .I(N__26515));
    Odrv4 I__5749 (
            .O(N__26523),
            .I(data_in_field_130));
    LocalMux I__5748 (
            .O(N__26518),
            .I(data_in_field_130));
    Odrv4 I__5747 (
            .O(N__26515),
            .I(data_in_field_130));
    CascadeMux I__5746 (
            .O(N__26508),
            .I(\c0.n9698_cascade_ ));
    InMux I__5745 (
            .O(N__26505),
            .I(N__26502));
    LocalMux I__5744 (
            .O(N__26502),
            .I(N__26497));
    InMux I__5743 (
            .O(N__26501),
            .I(N__26494));
    InMux I__5742 (
            .O(N__26500),
            .I(N__26491));
    Span4Mux_v I__5741 (
            .O(N__26497),
            .I(N__26486));
    LocalMux I__5740 (
            .O(N__26494),
            .I(N__26486));
    LocalMux I__5739 (
            .O(N__26491),
            .I(N__26481));
    Span4Mux_h I__5738 (
            .O(N__26486),
            .I(N__26478));
    InMux I__5737 (
            .O(N__26485),
            .I(N__26473));
    InMux I__5736 (
            .O(N__26484),
            .I(N__26473));
    Odrv4 I__5735 (
            .O(N__26481),
            .I(data_in_field_138));
    Odrv4 I__5734 (
            .O(N__26478),
            .I(data_in_field_138));
    LocalMux I__5733 (
            .O(N__26473),
            .I(data_in_field_138));
    CascadeMux I__5732 (
            .O(N__26466),
            .I(\c0.n9701_cascade_ ));
    InMux I__5731 (
            .O(N__26463),
            .I(N__26458));
    CascadeMux I__5730 (
            .O(N__26462),
            .I(N__26454));
    InMux I__5729 (
            .O(N__26461),
            .I(N__26451));
    LocalMux I__5728 (
            .O(N__26458),
            .I(N__26448));
    InMux I__5727 (
            .O(N__26457),
            .I(N__26445));
    InMux I__5726 (
            .O(N__26454),
            .I(N__26442));
    LocalMux I__5725 (
            .O(N__26451),
            .I(N__26438));
    Span4Mux_v I__5724 (
            .O(N__26448),
            .I(N__26433));
    LocalMux I__5723 (
            .O(N__26445),
            .I(N__26433));
    LocalMux I__5722 (
            .O(N__26442),
            .I(N__26430));
    InMux I__5721 (
            .O(N__26441),
            .I(N__26427));
    Span4Mux_h I__5720 (
            .O(N__26438),
            .I(N__26424));
    Span4Mux_h I__5719 (
            .O(N__26433),
            .I(N__26421));
    Span4Mux_v I__5718 (
            .O(N__26430),
            .I(N__26418));
    LocalMux I__5717 (
            .O(N__26427),
            .I(data_in_field_142));
    Odrv4 I__5716 (
            .O(N__26424),
            .I(data_in_field_142));
    Odrv4 I__5715 (
            .O(N__26421),
            .I(data_in_field_142));
    Odrv4 I__5714 (
            .O(N__26418),
            .I(data_in_field_142));
    InMux I__5713 (
            .O(N__26409),
            .I(N__26405));
    CascadeMux I__5712 (
            .O(N__26408),
            .I(N__26401));
    LocalMux I__5711 (
            .O(N__26405),
            .I(N__26398));
    InMux I__5710 (
            .O(N__26404),
            .I(N__26394));
    InMux I__5709 (
            .O(N__26401),
            .I(N__26391));
    Span4Mux_v I__5708 (
            .O(N__26398),
            .I(N__26388));
    InMux I__5707 (
            .O(N__26397),
            .I(N__26385));
    LocalMux I__5706 (
            .O(N__26394),
            .I(N__26382));
    LocalMux I__5705 (
            .O(N__26391),
            .I(N__26377));
    IoSpan4Mux I__5704 (
            .O(N__26388),
            .I(N__26374));
    LocalMux I__5703 (
            .O(N__26385),
            .I(N__26371));
    Span4Mux_s1_v I__5702 (
            .O(N__26382),
            .I(N__26368));
    InMux I__5701 (
            .O(N__26381),
            .I(N__26365));
    InMux I__5700 (
            .O(N__26380),
            .I(N__26362));
    Span4Mux_h I__5699 (
            .O(N__26377),
            .I(N__26353));
    Span4Mux_s3_h I__5698 (
            .O(N__26374),
            .I(N__26353));
    Span4Mux_v I__5697 (
            .O(N__26371),
            .I(N__26353));
    Span4Mux_v I__5696 (
            .O(N__26368),
            .I(N__26353));
    LocalMux I__5695 (
            .O(N__26365),
            .I(data_in_field_78));
    LocalMux I__5694 (
            .O(N__26362),
            .I(data_in_field_78));
    Odrv4 I__5693 (
            .O(N__26353),
            .I(data_in_field_78));
    InMux I__5692 (
            .O(N__26346),
            .I(N__26342));
    InMux I__5691 (
            .O(N__26345),
            .I(N__26339));
    LocalMux I__5690 (
            .O(N__26342),
            .I(N__26336));
    LocalMux I__5689 (
            .O(N__26339),
            .I(N__26333));
    Span4Mux_v I__5688 (
            .O(N__26336),
            .I(N__26330));
    Span4Mux_v I__5687 (
            .O(N__26333),
            .I(N__26326));
    Span4Mux_h I__5686 (
            .O(N__26330),
            .I(N__26323));
    InMux I__5685 (
            .O(N__26329),
            .I(N__26320));
    Odrv4 I__5684 (
            .O(N__26326),
            .I(\c0.n4215 ));
    Odrv4 I__5683 (
            .O(N__26323),
            .I(\c0.n4215 ));
    LocalMux I__5682 (
            .O(N__26320),
            .I(\c0.n4215 ));
    CascadeMux I__5681 (
            .O(N__26313),
            .I(N__26310));
    InMux I__5680 (
            .O(N__26310),
            .I(N__26307));
    LocalMux I__5679 (
            .O(N__26307),
            .I(N__26304));
    Span4Mux_v I__5678 (
            .O(N__26304),
            .I(N__26300));
    InMux I__5677 (
            .O(N__26303),
            .I(N__26297));
    Odrv4 I__5676 (
            .O(N__26300),
            .I(\c0.n8912 ));
    LocalMux I__5675 (
            .O(N__26297),
            .I(\c0.n8912 ));
    InMux I__5674 (
            .O(N__26292),
            .I(N__26288));
    InMux I__5673 (
            .O(N__26291),
            .I(N__26285));
    LocalMux I__5672 (
            .O(N__26288),
            .I(N__26282));
    LocalMux I__5671 (
            .O(N__26285),
            .I(N__26279));
    Odrv4 I__5670 (
            .O(N__26282),
            .I(\c0.n8954 ));
    Odrv12 I__5669 (
            .O(N__26279),
            .I(\c0.n8954 ));
    CascadeMux I__5668 (
            .O(N__26274),
            .I(\c0.n8819_cascade_ ));
    InMux I__5667 (
            .O(N__26271),
            .I(N__26268));
    LocalMux I__5666 (
            .O(N__26268),
            .I(N__26264));
    InMux I__5665 (
            .O(N__26267),
            .I(N__26261));
    Odrv4 I__5664 (
            .O(N__26264),
            .I(\c0.n4365 ));
    LocalMux I__5663 (
            .O(N__26261),
            .I(\c0.n4365 ));
    CascadeMux I__5662 (
            .O(N__26256),
            .I(\c0.n21_adj_1644_cascade_ ));
    InMux I__5661 (
            .O(N__26253),
            .I(N__26250));
    LocalMux I__5660 (
            .O(N__26250),
            .I(N__26247));
    Span4Mux_h I__5659 (
            .O(N__26247),
            .I(N__26244));
    Span4Mux_h I__5658 (
            .O(N__26244),
            .I(N__26241));
    Odrv4 I__5657 (
            .O(N__26241),
            .I(\c0.n19_adj_1643 ));
    CascadeMux I__5656 (
            .O(N__26238),
            .I(N__26235));
    InMux I__5655 (
            .O(N__26235),
            .I(N__26232));
    LocalMux I__5654 (
            .O(N__26232),
            .I(\c0.data_in_frame_19_2 ));
    InMux I__5653 (
            .O(N__26229),
            .I(N__26226));
    LocalMux I__5652 (
            .O(N__26226),
            .I(\c0.data_in_frame_19_0 ));
    InMux I__5651 (
            .O(N__26223),
            .I(N__26220));
    LocalMux I__5650 (
            .O(N__26220),
            .I(N__26216));
    InMux I__5649 (
            .O(N__26219),
            .I(N__26213));
    Span4Mux_h I__5648 (
            .O(N__26216),
            .I(N__26207));
    LocalMux I__5647 (
            .O(N__26213),
            .I(N__26207));
    InMux I__5646 (
            .O(N__26212),
            .I(N__26203));
    Span4Mux_h I__5645 (
            .O(N__26207),
            .I(N__26200));
    InMux I__5644 (
            .O(N__26206),
            .I(N__26197));
    LocalMux I__5643 (
            .O(N__26203),
            .I(data_in_field_136));
    Odrv4 I__5642 (
            .O(N__26200),
            .I(data_in_field_136));
    LocalMux I__5641 (
            .O(N__26197),
            .I(data_in_field_136));
    CascadeMux I__5640 (
            .O(N__26190),
            .I(\c0.n9536_cascade_ ));
    InMux I__5639 (
            .O(N__26187),
            .I(N__26183));
    InMux I__5638 (
            .O(N__26186),
            .I(N__26180));
    LocalMux I__5637 (
            .O(N__26183),
            .I(N__26176));
    LocalMux I__5636 (
            .O(N__26180),
            .I(N__26173));
    InMux I__5635 (
            .O(N__26179),
            .I(N__26169));
    Span4Mux_h I__5634 (
            .O(N__26176),
            .I(N__26164));
    Span4Mux_h I__5633 (
            .O(N__26173),
            .I(N__26164));
    InMux I__5632 (
            .O(N__26172),
            .I(N__26161));
    LocalMux I__5631 (
            .O(N__26169),
            .I(data_in_field_128));
    Odrv4 I__5630 (
            .O(N__26164),
            .I(data_in_field_128));
    LocalMux I__5629 (
            .O(N__26161),
            .I(data_in_field_128));
    CascadeMux I__5628 (
            .O(N__26154),
            .I(\c0.n9539_cascade_ ));
    InMux I__5627 (
            .O(N__26151),
            .I(N__26148));
    LocalMux I__5626 (
            .O(N__26148),
            .I(N__26143));
    InMux I__5625 (
            .O(N__26147),
            .I(N__26140));
    InMux I__5624 (
            .O(N__26146),
            .I(N__26137));
    Span4Mux_v I__5623 (
            .O(N__26143),
            .I(N__26132));
    LocalMux I__5622 (
            .O(N__26140),
            .I(N__26132));
    LocalMux I__5621 (
            .O(N__26137),
            .I(N__26127));
    Span4Mux_h I__5620 (
            .O(N__26132),
            .I(N__26127));
    Span4Mux_v I__5619 (
            .O(N__26127),
            .I(N__26123));
    InMux I__5618 (
            .O(N__26126),
            .I(N__26120));
    Odrv4 I__5617 (
            .O(N__26123),
            .I(rand_data_18));
    LocalMux I__5616 (
            .O(N__26120),
            .I(rand_data_18));
    InMux I__5615 (
            .O(N__26115),
            .I(N__26112));
    LocalMux I__5614 (
            .O(N__26112),
            .I(N__26109));
    Span4Mux_s2_v I__5613 (
            .O(N__26109),
            .I(N__26105));
    InMux I__5612 (
            .O(N__26108),
            .I(N__26102));
    Span4Mux_h I__5611 (
            .O(N__26105),
            .I(N__26097));
    LocalMux I__5610 (
            .O(N__26102),
            .I(N__26097));
    Span4Mux_v I__5609 (
            .O(N__26097),
            .I(N__26092));
    InMux I__5608 (
            .O(N__26096),
            .I(N__26087));
    InMux I__5607 (
            .O(N__26095),
            .I(N__26087));
    Odrv4 I__5606 (
            .O(N__26092),
            .I(data_in_field_114));
    LocalMux I__5605 (
            .O(N__26087),
            .I(data_in_field_114));
    InMux I__5604 (
            .O(N__26082),
            .I(N__26076));
    InMux I__5603 (
            .O(N__26081),
            .I(N__26073));
    InMux I__5602 (
            .O(N__26080),
            .I(N__26070));
    InMux I__5601 (
            .O(N__26079),
            .I(N__26067));
    LocalMux I__5600 (
            .O(N__26076),
            .I(N__26062));
    LocalMux I__5599 (
            .O(N__26073),
            .I(N__26062));
    LocalMux I__5598 (
            .O(N__26070),
            .I(N__26057));
    LocalMux I__5597 (
            .O(N__26067),
            .I(N__26054));
    Span4Mux_v I__5596 (
            .O(N__26062),
            .I(N__26051));
    InMux I__5595 (
            .O(N__26061),
            .I(N__26046));
    InMux I__5594 (
            .O(N__26060),
            .I(N__26046));
    Span4Mux_h I__5593 (
            .O(N__26057),
            .I(N__26043));
    Span4Mux_h I__5592 (
            .O(N__26054),
            .I(N__26038));
    Span4Mux_h I__5591 (
            .O(N__26051),
            .I(N__26038));
    LocalMux I__5590 (
            .O(N__26046),
            .I(data_in_field_144));
    Odrv4 I__5589 (
            .O(N__26043),
            .I(data_in_field_144));
    Odrv4 I__5588 (
            .O(N__26038),
            .I(data_in_field_144));
    InMux I__5587 (
            .O(N__26031),
            .I(N__26027));
    InMux I__5586 (
            .O(N__26030),
            .I(N__26024));
    LocalMux I__5585 (
            .O(N__26027),
            .I(N__26021));
    LocalMux I__5584 (
            .O(N__26024),
            .I(N__26018));
    Span4Mux_h I__5583 (
            .O(N__26021),
            .I(N__26015));
    Span4Mux_v I__5582 (
            .O(N__26018),
            .I(N__26012));
    Span4Mux_h I__5581 (
            .O(N__26015),
            .I(N__26009));
    Odrv4 I__5580 (
            .O(N__26012),
            .I(\c0.n8971 ));
    Odrv4 I__5579 (
            .O(N__26009),
            .I(\c0.n8971 ));
    InMux I__5578 (
            .O(N__26004),
            .I(N__26001));
    LocalMux I__5577 (
            .O(N__26001),
            .I(\c0.n6_adj_1628 ));
    InMux I__5576 (
            .O(N__25998),
            .I(N__25994));
    InMux I__5575 (
            .O(N__25997),
            .I(N__25991));
    LocalMux I__5574 (
            .O(N__25994),
            .I(N__25988));
    LocalMux I__5573 (
            .O(N__25991),
            .I(N__25984));
    Span4Mux_h I__5572 (
            .O(N__25988),
            .I(N__25981));
    InMux I__5571 (
            .O(N__25987),
            .I(N__25978));
    Span4Mux_v I__5570 (
            .O(N__25984),
            .I(N__25973));
    Span4Mux_v I__5569 (
            .O(N__25981),
            .I(N__25970));
    LocalMux I__5568 (
            .O(N__25978),
            .I(N__25967));
    InMux I__5567 (
            .O(N__25977),
            .I(N__25964));
    InMux I__5566 (
            .O(N__25976),
            .I(N__25961));
    Odrv4 I__5565 (
            .O(N__25973),
            .I(rand_data_0));
    Odrv4 I__5564 (
            .O(N__25970),
            .I(rand_data_0));
    Odrv4 I__5563 (
            .O(N__25967),
            .I(rand_data_0));
    LocalMux I__5562 (
            .O(N__25964),
            .I(rand_data_0));
    LocalMux I__5561 (
            .O(N__25961),
            .I(rand_data_0));
    InMux I__5560 (
            .O(N__25950),
            .I(N__25938));
    InMux I__5559 (
            .O(N__25949),
            .I(N__25938));
    InMux I__5558 (
            .O(N__25948),
            .I(N__25938));
    InMux I__5557 (
            .O(N__25947),
            .I(N__25938));
    LocalMux I__5556 (
            .O(N__25938),
            .I(n9077));
    InMux I__5555 (
            .O(N__25935),
            .I(N__25929));
    InMux I__5554 (
            .O(N__25934),
            .I(N__25929));
    LocalMux I__5553 (
            .O(N__25929),
            .I(n5185));
    InMux I__5552 (
            .O(N__25926),
            .I(N__25922));
    InMux I__5551 (
            .O(N__25925),
            .I(N__25919));
    LocalMux I__5550 (
            .O(N__25922),
            .I(N__25916));
    LocalMux I__5549 (
            .O(N__25919),
            .I(N__25913));
    Span4Mux_h I__5548 (
            .O(N__25916),
            .I(N__25910));
    Span4Mux_h I__5547 (
            .O(N__25913),
            .I(N__25907));
    Span4Mux_v I__5546 (
            .O(N__25910),
            .I(N__25903));
    Span4Mux_v I__5545 (
            .O(N__25907),
            .I(N__25900));
    CascadeMux I__5544 (
            .O(N__25906),
            .I(N__25897));
    Span4Mux_v I__5543 (
            .O(N__25903),
            .I(N__25892));
    Span4Mux_v I__5542 (
            .O(N__25900),
            .I(N__25889));
    InMux I__5541 (
            .O(N__25897),
            .I(N__25882));
    InMux I__5540 (
            .O(N__25896),
            .I(N__25882));
    InMux I__5539 (
            .O(N__25895),
            .I(N__25882));
    Odrv4 I__5538 (
            .O(N__25892),
            .I(r_Bit_Index_0_adj_1733));
    Odrv4 I__5537 (
            .O(N__25889),
            .I(r_Bit_Index_0_adj_1733));
    LocalMux I__5536 (
            .O(N__25882),
            .I(r_Bit_Index_0_adj_1733));
    InMux I__5535 (
            .O(N__25875),
            .I(N__25870));
    InMux I__5534 (
            .O(N__25874),
            .I(N__25867));
    InMux I__5533 (
            .O(N__25873),
            .I(N__25864));
    LocalMux I__5532 (
            .O(N__25870),
            .I(N__25860));
    LocalMux I__5531 (
            .O(N__25867),
            .I(N__25855));
    LocalMux I__5530 (
            .O(N__25864),
            .I(N__25855));
    InMux I__5529 (
            .O(N__25863),
            .I(N__25852));
    Span4Mux_v I__5528 (
            .O(N__25860),
            .I(N__25849));
    Span12Mux_s8_h I__5527 (
            .O(N__25855),
            .I(N__25844));
    LocalMux I__5526 (
            .O(N__25852),
            .I(N__25844));
    Span4Mux_v I__5525 (
            .O(N__25849),
            .I(N__25839));
    Span12Mux_v I__5524 (
            .O(N__25844),
            .I(N__25836));
    InMux I__5523 (
            .O(N__25843),
            .I(N__25831));
    InMux I__5522 (
            .O(N__25842),
            .I(N__25831));
    Odrv4 I__5521 (
            .O(N__25839),
            .I(r_Bit_Index_1_adj_1732));
    Odrv12 I__5520 (
            .O(N__25836),
            .I(r_Bit_Index_1_adj_1732));
    LocalMux I__5519 (
            .O(N__25831),
            .I(r_Bit_Index_1_adj_1732));
    InMux I__5518 (
            .O(N__25824),
            .I(N__25818));
    InMux I__5517 (
            .O(N__25823),
            .I(N__25818));
    LocalMux I__5516 (
            .O(N__25818),
            .I(N__25815));
    Span4Mux_v I__5515 (
            .O(N__25815),
            .I(N__25812));
    Odrv4 I__5514 (
            .O(N__25812),
            .I(n4_adj_1724));
    CascadeMux I__5513 (
            .O(N__25809),
            .I(N__25805));
    InMux I__5512 (
            .O(N__25808),
            .I(N__25801));
    InMux I__5511 (
            .O(N__25805),
            .I(N__25798));
    InMux I__5510 (
            .O(N__25804),
            .I(N__25795));
    LocalMux I__5509 (
            .O(N__25801),
            .I(N__25792));
    LocalMux I__5508 (
            .O(N__25798),
            .I(N__25788));
    LocalMux I__5507 (
            .O(N__25795),
            .I(N__25785));
    Span4Mux_v I__5506 (
            .O(N__25792),
            .I(N__25781));
    InMux I__5505 (
            .O(N__25791),
            .I(N__25778));
    Span4Mux_v I__5504 (
            .O(N__25788),
            .I(N__25773));
    Span4Mux_v I__5503 (
            .O(N__25785),
            .I(N__25773));
    InMux I__5502 (
            .O(N__25784),
            .I(N__25770));
    Span4Mux_v I__5501 (
            .O(N__25781),
            .I(N__25767));
    LocalMux I__5500 (
            .O(N__25778),
            .I(N__25764));
    Span4Mux_h I__5499 (
            .O(N__25773),
            .I(N__25761));
    LocalMux I__5498 (
            .O(N__25770),
            .I(data_in_field_134));
    Odrv4 I__5497 (
            .O(N__25767),
            .I(data_in_field_134));
    Odrv12 I__5496 (
            .O(N__25764),
            .I(data_in_field_134));
    Odrv4 I__5495 (
            .O(N__25761),
            .I(data_in_field_134));
    InMux I__5494 (
            .O(N__25752),
            .I(N__25749));
    LocalMux I__5493 (
            .O(N__25749),
            .I(N__25746));
    Span4Mux_v I__5492 (
            .O(N__25746),
            .I(N__25742));
    InMux I__5491 (
            .O(N__25745),
            .I(N__25737));
    Span4Mux_h I__5490 (
            .O(N__25742),
            .I(N__25734));
    InMux I__5489 (
            .O(N__25741),
            .I(N__25729));
    InMux I__5488 (
            .O(N__25740),
            .I(N__25729));
    LocalMux I__5487 (
            .O(N__25737),
            .I(data_in_field_119));
    Odrv4 I__5486 (
            .O(N__25734),
            .I(data_in_field_119));
    LocalMux I__5485 (
            .O(N__25729),
            .I(data_in_field_119));
    InMux I__5484 (
            .O(N__25722),
            .I(N__25719));
    LocalMux I__5483 (
            .O(N__25719),
            .I(N__25715));
    InMux I__5482 (
            .O(N__25718),
            .I(N__25712));
    Span4Mux_h I__5481 (
            .O(N__25715),
            .I(N__25706));
    LocalMux I__5480 (
            .O(N__25712),
            .I(N__25706));
    InMux I__5479 (
            .O(N__25711),
            .I(N__25703));
    Span4Mux_v I__5478 (
            .O(N__25706),
            .I(N__25700));
    LocalMux I__5477 (
            .O(N__25703),
            .I(N__25697));
    Span4Mux_s3_h I__5476 (
            .O(N__25700),
            .I(N__25694));
    Span4Mux_h I__5475 (
            .O(N__25697),
            .I(N__25691));
    Odrv4 I__5474 (
            .O(N__25694),
            .I(\c0.n8883 ));
    Odrv4 I__5473 (
            .O(N__25691),
            .I(\c0.n8883 ));
    InMux I__5472 (
            .O(N__25686),
            .I(N__25683));
    LocalMux I__5471 (
            .O(N__25683),
            .I(N__25680));
    Odrv4 I__5470 (
            .O(N__25680),
            .I(\c0.n8770 ));
    InMux I__5469 (
            .O(N__25677),
            .I(N__25674));
    LocalMux I__5468 (
            .O(N__25674),
            .I(N__25670));
    CascadeMux I__5467 (
            .O(N__25673),
            .I(N__25667));
    Span4Mux_v I__5466 (
            .O(N__25670),
            .I(N__25664));
    InMux I__5465 (
            .O(N__25667),
            .I(N__25661));
    Span4Mux_h I__5464 (
            .O(N__25664),
            .I(N__25656));
    LocalMux I__5463 (
            .O(N__25661),
            .I(N__25656));
    Span4Mux_h I__5462 (
            .O(N__25656),
            .I(N__25653));
    Span4Mux_v I__5461 (
            .O(N__25653),
            .I(N__25650));
    Odrv4 I__5460 (
            .O(N__25650),
            .I(\c0.n8810 ));
    InMux I__5459 (
            .O(N__25647),
            .I(N__25644));
    LocalMux I__5458 (
            .O(N__25644),
            .I(N__25641));
    Span4Mux_v I__5457 (
            .O(N__25641),
            .I(N__25637));
    InMux I__5456 (
            .O(N__25640),
            .I(N__25634));
    Span4Mux_h I__5455 (
            .O(N__25637),
            .I(N__25629));
    LocalMux I__5454 (
            .O(N__25634),
            .I(N__25629));
    Span4Mux_h I__5453 (
            .O(N__25629),
            .I(N__25626));
    Odrv4 I__5452 (
            .O(N__25626),
            .I(\c0.n8899 ));
    InMux I__5451 (
            .O(N__25623),
            .I(N__25620));
    LocalMux I__5450 (
            .O(N__25620),
            .I(\c0.n16_adj_1657 ));
    CascadeMux I__5449 (
            .O(N__25617),
            .I(\c0.n22_adj_1655_cascade_ ));
    InMux I__5448 (
            .O(N__25614),
            .I(N__25608));
    InMux I__5447 (
            .O(N__25613),
            .I(N__25605));
    CascadeMux I__5446 (
            .O(N__25612),
            .I(N__25600));
    CascadeMux I__5445 (
            .O(N__25611),
            .I(N__25597));
    LocalMux I__5444 (
            .O(N__25608),
            .I(N__25594));
    LocalMux I__5443 (
            .O(N__25605),
            .I(N__25591));
    InMux I__5442 (
            .O(N__25604),
            .I(N__25586));
    InMux I__5441 (
            .O(N__25603),
            .I(N__25586));
    InMux I__5440 (
            .O(N__25600),
            .I(N__25581));
    InMux I__5439 (
            .O(N__25597),
            .I(N__25581));
    Odrv12 I__5438 (
            .O(N__25594),
            .I(data_in_field_37));
    Odrv4 I__5437 (
            .O(N__25591),
            .I(data_in_field_37));
    LocalMux I__5436 (
            .O(N__25586),
            .I(data_in_field_37));
    LocalMux I__5435 (
            .O(N__25581),
            .I(data_in_field_37));
    InMux I__5434 (
            .O(N__25572),
            .I(N__25569));
    LocalMux I__5433 (
            .O(N__25569),
            .I(\c0.n24_adj_1658 ));
    CascadeMux I__5432 (
            .O(N__25566),
            .I(N__25563));
    InMux I__5431 (
            .O(N__25563),
            .I(N__25560));
    LocalMux I__5430 (
            .O(N__25560),
            .I(N__25557));
    Span4Mux_h I__5429 (
            .O(N__25557),
            .I(N__25554));
    Span4Mux_h I__5428 (
            .O(N__25554),
            .I(N__25550));
    InMux I__5427 (
            .O(N__25553),
            .I(N__25547));
    Odrv4 I__5426 (
            .O(N__25550),
            .I(\c0.n8939 ));
    LocalMux I__5425 (
            .O(N__25547),
            .I(\c0.n8939 ));
    InMux I__5424 (
            .O(N__25542),
            .I(N__25539));
    LocalMux I__5423 (
            .O(N__25539),
            .I(N__25536));
    Span4Mux_v I__5422 (
            .O(N__25536),
            .I(N__25533));
    Span4Mux_h I__5421 (
            .O(N__25533),
            .I(N__25530));
    Odrv4 I__5420 (
            .O(N__25530),
            .I(\c0.n20_adj_1659 ));
    InMux I__5419 (
            .O(N__25527),
            .I(N__25524));
    LocalMux I__5418 (
            .O(N__25524),
            .I(N__25520));
    InMux I__5417 (
            .O(N__25523),
            .I(N__25517));
    Span4Mux_h I__5416 (
            .O(N__25520),
            .I(N__25514));
    LocalMux I__5415 (
            .O(N__25517),
            .I(N__25508));
    IoSpan4Mux I__5414 (
            .O(N__25514),
            .I(N__25505));
    InMux I__5413 (
            .O(N__25513),
            .I(N__25500));
    InMux I__5412 (
            .O(N__25512),
            .I(N__25500));
    InMux I__5411 (
            .O(N__25511),
            .I(N__25497));
    Span4Mux_h I__5410 (
            .O(N__25508),
            .I(N__25494));
    Sp12to4 I__5409 (
            .O(N__25505),
            .I(N__25489));
    LocalMux I__5408 (
            .O(N__25500),
            .I(N__25489));
    LocalMux I__5407 (
            .O(N__25497),
            .I(data_in_field_68));
    Odrv4 I__5406 (
            .O(N__25494),
            .I(data_in_field_68));
    Odrv12 I__5405 (
            .O(N__25489),
            .I(data_in_field_68));
    CascadeMux I__5404 (
            .O(N__25482),
            .I(N__25477));
    InMux I__5403 (
            .O(N__25481),
            .I(N__25473));
    InMux I__5402 (
            .O(N__25480),
            .I(N__25470));
    InMux I__5401 (
            .O(N__25477),
            .I(N__25467));
    InMux I__5400 (
            .O(N__25476),
            .I(N__25464));
    LocalMux I__5399 (
            .O(N__25473),
            .I(N__25461));
    LocalMux I__5398 (
            .O(N__25470),
            .I(N__25458));
    LocalMux I__5397 (
            .O(N__25467),
            .I(N__25455));
    LocalMux I__5396 (
            .O(N__25464),
            .I(N__25445));
    Span4Mux_h I__5395 (
            .O(N__25461),
            .I(N__25445));
    Span4Mux_v I__5394 (
            .O(N__25458),
            .I(N__25445));
    Span4Mux_v I__5393 (
            .O(N__25455),
            .I(N__25445));
    InMux I__5392 (
            .O(N__25454),
            .I(N__25442));
    Odrv4 I__5391 (
            .O(N__25445),
            .I(data_in_field_76));
    LocalMux I__5390 (
            .O(N__25442),
            .I(data_in_field_76));
    InMux I__5389 (
            .O(N__25437),
            .I(N__25434));
    LocalMux I__5388 (
            .O(N__25434),
            .I(N__25431));
    Odrv4 I__5387 (
            .O(N__25431),
            .I(\c0.n9566 ));
    InMux I__5386 (
            .O(N__25428),
            .I(N__25425));
    LocalMux I__5385 (
            .O(N__25425),
            .I(N__25422));
    Odrv4 I__5384 (
            .O(N__25422),
            .I(\c0.n9171 ));
    CascadeMux I__5383 (
            .O(N__25419),
            .I(\c0.n9168_cascade_ ));
    InMux I__5382 (
            .O(N__25416),
            .I(N__25413));
    LocalMux I__5381 (
            .O(N__25413),
            .I(N__25410));
    Span4Mux_s2_v I__5380 (
            .O(N__25410),
            .I(N__25407));
    Odrv4 I__5379 (
            .O(N__25407),
            .I(\c0.n9165 ));
    CascadeMux I__5378 (
            .O(N__25404),
            .I(N__25401));
    InMux I__5377 (
            .O(N__25401),
            .I(N__25398));
    LocalMux I__5376 (
            .O(N__25398),
            .I(N__25395));
    Span4Mux_h I__5375 (
            .O(N__25395),
            .I(N__25392));
    Span4Mux_h I__5374 (
            .O(N__25392),
            .I(N__25389));
    Sp12to4 I__5373 (
            .O(N__25389),
            .I(N__25386));
    Odrv12 I__5372 (
            .O(N__25386),
            .I(\c0.n9162 ));
    InMux I__5371 (
            .O(N__25383),
            .I(N__25380));
    LocalMux I__5370 (
            .O(N__25380),
            .I(\c0.n9554 ));
    InMux I__5369 (
            .O(N__25377),
            .I(N__25374));
    LocalMux I__5368 (
            .O(N__25374),
            .I(N__25371));
    Odrv4 I__5367 (
            .O(N__25371),
            .I(\c0.n22_adj_1679 ));
    CascadeMux I__5366 (
            .O(N__25368),
            .I(\c0.n9557_cascade_ ));
    InMux I__5365 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__5364 (
            .O(N__25362),
            .I(N__25359));
    Span4Mux_s1_v I__5363 (
            .O(N__25359),
            .I(N__25356));
    Span4Mux_h I__5362 (
            .O(N__25356),
            .I(N__25353));
    Odrv4 I__5361 (
            .O(N__25353),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CascadeMux I__5360 (
            .O(N__25350),
            .I(n5185_cascade_));
    InMux I__5359 (
            .O(N__25347),
            .I(N__25343));
    InMux I__5358 (
            .O(N__25346),
            .I(N__25340));
    LocalMux I__5357 (
            .O(N__25343),
            .I(N__25335));
    LocalMux I__5356 (
            .O(N__25340),
            .I(N__25331));
    InMux I__5355 (
            .O(N__25339),
            .I(N__25328));
    InMux I__5354 (
            .O(N__25338),
            .I(N__25325));
    Span4Mux_v I__5353 (
            .O(N__25335),
            .I(N__25322));
    InMux I__5352 (
            .O(N__25334),
            .I(N__25319));
    Span4Mux_h I__5351 (
            .O(N__25331),
            .I(N__25315));
    LocalMux I__5350 (
            .O(N__25328),
            .I(N__25310));
    LocalMux I__5349 (
            .O(N__25325),
            .I(N__25310));
    Span4Mux_v I__5348 (
            .O(N__25322),
            .I(N__25307));
    LocalMux I__5347 (
            .O(N__25319),
            .I(N__25304));
    InMux I__5346 (
            .O(N__25318),
            .I(N__25300));
    Span4Mux_h I__5345 (
            .O(N__25315),
            .I(N__25295));
    Span4Mux_v I__5344 (
            .O(N__25310),
            .I(N__25295));
    Sp12to4 I__5343 (
            .O(N__25307),
            .I(N__25290));
    Span12Mux_s8_v I__5342 (
            .O(N__25304),
            .I(N__25290));
    InMux I__5341 (
            .O(N__25303),
            .I(N__25287));
    LocalMux I__5340 (
            .O(N__25300),
            .I(data_in_field_150));
    Odrv4 I__5339 (
            .O(N__25295),
            .I(data_in_field_150));
    Odrv12 I__5338 (
            .O(N__25290),
            .I(data_in_field_150));
    LocalMux I__5337 (
            .O(N__25287),
            .I(data_in_field_150));
    InMux I__5336 (
            .O(N__25278),
            .I(N__25272));
    InMux I__5335 (
            .O(N__25277),
            .I(N__25269));
    InMux I__5334 (
            .O(N__25276),
            .I(N__25266));
    InMux I__5333 (
            .O(N__25275),
            .I(N__25263));
    LocalMux I__5332 (
            .O(N__25272),
            .I(N__25259));
    LocalMux I__5331 (
            .O(N__25269),
            .I(N__25256));
    LocalMux I__5330 (
            .O(N__25266),
            .I(N__25251));
    LocalMux I__5329 (
            .O(N__25263),
            .I(N__25251));
    InMux I__5328 (
            .O(N__25262),
            .I(N__25247));
    Span12Mux_s7_v I__5327 (
            .O(N__25259),
            .I(N__25244));
    Span4Mux_v I__5326 (
            .O(N__25256),
            .I(N__25241));
    Span4Mux_v I__5325 (
            .O(N__25251),
            .I(N__25238));
    InMux I__5324 (
            .O(N__25250),
            .I(N__25235));
    LocalMux I__5323 (
            .O(N__25247),
            .I(data_in_field_52));
    Odrv12 I__5322 (
            .O(N__25244),
            .I(data_in_field_52));
    Odrv4 I__5321 (
            .O(N__25241),
            .I(data_in_field_52));
    Odrv4 I__5320 (
            .O(N__25238),
            .I(data_in_field_52));
    LocalMux I__5319 (
            .O(N__25235),
            .I(data_in_field_52));
    CascadeMux I__5318 (
            .O(N__25224),
            .I(N__25221));
    InMux I__5317 (
            .O(N__25221),
            .I(N__25215));
    InMux I__5316 (
            .O(N__25220),
            .I(N__25210));
    InMux I__5315 (
            .O(N__25219),
            .I(N__25207));
    InMux I__5314 (
            .O(N__25218),
            .I(N__25204));
    LocalMux I__5313 (
            .O(N__25215),
            .I(N__25201));
    InMux I__5312 (
            .O(N__25214),
            .I(N__25198));
    InMux I__5311 (
            .O(N__25213),
            .I(N__25195));
    LocalMux I__5310 (
            .O(N__25210),
            .I(N__25190));
    LocalMux I__5309 (
            .O(N__25207),
            .I(N__25190));
    LocalMux I__5308 (
            .O(N__25204),
            .I(N__25183));
    Span4Mux_h I__5307 (
            .O(N__25201),
            .I(N__25183));
    LocalMux I__5306 (
            .O(N__25198),
            .I(N__25183));
    LocalMux I__5305 (
            .O(N__25195),
            .I(N__25180));
    Span4Mux_v I__5304 (
            .O(N__25190),
            .I(N__25177));
    Span4Mux_v I__5303 (
            .O(N__25183),
            .I(N__25174));
    Span4Mux_h I__5302 (
            .O(N__25180),
            .I(N__25171));
    Span4Mux_v I__5301 (
            .O(N__25177),
            .I(N__25167));
    Span4Mux_h I__5300 (
            .O(N__25174),
            .I(N__25161));
    Span4Mux_v I__5299 (
            .O(N__25171),
            .I(N__25161));
    InMux I__5298 (
            .O(N__25170),
            .I(N__25158));
    Span4Mux_h I__5297 (
            .O(N__25167),
            .I(N__25155));
    InMux I__5296 (
            .O(N__25166),
            .I(N__25152));
    Span4Mux_v I__5295 (
            .O(N__25161),
            .I(N__25149));
    LocalMux I__5294 (
            .O(N__25158),
            .I(data_in_field_151));
    Odrv4 I__5293 (
            .O(N__25155),
            .I(data_in_field_151));
    LocalMux I__5292 (
            .O(N__25152),
            .I(data_in_field_151));
    Odrv4 I__5291 (
            .O(N__25149),
            .I(data_in_field_151));
    InMux I__5290 (
            .O(N__25140),
            .I(N__25135));
    InMux I__5289 (
            .O(N__25139),
            .I(N__25132));
    CascadeMux I__5288 (
            .O(N__25138),
            .I(N__25129));
    LocalMux I__5287 (
            .O(N__25135),
            .I(N__25125));
    LocalMux I__5286 (
            .O(N__25132),
            .I(N__25122));
    InMux I__5285 (
            .O(N__25129),
            .I(N__25119));
    InMux I__5284 (
            .O(N__25128),
            .I(N__25115));
    Span4Mux_s2_v I__5283 (
            .O(N__25125),
            .I(N__25112));
    Span4Mux_s2_v I__5282 (
            .O(N__25122),
            .I(N__25109));
    LocalMux I__5281 (
            .O(N__25119),
            .I(N__25106));
    InMux I__5280 (
            .O(N__25118),
            .I(N__25103));
    LocalMux I__5279 (
            .O(N__25115),
            .I(N__25100));
    Span4Mux_v I__5278 (
            .O(N__25112),
            .I(N__25095));
    Span4Mux_v I__5277 (
            .O(N__25109),
            .I(N__25095));
    Span4Mux_s3_v I__5276 (
            .O(N__25106),
            .I(N__25092));
    LocalMux I__5275 (
            .O(N__25103),
            .I(data_in_field_86));
    Odrv12 I__5274 (
            .O(N__25100),
            .I(data_in_field_86));
    Odrv4 I__5273 (
            .O(N__25095),
            .I(data_in_field_86));
    Odrv4 I__5272 (
            .O(N__25092),
            .I(data_in_field_86));
    InMux I__5271 (
            .O(N__25083),
            .I(N__25080));
    LocalMux I__5270 (
            .O(N__25080),
            .I(N__25076));
    CascadeMux I__5269 (
            .O(N__25079),
            .I(N__25073));
    Span4Mux_h I__5268 (
            .O(N__25076),
            .I(N__25070));
    InMux I__5267 (
            .O(N__25073),
            .I(N__25067));
    Span4Mux_h I__5266 (
            .O(N__25070),
            .I(N__25062));
    LocalMux I__5265 (
            .O(N__25067),
            .I(N__25062));
    Odrv4 I__5264 (
            .O(N__25062),
            .I(\c0.n8915 ));
    InMux I__5263 (
            .O(N__25059),
            .I(N__25056));
    LocalMux I__5262 (
            .O(N__25056),
            .I(N__25053));
    Span4Mux_v I__5261 (
            .O(N__25053),
            .I(N__25050));
    Span4Mux_h I__5260 (
            .O(N__25050),
            .I(N__25047));
    Odrv4 I__5259 (
            .O(N__25047),
            .I(\c0.n8788 ));
    CascadeMux I__5258 (
            .O(N__25044),
            .I(N__25041));
    InMux I__5257 (
            .O(N__25041),
            .I(N__25038));
    LocalMux I__5256 (
            .O(N__25038),
            .I(N__25035));
    Span4Mux_v I__5255 (
            .O(N__25035),
            .I(N__25031));
    InMux I__5254 (
            .O(N__25034),
            .I(N__25028));
    Odrv4 I__5253 (
            .O(N__25031),
            .I(\c0.n8828 ));
    LocalMux I__5252 (
            .O(N__25028),
            .I(\c0.n8828 ));
    InMux I__5251 (
            .O(N__25023),
            .I(N__25020));
    LocalMux I__5250 (
            .O(N__25020),
            .I(N__25016));
    InMux I__5249 (
            .O(N__25019),
            .I(N__25013));
    Span4Mux_v I__5248 (
            .O(N__25016),
            .I(N__25010));
    LocalMux I__5247 (
            .O(N__25013),
            .I(N__25007));
    Span4Mux_h I__5246 (
            .O(N__25010),
            .I(N__25002));
    Span4Mux_v I__5245 (
            .O(N__25007),
            .I(N__25002));
    Odrv4 I__5244 (
            .O(N__25002),
            .I(\c0.n8855 ));
    InMux I__5243 (
            .O(N__24999),
            .I(N__24996));
    LocalMux I__5242 (
            .O(N__24996),
            .I(N__24993));
    Span12Mux_s3_v I__5241 (
            .O(N__24993),
            .I(N__24990));
    Odrv12 I__5240 (
            .O(N__24990),
            .I(\c0.n35 ));
    CascadeMux I__5239 (
            .O(N__24987),
            .I(N__24981));
    InMux I__5238 (
            .O(N__24986),
            .I(N__24975));
    InMux I__5237 (
            .O(N__24985),
            .I(N__24975));
    InMux I__5236 (
            .O(N__24984),
            .I(N__24970));
    InMux I__5235 (
            .O(N__24981),
            .I(N__24970));
    InMux I__5234 (
            .O(N__24980),
            .I(N__24967));
    LocalMux I__5233 (
            .O(N__24975),
            .I(data_in_field_84));
    LocalMux I__5232 (
            .O(N__24970),
            .I(data_in_field_84));
    LocalMux I__5231 (
            .O(N__24967),
            .I(data_in_field_84));
    CascadeMux I__5230 (
            .O(N__24960),
            .I(N__24955));
    InMux I__5229 (
            .O(N__24959),
            .I(N__24952));
    InMux I__5228 (
            .O(N__24958),
            .I(N__24949));
    InMux I__5227 (
            .O(N__24955),
            .I(N__24945));
    LocalMux I__5226 (
            .O(N__24952),
            .I(N__24938));
    LocalMux I__5225 (
            .O(N__24949),
            .I(N__24938));
    InMux I__5224 (
            .O(N__24948),
            .I(N__24935));
    LocalMux I__5223 (
            .O(N__24945),
            .I(N__24932));
    InMux I__5222 (
            .O(N__24944),
            .I(N__24929));
    InMux I__5221 (
            .O(N__24943),
            .I(N__24926));
    Span4Mux_h I__5220 (
            .O(N__24938),
            .I(N__24923));
    LocalMux I__5219 (
            .O(N__24935),
            .I(N__24918));
    Span4Mux_h I__5218 (
            .O(N__24932),
            .I(N__24918));
    LocalMux I__5217 (
            .O(N__24929),
            .I(data_in_field_92));
    LocalMux I__5216 (
            .O(N__24926),
            .I(data_in_field_92));
    Odrv4 I__5215 (
            .O(N__24923),
            .I(data_in_field_92));
    Odrv4 I__5214 (
            .O(N__24918),
            .I(data_in_field_92));
    InMux I__5213 (
            .O(N__24909),
            .I(N__24906));
    LocalMux I__5212 (
            .O(N__24906),
            .I(\c0.n9560 ));
    InMux I__5211 (
            .O(N__24903),
            .I(N__24899));
    InMux I__5210 (
            .O(N__24902),
            .I(N__24896));
    LocalMux I__5209 (
            .O(N__24899),
            .I(N__24893));
    LocalMux I__5208 (
            .O(N__24896),
            .I(N__24890));
    Span4Mux_h I__5207 (
            .O(N__24893),
            .I(N__24882));
    Span4Mux_h I__5206 (
            .O(N__24890),
            .I(N__24882));
    InMux I__5205 (
            .O(N__24889),
            .I(N__24877));
    InMux I__5204 (
            .O(N__24888),
            .I(N__24877));
    InMux I__5203 (
            .O(N__24887),
            .I(N__24874));
    Span4Mux_v I__5202 (
            .O(N__24882),
            .I(N__24871));
    LocalMux I__5201 (
            .O(N__24877),
            .I(N__24868));
    LocalMux I__5200 (
            .O(N__24874),
            .I(data_in_field_108));
    Odrv4 I__5199 (
            .O(N__24871),
            .I(data_in_field_108));
    Odrv12 I__5198 (
            .O(N__24868),
            .I(data_in_field_108));
    InMux I__5197 (
            .O(N__24861),
            .I(N__24857));
    InMux I__5196 (
            .O(N__24860),
            .I(N__24853));
    LocalMux I__5195 (
            .O(N__24857),
            .I(N__24850));
    InMux I__5194 (
            .O(N__24856),
            .I(N__24847));
    LocalMux I__5193 (
            .O(N__24853),
            .I(N__24842));
    Span4Mux_v I__5192 (
            .O(N__24850),
            .I(N__24839));
    LocalMux I__5191 (
            .O(N__24847),
            .I(N__24836));
    InMux I__5190 (
            .O(N__24846),
            .I(N__24833));
    InMux I__5189 (
            .O(N__24845),
            .I(N__24830));
    Span4Mux_v I__5188 (
            .O(N__24842),
            .I(N__24827));
    Span4Mux_h I__5187 (
            .O(N__24839),
            .I(N__24820));
    Span4Mux_v I__5186 (
            .O(N__24836),
            .I(N__24820));
    LocalMux I__5185 (
            .O(N__24833),
            .I(N__24820));
    LocalMux I__5184 (
            .O(N__24830),
            .I(data_in_field_100));
    Odrv4 I__5183 (
            .O(N__24827),
            .I(data_in_field_100));
    Odrv4 I__5182 (
            .O(N__24820),
            .I(data_in_field_100));
    InMux I__5181 (
            .O(N__24813),
            .I(N__24810));
    LocalMux I__5180 (
            .O(N__24810),
            .I(N__24807));
    Span12Mux_h I__5179 (
            .O(N__24807),
            .I(N__24804));
    Odrv12 I__5178 (
            .O(N__24804),
            .I(\c0.n8927 ));
    InMux I__5177 (
            .O(N__24801),
            .I(N__24795));
    InMux I__5176 (
            .O(N__24800),
            .I(N__24795));
    LocalMux I__5175 (
            .O(N__24795),
            .I(N__24792));
    Odrv12 I__5174 (
            .O(N__24792),
            .I(\c0.n8837 ));
    InMux I__5173 (
            .O(N__24789),
            .I(N__24786));
    LocalMux I__5172 (
            .O(N__24786),
            .I(N__24782));
    InMux I__5171 (
            .O(N__24785),
            .I(N__24777));
    Span4Mux_v I__5170 (
            .O(N__24782),
            .I(N__24773));
    InMux I__5169 (
            .O(N__24781),
            .I(N__24770));
    InMux I__5168 (
            .O(N__24780),
            .I(N__24767));
    LocalMux I__5167 (
            .O(N__24777),
            .I(N__24764));
    InMux I__5166 (
            .O(N__24776),
            .I(N__24761));
    Span4Mux_h I__5165 (
            .O(N__24773),
            .I(N__24756));
    LocalMux I__5164 (
            .O(N__24770),
            .I(N__24756));
    LocalMux I__5163 (
            .O(N__24767),
            .I(N__24751));
    Span4Mux_h I__5162 (
            .O(N__24764),
            .I(N__24748));
    LocalMux I__5161 (
            .O(N__24761),
            .I(N__24743));
    Span4Mux_v I__5160 (
            .O(N__24756),
            .I(N__24743));
    InMux I__5159 (
            .O(N__24755),
            .I(N__24738));
    InMux I__5158 (
            .O(N__24754),
            .I(N__24738));
    Odrv12 I__5157 (
            .O(N__24751),
            .I(data_in_field_41));
    Odrv4 I__5156 (
            .O(N__24748),
            .I(data_in_field_41));
    Odrv4 I__5155 (
            .O(N__24743),
            .I(data_in_field_41));
    LocalMux I__5154 (
            .O(N__24738),
            .I(data_in_field_41));
    InMux I__5153 (
            .O(N__24729),
            .I(N__24726));
    LocalMux I__5152 (
            .O(N__24726),
            .I(N__24723));
    Odrv4 I__5151 (
            .O(N__24723),
            .I(\c0.n16_adj_1629 ));
    CascadeMux I__5150 (
            .O(N__24720),
            .I(N__24717));
    InMux I__5149 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__5148 (
            .O(N__24714),
            .I(N__24710));
    InMux I__5147 (
            .O(N__24713),
            .I(N__24707));
    Span4Mux_v I__5146 (
            .O(N__24710),
            .I(N__24704));
    LocalMux I__5145 (
            .O(N__24707),
            .I(N__24701));
    Span4Mux_h I__5144 (
            .O(N__24704),
            .I(N__24698));
    Span4Mux_s3_v I__5143 (
            .O(N__24701),
            .I(N__24695));
    Odrv4 I__5142 (
            .O(N__24698),
            .I(\c0.n8977 ));
    Odrv4 I__5141 (
            .O(N__24695),
            .I(\c0.n8977 ));
    InMux I__5140 (
            .O(N__24690),
            .I(N__24687));
    LocalMux I__5139 (
            .O(N__24687),
            .I(\c0.n17_adj_1630 ));
    CascadeMux I__5138 (
            .O(N__24684),
            .I(N__24681));
    InMux I__5137 (
            .O(N__24681),
            .I(N__24678));
    LocalMux I__5136 (
            .O(N__24678),
            .I(\c0.data_in_frame_19_4 ));
    CascadeMux I__5135 (
            .O(N__24675),
            .I(N__24672));
    InMux I__5134 (
            .O(N__24672),
            .I(N__24669));
    LocalMux I__5133 (
            .O(N__24669),
            .I(N__24666));
    Span4Mux_s3_v I__5132 (
            .O(N__24666),
            .I(N__24663));
    Span4Mux_h I__5131 (
            .O(N__24663),
            .I(N__24660));
    Odrv4 I__5130 (
            .O(N__24660),
            .I(\c0.data_in_frame_20_4 ));
    InMux I__5129 (
            .O(N__24657),
            .I(N__24651));
    InMux I__5128 (
            .O(N__24656),
            .I(N__24648));
    InMux I__5127 (
            .O(N__24655),
            .I(N__24645));
    InMux I__5126 (
            .O(N__24654),
            .I(N__24642));
    LocalMux I__5125 (
            .O(N__24651),
            .I(N__24639));
    LocalMux I__5124 (
            .O(N__24648),
            .I(N__24636));
    LocalMux I__5123 (
            .O(N__24645),
            .I(N__24633));
    LocalMux I__5122 (
            .O(N__24642),
            .I(N__24630));
    Span4Mux_v I__5121 (
            .O(N__24639),
            .I(N__24626));
    Span4Mux_h I__5120 (
            .O(N__24636),
            .I(N__24623));
    Span4Mux_v I__5119 (
            .O(N__24633),
            .I(N__24618));
    Span4Mux_h I__5118 (
            .O(N__24630),
            .I(N__24618));
    InMux I__5117 (
            .O(N__24629),
            .I(N__24615));
    Odrv4 I__5116 (
            .O(N__24626),
            .I(rand_data_6));
    Odrv4 I__5115 (
            .O(N__24623),
            .I(rand_data_6));
    Odrv4 I__5114 (
            .O(N__24618),
            .I(rand_data_6));
    LocalMux I__5113 (
            .O(N__24615),
            .I(rand_data_6));
    InMux I__5112 (
            .O(N__24606),
            .I(N__24601));
    InMux I__5111 (
            .O(N__24605),
            .I(N__24598));
    InMux I__5110 (
            .O(N__24604),
            .I(N__24595));
    LocalMux I__5109 (
            .O(N__24601),
            .I(N__24590));
    LocalMux I__5108 (
            .O(N__24598),
            .I(N__24590));
    LocalMux I__5107 (
            .O(N__24595),
            .I(N__24587));
    Span4Mux_h I__5106 (
            .O(N__24590),
            .I(N__24584));
    Span4Mux_s1_v I__5105 (
            .O(N__24587),
            .I(N__24581));
    Span4Mux_h I__5104 (
            .O(N__24584),
            .I(N__24576));
    Span4Mux_v I__5103 (
            .O(N__24581),
            .I(N__24573));
    InMux I__5102 (
            .O(N__24580),
            .I(N__24568));
    InMux I__5101 (
            .O(N__24579),
            .I(N__24568));
    Odrv4 I__5100 (
            .O(N__24576),
            .I(data_in_field_102));
    Odrv4 I__5099 (
            .O(N__24573),
            .I(data_in_field_102));
    LocalMux I__5098 (
            .O(N__24568),
            .I(data_in_field_102));
    InMux I__5097 (
            .O(N__24561),
            .I(N__24556));
    InMux I__5096 (
            .O(N__24560),
            .I(N__24553));
    CascadeMux I__5095 (
            .O(N__24559),
            .I(N__24550));
    LocalMux I__5094 (
            .O(N__24556),
            .I(N__24546));
    LocalMux I__5093 (
            .O(N__24553),
            .I(N__24543));
    InMux I__5092 (
            .O(N__24550),
            .I(N__24540));
    InMux I__5091 (
            .O(N__24549),
            .I(N__24536));
    Span4Mux_v I__5090 (
            .O(N__24546),
            .I(N__24533));
    Span4Mux_s2_h I__5089 (
            .O(N__24543),
            .I(N__24530));
    LocalMux I__5088 (
            .O(N__24540),
            .I(N__24527));
    InMux I__5087 (
            .O(N__24539),
            .I(N__24524));
    LocalMux I__5086 (
            .O(N__24536),
            .I(N__24521));
    Span4Mux_h I__5085 (
            .O(N__24533),
            .I(N__24518));
    Span4Mux_h I__5084 (
            .O(N__24530),
            .I(N__24513));
    Span4Mux_s2_v I__5083 (
            .O(N__24527),
            .I(N__24513));
    LocalMux I__5082 (
            .O(N__24524),
            .I(data_in_field_125));
    Odrv4 I__5081 (
            .O(N__24521),
            .I(data_in_field_125));
    Odrv4 I__5080 (
            .O(N__24518),
            .I(data_in_field_125));
    Odrv4 I__5079 (
            .O(N__24513),
            .I(data_in_field_125));
    InMux I__5078 (
            .O(N__24504),
            .I(N__24500));
    CascadeMux I__5077 (
            .O(N__24503),
            .I(N__24497));
    LocalMux I__5076 (
            .O(N__24500),
            .I(N__24494));
    InMux I__5075 (
            .O(N__24497),
            .I(N__24491));
    Span4Mux_v I__5074 (
            .O(N__24494),
            .I(N__24485));
    LocalMux I__5073 (
            .O(N__24491),
            .I(N__24482));
    InMux I__5072 (
            .O(N__24490),
            .I(N__24479));
    InMux I__5071 (
            .O(N__24489),
            .I(N__24476));
    InMux I__5070 (
            .O(N__24488),
            .I(N__24473));
    Span4Mux_h I__5069 (
            .O(N__24485),
            .I(N__24466));
    Span4Mux_v I__5068 (
            .O(N__24482),
            .I(N__24466));
    LocalMux I__5067 (
            .O(N__24479),
            .I(N__24466));
    LocalMux I__5066 (
            .O(N__24476),
            .I(data_in_field_73));
    LocalMux I__5065 (
            .O(N__24473),
            .I(data_in_field_73));
    Odrv4 I__5064 (
            .O(N__24466),
            .I(data_in_field_73));
    CascadeMux I__5063 (
            .O(N__24459),
            .I(N__24456));
    InMux I__5062 (
            .O(N__24456),
            .I(N__24453));
    LocalMux I__5061 (
            .O(N__24453),
            .I(\c0.n18_adj_1618 ));
    InMux I__5060 (
            .O(N__24450),
            .I(N__24446));
    InMux I__5059 (
            .O(N__24449),
            .I(N__24443));
    LocalMux I__5058 (
            .O(N__24446),
            .I(N__24438));
    LocalMux I__5057 (
            .O(N__24443),
            .I(N__24434));
    InMux I__5056 (
            .O(N__24442),
            .I(N__24429));
    InMux I__5055 (
            .O(N__24441),
            .I(N__24429));
    Span4Mux_h I__5054 (
            .O(N__24438),
            .I(N__24426));
    InMux I__5053 (
            .O(N__24437),
            .I(N__24423));
    Span4Mux_h I__5052 (
            .O(N__24434),
            .I(N__24420));
    LocalMux I__5051 (
            .O(N__24429),
            .I(N__24417));
    Span4Mux_v I__5050 (
            .O(N__24426),
            .I(N__24414));
    LocalMux I__5049 (
            .O(N__24423),
            .I(N__24407));
    Span4Mux_v I__5048 (
            .O(N__24420),
            .I(N__24407));
    Span4Mux_v I__5047 (
            .O(N__24417),
            .I(N__24407));
    Odrv4 I__5046 (
            .O(N__24414),
            .I(data_in_field_54));
    Odrv4 I__5045 (
            .O(N__24407),
            .I(data_in_field_54));
    InMux I__5044 (
            .O(N__24402),
            .I(N__24399));
    LocalMux I__5043 (
            .O(N__24399),
            .I(N__24395));
    InMux I__5042 (
            .O(N__24398),
            .I(N__24392));
    Span4Mux_h I__5041 (
            .O(N__24395),
            .I(N__24387));
    LocalMux I__5040 (
            .O(N__24392),
            .I(N__24384));
    InMux I__5039 (
            .O(N__24391),
            .I(N__24379));
    InMux I__5038 (
            .O(N__24390),
            .I(N__24379));
    Odrv4 I__5037 (
            .O(N__24387),
            .I(data_in_field_69));
    Odrv4 I__5036 (
            .O(N__24384),
            .I(data_in_field_69));
    LocalMux I__5035 (
            .O(N__24379),
            .I(data_in_field_69));
    InMux I__5034 (
            .O(N__24372),
            .I(N__24369));
    LocalMux I__5033 (
            .O(N__24369),
            .I(N__24366));
    Span4Mux_v I__5032 (
            .O(N__24366),
            .I(N__24362));
    InMux I__5031 (
            .O(N__24365),
            .I(N__24359));
    Span4Mux_h I__5030 (
            .O(N__24362),
            .I(N__24354));
    LocalMux I__5029 (
            .O(N__24359),
            .I(N__24354));
    Odrv4 I__5028 (
            .O(N__24354),
            .I(\c0.n8998 ));
    InMux I__5027 (
            .O(N__24351),
            .I(N__24348));
    LocalMux I__5026 (
            .O(N__24348),
            .I(N__24345));
    Span4Mux_s3_h I__5025 (
            .O(N__24345),
            .I(N__24342));
    Span4Mux_h I__5024 (
            .O(N__24342),
            .I(N__24339));
    Odrv4 I__5023 (
            .O(N__24339),
            .I(\c0.n16_adj_1591 ));
    InMux I__5022 (
            .O(N__24336),
            .I(N__24333));
    LocalMux I__5021 (
            .O(N__24333),
            .I(N__24328));
    InMux I__5020 (
            .O(N__24332),
            .I(N__24323));
    InMux I__5019 (
            .O(N__24331),
            .I(N__24323));
    Span4Mux_v I__5018 (
            .O(N__24328),
            .I(N__24320));
    LocalMux I__5017 (
            .O(N__24323),
            .I(N__24317));
    Span4Mux_v I__5016 (
            .O(N__24320),
            .I(N__24314));
    Span4Mux_v I__5015 (
            .O(N__24317),
            .I(N__24308));
    Span4Mux_h I__5014 (
            .O(N__24314),
            .I(N__24308));
    InMux I__5013 (
            .O(N__24313),
            .I(N__24305));
    Odrv4 I__5012 (
            .O(N__24308),
            .I(rand_data_20));
    LocalMux I__5011 (
            .O(N__24305),
            .I(rand_data_20));
    InMux I__5010 (
            .O(N__24300),
            .I(N__24293));
    InMux I__5009 (
            .O(N__24299),
            .I(N__24293));
    InMux I__5008 (
            .O(N__24298),
            .I(N__24288));
    LocalMux I__5007 (
            .O(N__24293),
            .I(N__24285));
    InMux I__5006 (
            .O(N__24292),
            .I(N__24282));
    InMux I__5005 (
            .O(N__24291),
            .I(N__24278));
    LocalMux I__5004 (
            .O(N__24288),
            .I(N__24273));
    Span4Mux_h I__5003 (
            .O(N__24285),
            .I(N__24273));
    LocalMux I__5002 (
            .O(N__24282),
            .I(N__24270));
    InMux I__5001 (
            .O(N__24281),
            .I(N__24267));
    LocalMux I__5000 (
            .O(N__24278),
            .I(N__24264));
    Span4Mux_v I__4999 (
            .O(N__24273),
            .I(N__24261));
    Span4Mux_h I__4998 (
            .O(N__24270),
            .I(N__24258));
    LocalMux I__4997 (
            .O(N__24267),
            .I(data_in_field_124));
    Odrv4 I__4996 (
            .O(N__24264),
            .I(data_in_field_124));
    Odrv4 I__4995 (
            .O(N__24261),
            .I(data_in_field_124));
    Odrv4 I__4994 (
            .O(N__24258),
            .I(data_in_field_124));
    InMux I__4993 (
            .O(N__24249),
            .I(N__24246));
    LocalMux I__4992 (
            .O(N__24246),
            .I(N__24243));
    Span4Mux_h I__4991 (
            .O(N__24243),
            .I(N__24237));
    InMux I__4990 (
            .O(N__24242),
            .I(N__24230));
    InMux I__4989 (
            .O(N__24241),
            .I(N__24230));
    InMux I__4988 (
            .O(N__24240),
            .I(N__24230));
    Odrv4 I__4987 (
            .O(N__24237),
            .I(data_in_field_116));
    LocalMux I__4986 (
            .O(N__24230),
            .I(data_in_field_116));
    InMux I__4985 (
            .O(N__24225),
            .I(N__24220));
    InMux I__4984 (
            .O(N__24224),
            .I(N__24217));
    InMux I__4983 (
            .O(N__24223),
            .I(N__24214));
    LocalMux I__4982 (
            .O(N__24220),
            .I(N__24208));
    LocalMux I__4981 (
            .O(N__24217),
            .I(N__24208));
    LocalMux I__4980 (
            .O(N__24214),
            .I(N__24205));
    InMux I__4979 (
            .O(N__24213),
            .I(N__24202));
    Span4Mux_v I__4978 (
            .O(N__24208),
            .I(N__24199));
    Span4Mux_v I__4977 (
            .O(N__24205),
            .I(N__24196));
    LocalMux I__4976 (
            .O(N__24202),
            .I(data_in_field_56));
    Odrv4 I__4975 (
            .O(N__24199),
            .I(data_in_field_56));
    Odrv4 I__4974 (
            .O(N__24196),
            .I(data_in_field_56));
    CascadeMux I__4973 (
            .O(N__24189),
            .I(N__24185));
    InMux I__4972 (
            .O(N__24188),
            .I(N__24180));
    InMux I__4971 (
            .O(N__24185),
            .I(N__24177));
    InMux I__4970 (
            .O(N__24184),
            .I(N__24174));
    InMux I__4969 (
            .O(N__24183),
            .I(N__24171));
    LocalMux I__4968 (
            .O(N__24180),
            .I(N__24168));
    LocalMux I__4967 (
            .O(N__24177),
            .I(N__24165));
    LocalMux I__4966 (
            .O(N__24174),
            .I(N__24162));
    LocalMux I__4965 (
            .O(N__24171),
            .I(N__24159));
    Span4Mux_s2_v I__4964 (
            .O(N__24168),
            .I(N__24155));
    Span4Mux_v I__4963 (
            .O(N__24165),
            .I(N__24150));
    Span4Mux_v I__4962 (
            .O(N__24162),
            .I(N__24150));
    Span4Mux_h I__4961 (
            .O(N__24159),
            .I(N__24147));
    InMux I__4960 (
            .O(N__24158),
            .I(N__24144));
    Span4Mux_h I__4959 (
            .O(N__24155),
            .I(N__24141));
    Span4Mux_h I__4958 (
            .O(N__24150),
            .I(N__24136));
    Span4Mux_v I__4957 (
            .O(N__24147),
            .I(N__24136));
    LocalMux I__4956 (
            .O(N__24144),
            .I(data_in_field_101));
    Odrv4 I__4955 (
            .O(N__24141),
            .I(data_in_field_101));
    Odrv4 I__4954 (
            .O(N__24136),
            .I(data_in_field_101));
    InMux I__4953 (
            .O(N__24129),
            .I(N__24124));
    InMux I__4952 (
            .O(N__24128),
            .I(N__24121));
    InMux I__4951 (
            .O(N__24127),
            .I(N__24118));
    LocalMux I__4950 (
            .O(N__24124),
            .I(N__24113));
    LocalMux I__4949 (
            .O(N__24121),
            .I(N__24113));
    LocalMux I__4948 (
            .O(N__24118),
            .I(N__24110));
    Span4Mux_v I__4947 (
            .O(N__24113),
            .I(N__24107));
    Span4Mux_v I__4946 (
            .O(N__24110),
            .I(N__24103));
    Span4Mux_h I__4945 (
            .O(N__24107),
            .I(N__24100));
    InMux I__4944 (
            .O(N__24106),
            .I(N__24097));
    Odrv4 I__4943 (
            .O(N__24103),
            .I(rand_data_16));
    Odrv4 I__4942 (
            .O(N__24100),
            .I(rand_data_16));
    LocalMux I__4941 (
            .O(N__24097),
            .I(rand_data_16));
    InMux I__4940 (
            .O(N__24090),
            .I(N__24086));
    InMux I__4939 (
            .O(N__24089),
            .I(N__24083));
    LocalMux I__4938 (
            .O(N__24086),
            .I(N__24077));
    LocalMux I__4937 (
            .O(N__24083),
            .I(N__24077));
    InMux I__4936 (
            .O(N__24082),
            .I(N__24074));
    Span4Mux_v I__4935 (
            .O(N__24077),
            .I(N__24071));
    LocalMux I__4934 (
            .O(N__24074),
            .I(N__24067));
    Span4Mux_v I__4933 (
            .O(N__24071),
            .I(N__24064));
    InMux I__4932 (
            .O(N__24070),
            .I(N__24061));
    Span12Mux_h I__4931 (
            .O(N__24067),
            .I(N__24058));
    Span4Mux_s2_v I__4930 (
            .O(N__24064),
            .I(N__24055));
    LocalMux I__4929 (
            .O(N__24061),
            .I(rand_data_26));
    Odrv12 I__4928 (
            .O(N__24058),
            .I(rand_data_26));
    Odrv4 I__4927 (
            .O(N__24055),
            .I(rand_data_26));
    InMux I__4926 (
            .O(N__24048),
            .I(N__24044));
    InMux I__4925 (
            .O(N__24047),
            .I(N__24041));
    LocalMux I__4924 (
            .O(N__24044),
            .I(N__24037));
    LocalMux I__4923 (
            .O(N__24041),
            .I(N__24034));
    InMux I__4922 (
            .O(N__24040),
            .I(N__24030));
    Span4Mux_v I__4921 (
            .O(N__24037),
            .I(N__24027));
    Sp12to4 I__4920 (
            .O(N__24034),
            .I(N__24024));
    InMux I__4919 (
            .O(N__24033),
            .I(N__24021));
    LocalMux I__4918 (
            .O(N__24030),
            .I(data_in_field_58));
    Odrv4 I__4917 (
            .O(N__24027),
            .I(data_in_field_58));
    Odrv12 I__4916 (
            .O(N__24024),
            .I(data_in_field_58));
    LocalMux I__4915 (
            .O(N__24021),
            .I(data_in_field_58));
    InMux I__4914 (
            .O(N__24012),
            .I(N__24007));
    InMux I__4913 (
            .O(N__24011),
            .I(N__24004));
    CascadeMux I__4912 (
            .O(N__24010),
            .I(N__24000));
    LocalMux I__4911 (
            .O(N__24007),
            .I(N__23997));
    LocalMux I__4910 (
            .O(N__24004),
            .I(N__23994));
    InMux I__4909 (
            .O(N__24003),
            .I(N__23991));
    InMux I__4908 (
            .O(N__24000),
            .I(N__23988));
    Span4Mux_h I__4907 (
            .O(N__23997),
            .I(N__23985));
    Span12Mux_s1_v I__4906 (
            .O(N__23994),
            .I(N__23980));
    LocalMux I__4905 (
            .O(N__23991),
            .I(N__23980));
    LocalMux I__4904 (
            .O(N__23988),
            .I(data_in_field_118));
    Odrv4 I__4903 (
            .O(N__23985),
            .I(data_in_field_118));
    Odrv12 I__4902 (
            .O(N__23980),
            .I(data_in_field_118));
    CascadeMux I__4901 (
            .O(N__23973),
            .I(N__23970));
    InMux I__4900 (
            .O(N__23970),
            .I(N__23967));
    LocalMux I__4899 (
            .O(N__23967),
            .I(\c0.n4534 ));
    InMux I__4898 (
            .O(N__23964),
            .I(N__23961));
    LocalMux I__4897 (
            .O(N__23961),
            .I(N__23958));
    Span4Mux_h I__4896 (
            .O(N__23958),
            .I(N__23955));
    Odrv4 I__4895 (
            .O(N__23955),
            .I(\c0.n27_adj_1621 ));
    InMux I__4894 (
            .O(N__23952),
            .I(N__23948));
    InMux I__4893 (
            .O(N__23951),
            .I(N__23945));
    LocalMux I__4892 (
            .O(N__23948),
            .I(N__23938));
    LocalMux I__4891 (
            .O(N__23945),
            .I(N__23938));
    InMux I__4890 (
            .O(N__23944),
            .I(N__23933));
    InMux I__4889 (
            .O(N__23943),
            .I(N__23933));
    Span12Mux_h I__4888 (
            .O(N__23938),
            .I(N__23929));
    LocalMux I__4887 (
            .O(N__23933),
            .I(N__23926));
    InMux I__4886 (
            .O(N__23932),
            .I(N__23923));
    Odrv12 I__4885 (
            .O(N__23929),
            .I(rand_data_10));
    Odrv4 I__4884 (
            .O(N__23926),
            .I(rand_data_10));
    LocalMux I__4883 (
            .O(N__23923),
            .I(rand_data_10));
    CascadeMux I__4882 (
            .O(N__23916),
            .I(N__23913));
    InMux I__4881 (
            .O(N__23913),
            .I(N__23910));
    LocalMux I__4880 (
            .O(N__23910),
            .I(N__23907));
    Span12Mux_s5_v I__4879 (
            .O(N__23907),
            .I(N__23904));
    Odrv12 I__4878 (
            .O(N__23904),
            .I(\c0.n4473 ));
    CascadeMux I__4877 (
            .O(N__23901),
            .I(\c0.n4473_cascade_ ));
    InMux I__4876 (
            .O(N__23898),
            .I(N__23895));
    LocalMux I__4875 (
            .O(N__23895),
            .I(N__23891));
    InMux I__4874 (
            .O(N__23894),
            .I(N__23888));
    Span4Mux_h I__4873 (
            .O(N__23891),
            .I(N__23885));
    LocalMux I__4872 (
            .O(N__23888),
            .I(\c0.n9010 ));
    Odrv4 I__4871 (
            .O(N__23885),
            .I(\c0.n9010 ));
    CascadeMux I__4870 (
            .O(N__23880),
            .I(\c0.n4244_cascade_ ));
    InMux I__4869 (
            .O(N__23877),
            .I(N__23874));
    LocalMux I__4868 (
            .O(N__23874),
            .I(N__23871));
    Span4Mux_v I__4867 (
            .O(N__23871),
            .I(N__23868));
    Span4Mux_h I__4866 (
            .O(N__23868),
            .I(N__23865));
    Odrv4 I__4865 (
            .O(N__23865),
            .I(\c0.n4479 ));
    CascadeMux I__4864 (
            .O(N__23862),
            .I(\c0.n4235_cascade_ ));
    InMux I__4863 (
            .O(N__23859),
            .I(N__23856));
    LocalMux I__4862 (
            .O(N__23856),
            .I(\c0.n4562 ));
    CascadeMux I__4861 (
            .O(N__23853),
            .I(N__23846));
    InMux I__4860 (
            .O(N__23852),
            .I(N__23842));
    InMux I__4859 (
            .O(N__23851),
            .I(N__23839));
    InMux I__4858 (
            .O(N__23850),
            .I(N__23834));
    InMux I__4857 (
            .O(N__23849),
            .I(N__23834));
    InMux I__4856 (
            .O(N__23846),
            .I(N__23831));
    InMux I__4855 (
            .O(N__23845),
            .I(N__23828));
    LocalMux I__4854 (
            .O(N__23842),
            .I(N__23825));
    LocalMux I__4853 (
            .O(N__23839),
            .I(N__23821));
    LocalMux I__4852 (
            .O(N__23834),
            .I(N__23818));
    LocalMux I__4851 (
            .O(N__23831),
            .I(N__23815));
    LocalMux I__4850 (
            .O(N__23828),
            .I(N__23810));
    Span4Mux_s3_h I__4849 (
            .O(N__23825),
            .I(N__23810));
    InMux I__4848 (
            .O(N__23824),
            .I(N__23807));
    Span4Mux_h I__4847 (
            .O(N__23821),
            .I(N__23804));
    Span4Mux_h I__4846 (
            .O(N__23818),
            .I(N__23799));
    Span4Mux_h I__4845 (
            .O(N__23815),
            .I(N__23799));
    Span4Mux_v I__4844 (
            .O(N__23810),
            .I(N__23796));
    LocalMux I__4843 (
            .O(N__23807),
            .I(data_in_field_99));
    Odrv4 I__4842 (
            .O(N__23804),
            .I(data_in_field_99));
    Odrv4 I__4841 (
            .O(N__23799),
            .I(data_in_field_99));
    Odrv4 I__4840 (
            .O(N__23796),
            .I(data_in_field_99));
    CascadeMux I__4839 (
            .O(N__23787),
            .I(N__23783));
    InMux I__4838 (
            .O(N__23786),
            .I(N__23776));
    InMux I__4837 (
            .O(N__23783),
            .I(N__23776));
    InMux I__4836 (
            .O(N__23782),
            .I(N__23772));
    InMux I__4835 (
            .O(N__23781),
            .I(N__23769));
    LocalMux I__4834 (
            .O(N__23776),
            .I(N__23766));
    CascadeMux I__4833 (
            .O(N__23775),
            .I(N__23763));
    LocalMux I__4832 (
            .O(N__23772),
            .I(N__23759));
    LocalMux I__4831 (
            .O(N__23769),
            .I(N__23756));
    Span4Mux_v I__4830 (
            .O(N__23766),
            .I(N__23753));
    InMux I__4829 (
            .O(N__23763),
            .I(N__23748));
    InMux I__4828 (
            .O(N__23762),
            .I(N__23748));
    Span4Mux_s3_h I__4827 (
            .O(N__23759),
            .I(N__23745));
    Span4Mux_v I__4826 (
            .O(N__23756),
            .I(N__23740));
    Span4Mux_h I__4825 (
            .O(N__23753),
            .I(N__23740));
    LocalMux I__4824 (
            .O(N__23748),
            .I(data_in_field_131));
    Odrv4 I__4823 (
            .O(N__23745),
            .I(data_in_field_131));
    Odrv4 I__4822 (
            .O(N__23740),
            .I(data_in_field_131));
    InMux I__4821 (
            .O(N__23733),
            .I(N__23730));
    LocalMux I__4820 (
            .O(N__23730),
            .I(N__23727));
    Span4Mux_h I__4819 (
            .O(N__23727),
            .I(N__23724));
    Odrv4 I__4818 (
            .O(N__23724),
            .I(\c0.n8846 ));
    InMux I__4817 (
            .O(N__23721),
            .I(N__23715));
    InMux I__4816 (
            .O(N__23720),
            .I(N__23715));
    LocalMux I__4815 (
            .O(N__23715),
            .I(N__23711));
    InMux I__4814 (
            .O(N__23714),
            .I(N__23708));
    Span4Mux_v I__4813 (
            .O(N__23711),
            .I(N__23703));
    LocalMux I__4812 (
            .O(N__23708),
            .I(N__23700));
    InMux I__4811 (
            .O(N__23707),
            .I(N__23697));
    InMux I__4810 (
            .O(N__23706),
            .I(N__23694));
    Odrv4 I__4809 (
            .O(N__23703),
            .I(rand_data_2));
    Odrv12 I__4808 (
            .O(N__23700),
            .I(rand_data_2));
    LocalMux I__4807 (
            .O(N__23697),
            .I(rand_data_2));
    LocalMux I__4806 (
            .O(N__23694),
            .I(rand_data_2));
    InMux I__4805 (
            .O(N__23685),
            .I(N__23682));
    LocalMux I__4804 (
            .O(N__23682),
            .I(N__23679));
    Odrv12 I__4803 (
            .O(N__23679),
            .I(\c0.n30 ));
    InMux I__4802 (
            .O(N__23676),
            .I(N__23673));
    LocalMux I__4801 (
            .O(N__23673),
            .I(N__23670));
    Span4Mux_v I__4800 (
            .O(N__23670),
            .I(N__23664));
    InMux I__4799 (
            .O(N__23669),
            .I(N__23656));
    InMux I__4798 (
            .O(N__23668),
            .I(N__23653));
    InMux I__4797 (
            .O(N__23667),
            .I(N__23650));
    Span4Mux_h I__4796 (
            .O(N__23664),
            .I(N__23647));
    InMux I__4795 (
            .O(N__23663),
            .I(N__23640));
    InMux I__4794 (
            .O(N__23662),
            .I(N__23640));
    InMux I__4793 (
            .O(N__23661),
            .I(N__23640));
    InMux I__4792 (
            .O(N__23660),
            .I(N__23635));
    InMux I__4791 (
            .O(N__23659),
            .I(N__23635));
    LocalMux I__4790 (
            .O(N__23656),
            .I(N__23630));
    LocalMux I__4789 (
            .O(N__23653),
            .I(N__23630));
    LocalMux I__4788 (
            .O(N__23650),
            .I(N__23623));
    Span4Mux_h I__4787 (
            .O(N__23647),
            .I(N__23623));
    LocalMux I__4786 (
            .O(N__23640),
            .I(N__23623));
    LocalMux I__4785 (
            .O(N__23635),
            .I(FRAME_MATCHER_state_2));
    Odrv12 I__4784 (
            .O(N__23630),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__4783 (
            .O(N__23623),
            .I(FRAME_MATCHER_state_2));
    InMux I__4782 (
            .O(N__23616),
            .I(N__23613));
    LocalMux I__4781 (
            .O(N__23613),
            .I(N__23610));
    Span4Mux_s2_h I__4780 (
            .O(N__23610),
            .I(N__23606));
    InMux I__4779 (
            .O(N__23609),
            .I(N__23603));
    Span4Mux_h I__4778 (
            .O(N__23606),
            .I(N__23600));
    LocalMux I__4777 (
            .O(N__23603),
            .I(N__23597));
    Span4Mux_v I__4776 (
            .O(N__23600),
            .I(N__23594));
    Odrv4 I__4775 (
            .O(N__23597),
            .I(\c0.n7194 ));
    Odrv4 I__4774 (
            .O(N__23594),
            .I(\c0.n7194 ));
    InMux I__4773 (
            .O(N__23589),
            .I(N__23586));
    LocalMux I__4772 (
            .O(N__23586),
            .I(N__23583));
    Span4Mux_h I__4771 (
            .O(N__23583),
            .I(N__23580));
    Odrv4 I__4770 (
            .O(N__23580),
            .I(n9262));
    InMux I__4769 (
            .O(N__23577),
            .I(N__23568));
    InMux I__4768 (
            .O(N__23576),
            .I(N__23568));
    InMux I__4767 (
            .O(N__23575),
            .I(N__23568));
    LocalMux I__4766 (
            .O(N__23568),
            .I(data_in_6_2));
    CascadeMux I__4765 (
            .O(N__23565),
            .I(N__23555));
    InMux I__4764 (
            .O(N__23564),
            .I(N__23537));
    InMux I__4763 (
            .O(N__23563),
            .I(N__23528));
    InMux I__4762 (
            .O(N__23562),
            .I(N__23528));
    InMux I__4761 (
            .O(N__23561),
            .I(N__23528));
    InMux I__4760 (
            .O(N__23560),
            .I(N__23528));
    CascadeMux I__4759 (
            .O(N__23559),
            .I(N__23521));
    CascadeMux I__4758 (
            .O(N__23558),
            .I(N__23517));
    InMux I__4757 (
            .O(N__23555),
            .I(N__23509));
    InMux I__4756 (
            .O(N__23554),
            .I(N__23509));
    InMux I__4755 (
            .O(N__23553),
            .I(N__23509));
    CascadeMux I__4754 (
            .O(N__23552),
            .I(N__23503));
    InMux I__4753 (
            .O(N__23551),
            .I(N__23494));
    InMux I__4752 (
            .O(N__23550),
            .I(N__23494));
    InMux I__4751 (
            .O(N__23549),
            .I(N__23494));
    CascadeMux I__4750 (
            .O(N__23548),
            .I(N__23490));
    CascadeMux I__4749 (
            .O(N__23547),
            .I(N__23487));
    CascadeMux I__4748 (
            .O(N__23546),
            .I(N__23474));
    CascadeMux I__4747 (
            .O(N__23545),
            .I(N__23465));
    InMux I__4746 (
            .O(N__23544),
            .I(N__23460));
    InMux I__4745 (
            .O(N__23543),
            .I(N__23460));
    InMux I__4744 (
            .O(N__23542),
            .I(N__23457));
    InMux I__4743 (
            .O(N__23541),
            .I(N__23452));
    InMux I__4742 (
            .O(N__23540),
            .I(N__23452));
    LocalMux I__4741 (
            .O(N__23537),
            .I(N__23448));
    LocalMux I__4740 (
            .O(N__23528),
            .I(N__23445));
    InMux I__4739 (
            .O(N__23527),
            .I(N__23438));
    InMux I__4738 (
            .O(N__23526),
            .I(N__23438));
    InMux I__4737 (
            .O(N__23525),
            .I(N__23438));
    InMux I__4736 (
            .O(N__23524),
            .I(N__23433));
    InMux I__4735 (
            .O(N__23521),
            .I(N__23433));
    InMux I__4734 (
            .O(N__23520),
            .I(N__23430));
    InMux I__4733 (
            .O(N__23517),
            .I(N__23424));
    InMux I__4732 (
            .O(N__23516),
            .I(N__23424));
    LocalMux I__4731 (
            .O(N__23509),
            .I(N__23421));
    InMux I__4730 (
            .O(N__23508),
            .I(N__23415));
    InMux I__4729 (
            .O(N__23507),
            .I(N__23410));
    InMux I__4728 (
            .O(N__23506),
            .I(N__23410));
    InMux I__4727 (
            .O(N__23503),
            .I(N__23403));
    InMux I__4726 (
            .O(N__23502),
            .I(N__23403));
    InMux I__4725 (
            .O(N__23501),
            .I(N__23403));
    LocalMux I__4724 (
            .O(N__23494),
            .I(N__23397));
    InMux I__4723 (
            .O(N__23493),
            .I(N__23386));
    InMux I__4722 (
            .O(N__23490),
            .I(N__23386));
    InMux I__4721 (
            .O(N__23487),
            .I(N__23386));
    InMux I__4720 (
            .O(N__23486),
            .I(N__23386));
    InMux I__4719 (
            .O(N__23485),
            .I(N__23386));
    InMux I__4718 (
            .O(N__23484),
            .I(N__23383));
    InMux I__4717 (
            .O(N__23483),
            .I(N__23372));
    InMux I__4716 (
            .O(N__23482),
            .I(N__23372));
    InMux I__4715 (
            .O(N__23481),
            .I(N__23372));
    InMux I__4714 (
            .O(N__23480),
            .I(N__23372));
    InMux I__4713 (
            .O(N__23479),
            .I(N__23372));
    InMux I__4712 (
            .O(N__23478),
            .I(N__23361));
    InMux I__4711 (
            .O(N__23477),
            .I(N__23361));
    InMux I__4710 (
            .O(N__23474),
            .I(N__23361));
    InMux I__4709 (
            .O(N__23473),
            .I(N__23361));
    InMux I__4708 (
            .O(N__23472),
            .I(N__23361));
    InMux I__4707 (
            .O(N__23471),
            .I(N__23350));
    InMux I__4706 (
            .O(N__23470),
            .I(N__23350));
    InMux I__4705 (
            .O(N__23469),
            .I(N__23350));
    InMux I__4704 (
            .O(N__23468),
            .I(N__23350));
    InMux I__4703 (
            .O(N__23465),
            .I(N__23350));
    LocalMux I__4702 (
            .O(N__23460),
            .I(N__23345));
    LocalMux I__4701 (
            .O(N__23457),
            .I(N__23345));
    LocalMux I__4700 (
            .O(N__23452),
            .I(N__23342));
    InMux I__4699 (
            .O(N__23451),
            .I(N__23339));
    Span4Mux_v I__4698 (
            .O(N__23448),
            .I(N__23332));
    Span4Mux_v I__4697 (
            .O(N__23445),
            .I(N__23332));
    LocalMux I__4696 (
            .O(N__23438),
            .I(N__23332));
    LocalMux I__4695 (
            .O(N__23433),
            .I(N__23327));
    LocalMux I__4694 (
            .O(N__23430),
            .I(N__23327));
    InMux I__4693 (
            .O(N__23429),
            .I(N__23322));
    LocalMux I__4692 (
            .O(N__23424),
            .I(N__23319));
    Span4Mux_v I__4691 (
            .O(N__23421),
            .I(N__23316));
    InMux I__4690 (
            .O(N__23420),
            .I(N__23313));
    InMux I__4689 (
            .O(N__23419),
            .I(N__23308));
    InMux I__4688 (
            .O(N__23418),
            .I(N__23308));
    LocalMux I__4687 (
            .O(N__23415),
            .I(N__23301));
    LocalMux I__4686 (
            .O(N__23410),
            .I(N__23301));
    LocalMux I__4685 (
            .O(N__23403),
            .I(N__23301));
    InMux I__4684 (
            .O(N__23402),
            .I(N__23294));
    InMux I__4683 (
            .O(N__23401),
            .I(N__23294));
    InMux I__4682 (
            .O(N__23400),
            .I(N__23294));
    Span4Mux_v I__4681 (
            .O(N__23397),
            .I(N__23291));
    LocalMux I__4680 (
            .O(N__23386),
            .I(N__23286));
    LocalMux I__4679 (
            .O(N__23383),
            .I(N__23286));
    LocalMux I__4678 (
            .O(N__23372),
            .I(N__23275));
    LocalMux I__4677 (
            .O(N__23361),
            .I(N__23275));
    LocalMux I__4676 (
            .O(N__23350),
            .I(N__23275));
    Span4Mux_h I__4675 (
            .O(N__23345),
            .I(N__23275));
    Span4Mux_v I__4674 (
            .O(N__23342),
            .I(N__23275));
    LocalMux I__4673 (
            .O(N__23339),
            .I(N__23268));
    Span4Mux_v I__4672 (
            .O(N__23332),
            .I(N__23268));
    Span4Mux_v I__4671 (
            .O(N__23327),
            .I(N__23268));
    CascadeMux I__4670 (
            .O(N__23326),
            .I(N__23263));
    InMux I__4669 (
            .O(N__23325),
            .I(N__23259));
    LocalMux I__4668 (
            .O(N__23322),
            .I(N__23248));
    Span4Mux_v I__4667 (
            .O(N__23319),
            .I(N__23248));
    Span4Mux_h I__4666 (
            .O(N__23316),
            .I(N__23248));
    LocalMux I__4665 (
            .O(N__23313),
            .I(N__23248));
    LocalMux I__4664 (
            .O(N__23308),
            .I(N__23248));
    Span4Mux_v I__4663 (
            .O(N__23301),
            .I(N__23241));
    LocalMux I__4662 (
            .O(N__23294),
            .I(N__23241));
    Span4Mux_h I__4661 (
            .O(N__23291),
            .I(N__23241));
    Span4Mux_s3_h I__4660 (
            .O(N__23286),
            .I(N__23234));
    Span4Mux_v I__4659 (
            .O(N__23275),
            .I(N__23234));
    Span4Mux_h I__4658 (
            .O(N__23268),
            .I(N__23234));
    InMux I__4657 (
            .O(N__23267),
            .I(N__23229));
    InMux I__4656 (
            .O(N__23266),
            .I(N__23229));
    InMux I__4655 (
            .O(N__23263),
            .I(N__23224));
    InMux I__4654 (
            .O(N__23262),
            .I(N__23224));
    LocalMux I__4653 (
            .O(N__23259),
            .I(N__23219));
    Sp12to4 I__4652 (
            .O(N__23248),
            .I(N__23219));
    Span4Mux_v I__4651 (
            .O(N__23241),
            .I(N__23216));
    Span4Mux_v I__4650 (
            .O(N__23234),
            .I(N__23213));
    LocalMux I__4649 (
            .O(N__23229),
            .I(FRAME_MATCHER_state_0));
    LocalMux I__4648 (
            .O(N__23224),
            .I(FRAME_MATCHER_state_0));
    Odrv12 I__4647 (
            .O(N__23219),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__4646 (
            .O(N__23216),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__4645 (
            .O(N__23213),
            .I(FRAME_MATCHER_state_0));
    InMux I__4644 (
            .O(N__23202),
            .I(N__23199));
    LocalMux I__4643 (
            .O(N__23199),
            .I(N__23196));
    Span4Mux_h I__4642 (
            .O(N__23196),
            .I(N__23193));
    Odrv4 I__4641 (
            .O(N__23193),
            .I(n1893));
    InMux I__4640 (
            .O(N__23190),
            .I(N__23184));
    InMux I__4639 (
            .O(N__23189),
            .I(N__23184));
    LocalMux I__4638 (
            .O(N__23184),
            .I(data_in_7_2));
    InMux I__4637 (
            .O(N__23181),
            .I(N__23175));
    InMux I__4636 (
            .O(N__23180),
            .I(N__23175));
    LocalMux I__4635 (
            .O(N__23175),
            .I(data_in_8_2));
    InMux I__4634 (
            .O(N__23172),
            .I(N__23169));
    LocalMux I__4633 (
            .O(N__23169),
            .I(N__23166));
    Span4Mux_v I__4632 (
            .O(N__23166),
            .I(N__23162));
    InMux I__4631 (
            .O(N__23165),
            .I(N__23159));
    Odrv4 I__4630 (
            .O(N__23162),
            .I(data_in_10_2));
    LocalMux I__4629 (
            .O(N__23159),
            .I(data_in_10_2));
    InMux I__4628 (
            .O(N__23154),
            .I(N__23148));
    InMux I__4627 (
            .O(N__23153),
            .I(N__23148));
    LocalMux I__4626 (
            .O(N__23148),
            .I(data_in_9_2));
    InMux I__4625 (
            .O(N__23145),
            .I(N__23141));
    InMux I__4624 (
            .O(N__23144),
            .I(N__23138));
    LocalMux I__4623 (
            .O(N__23141),
            .I(N__23135));
    LocalMux I__4622 (
            .O(N__23138),
            .I(N__23132));
    Span4Mux_v I__4621 (
            .O(N__23135),
            .I(N__23129));
    Span4Mux_v I__4620 (
            .O(N__23132),
            .I(N__23126));
    Sp12to4 I__4619 (
            .O(N__23129),
            .I(N__23121));
    Sp12to4 I__4618 (
            .O(N__23126),
            .I(N__23121));
    Odrv12 I__4617 (
            .O(N__23121),
            .I(\c0.n8921 ));
    CascadeMux I__4616 (
            .O(N__23118),
            .I(\c0.n4562_cascade_ ));
    InMux I__4615 (
            .O(N__23115),
            .I(N__23109));
    InMux I__4614 (
            .O(N__23114),
            .I(N__23109));
    LocalMux I__4613 (
            .O(N__23109),
            .I(data_in_16_2));
    InMux I__4612 (
            .O(N__23106),
            .I(N__23100));
    InMux I__4611 (
            .O(N__23105),
            .I(N__23100));
    LocalMux I__4610 (
            .O(N__23100),
            .I(data_in_18_2));
    InMux I__4609 (
            .O(N__23097),
            .I(N__23093));
    InMux I__4608 (
            .O(N__23096),
            .I(N__23090));
    LocalMux I__4607 (
            .O(N__23093),
            .I(data_in_17_2));
    LocalMux I__4606 (
            .O(N__23090),
            .I(data_in_17_2));
    InMux I__4605 (
            .O(N__23085),
            .I(N__23082));
    LocalMux I__4604 (
            .O(N__23082),
            .I(N__23079));
    Span4Mux_h I__4603 (
            .O(N__23079),
            .I(N__23075));
    InMux I__4602 (
            .O(N__23078),
            .I(N__23072));
    Odrv4 I__4601 (
            .O(N__23075),
            .I(data_in_20_2));
    LocalMux I__4600 (
            .O(N__23072),
            .I(data_in_20_2));
    InMux I__4599 (
            .O(N__23067),
            .I(N__23061));
    InMux I__4598 (
            .O(N__23066),
            .I(N__23061));
    LocalMux I__4597 (
            .O(N__23061),
            .I(data_in_19_2));
    InMux I__4596 (
            .O(N__23058),
            .I(N__23052));
    InMux I__4595 (
            .O(N__23057),
            .I(N__23052));
    LocalMux I__4594 (
            .O(N__23052),
            .I(N__23049));
    Span4Mux_h I__4593 (
            .O(N__23049),
            .I(N__23046));
    Odrv4 I__4592 (
            .O(N__23046),
            .I(n7171));
    InMux I__4591 (
            .O(N__23043),
            .I(N__23040));
    LocalMux I__4590 (
            .O(N__23040),
            .I(N__23037));
    Odrv4 I__4589 (
            .O(N__23037),
            .I(\c0.n9668 ));
    InMux I__4588 (
            .O(N__23034),
            .I(N__23031));
    LocalMux I__4587 (
            .O(N__23031),
            .I(N__23028));
    Span12Mux_h I__4586 (
            .O(N__23028),
            .I(N__23024));
    InMux I__4585 (
            .O(N__23027),
            .I(N__23021));
    Odrv12 I__4584 (
            .O(N__23024),
            .I(\c0.n8878 ));
    LocalMux I__4583 (
            .O(N__23021),
            .I(\c0.n8878 ));
    InMux I__4582 (
            .O(N__23016),
            .I(N__23013));
    LocalMux I__4581 (
            .O(N__23013),
            .I(N__23009));
    InMux I__4580 (
            .O(N__23012),
            .I(N__23006));
    Span4Mux_h I__4579 (
            .O(N__23009),
            .I(N__23003));
    LocalMux I__4578 (
            .O(N__23006),
            .I(N__23000));
    Odrv4 I__4577 (
            .O(N__23003),
            .I(\c0.n8813 ));
    Odrv4 I__4576 (
            .O(N__23000),
            .I(\c0.n8813 ));
    InMux I__4575 (
            .O(N__22995),
            .I(N__22992));
    LocalMux I__4574 (
            .O(N__22992),
            .I(N__22988));
    InMux I__4573 (
            .O(N__22991),
            .I(N__22985));
    Span4Mux_h I__4572 (
            .O(N__22988),
            .I(N__22978));
    LocalMux I__4571 (
            .O(N__22985),
            .I(N__22978));
    CascadeMux I__4570 (
            .O(N__22984),
            .I(N__22973));
    InMux I__4569 (
            .O(N__22983),
            .I(N__22969));
    Span4Mux_h I__4568 (
            .O(N__22978),
            .I(N__22966));
    InMux I__4567 (
            .O(N__22977),
            .I(N__22957));
    InMux I__4566 (
            .O(N__22976),
            .I(N__22957));
    InMux I__4565 (
            .O(N__22973),
            .I(N__22957));
    InMux I__4564 (
            .O(N__22972),
            .I(N__22957));
    LocalMux I__4563 (
            .O(N__22969),
            .I(data_in_field_43));
    Odrv4 I__4562 (
            .O(N__22966),
            .I(data_in_field_43));
    LocalMux I__4561 (
            .O(N__22957),
            .I(data_in_field_43));
    InMux I__4560 (
            .O(N__22950),
            .I(N__22947));
    LocalMux I__4559 (
            .O(N__22947),
            .I(N__22944));
    Span4Mux_v I__4558 (
            .O(N__22944),
            .I(N__22941));
    Odrv4 I__4557 (
            .O(N__22941),
            .I(\c0.n28_adj_1619 ));
    CascadeMux I__4556 (
            .O(N__22938),
            .I(\c0.n29_adj_1620_cascade_ ));
    CascadeMux I__4555 (
            .O(N__22935),
            .I(N__22932));
    InMux I__4554 (
            .O(N__22932),
            .I(N__22929));
    LocalMux I__4553 (
            .O(N__22929),
            .I(N__22926));
    Odrv12 I__4552 (
            .O(N__22926),
            .I(\c0.data_in_frame_19_6 ));
    InMux I__4551 (
            .O(N__22923),
            .I(N__22920));
    LocalMux I__4550 (
            .O(N__22920),
            .I(N__22917));
    Span4Mux_h I__4549 (
            .O(N__22917),
            .I(N__22914));
    Odrv4 I__4548 (
            .O(N__22914),
            .I(n1901));
    InMux I__4547 (
            .O(N__22911),
            .I(N__22908));
    LocalMux I__4546 (
            .O(N__22908),
            .I(\c0.n9141 ));
    CascadeMux I__4545 (
            .O(N__22905),
            .I(\c0.n9138_cascade_ ));
    InMux I__4544 (
            .O(N__22902),
            .I(N__22899));
    LocalMux I__4543 (
            .O(N__22899),
            .I(N__22896));
    Span4Mux_h I__4542 (
            .O(N__22896),
            .I(N__22893));
    Span4Mux_v I__4541 (
            .O(N__22893),
            .I(N__22890));
    Span4Mux_v I__4540 (
            .O(N__22890),
            .I(N__22887));
    Odrv4 I__4539 (
            .O(N__22887),
            .I(\c0.n9132 ));
    InMux I__4538 (
            .O(N__22884),
            .I(N__22881));
    LocalMux I__4537 (
            .O(N__22881),
            .I(\c0.n9135 ));
    CascadeMux I__4536 (
            .O(N__22878),
            .I(\c0.n9614_cascade_ ));
    CascadeMux I__4535 (
            .O(N__22875),
            .I(\c0.n9617_cascade_ ));
    InMux I__4534 (
            .O(N__22872),
            .I(N__22869));
    LocalMux I__4533 (
            .O(N__22869),
            .I(N__22866));
    Odrv4 I__4532 (
            .O(N__22866),
            .I(\c0.tx2.r_Tx_Data_6 ));
    InMux I__4531 (
            .O(N__22863),
            .I(N__22857));
    InMux I__4530 (
            .O(N__22862),
            .I(N__22857));
    LocalMux I__4529 (
            .O(N__22857),
            .I(data_in_11_2));
    InMux I__4528 (
            .O(N__22854),
            .I(N__22848));
    InMux I__4527 (
            .O(N__22853),
            .I(N__22848));
    LocalMux I__4526 (
            .O(N__22848),
            .I(data_in_12_2));
    InMux I__4525 (
            .O(N__22845),
            .I(N__22839));
    InMux I__4524 (
            .O(N__22844),
            .I(N__22839));
    LocalMux I__4523 (
            .O(N__22839),
            .I(data_in_13_2));
    InMux I__4522 (
            .O(N__22836),
            .I(N__22830));
    InMux I__4521 (
            .O(N__22835),
            .I(N__22830));
    LocalMux I__4520 (
            .O(N__22830),
            .I(data_in_14_2));
    InMux I__4519 (
            .O(N__22827),
            .I(N__22821));
    InMux I__4518 (
            .O(N__22826),
            .I(N__22821));
    LocalMux I__4517 (
            .O(N__22821),
            .I(data_in_15_2));
    InMux I__4516 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__4515 (
            .O(N__22815),
            .I(N__22812));
    Odrv12 I__4514 (
            .O(N__22812),
            .I(\c0.n18_adj_1666 ));
    CascadeMux I__4513 (
            .O(N__22809),
            .I(N__22806));
    InMux I__4512 (
            .O(N__22806),
            .I(N__22801));
    InMux I__4511 (
            .O(N__22805),
            .I(N__22798));
    CascadeMux I__4510 (
            .O(N__22804),
            .I(N__22795));
    LocalMux I__4509 (
            .O(N__22801),
            .I(N__22792));
    LocalMux I__4508 (
            .O(N__22798),
            .I(N__22789));
    InMux I__4507 (
            .O(N__22795),
            .I(N__22786));
    Span4Mux_h I__4506 (
            .O(N__22792),
            .I(N__22783));
    Span4Mux_h I__4505 (
            .O(N__22789),
            .I(N__22780));
    LocalMux I__4504 (
            .O(N__22786),
            .I(N__22774));
    Span4Mux_v I__4503 (
            .O(N__22783),
            .I(N__22771));
    Span4Mux_v I__4502 (
            .O(N__22780),
            .I(N__22768));
    InMux I__4501 (
            .O(N__22779),
            .I(N__22765));
    InMux I__4500 (
            .O(N__22778),
            .I(N__22760));
    InMux I__4499 (
            .O(N__22777),
            .I(N__22760));
    Odrv4 I__4498 (
            .O(N__22774),
            .I(data_in_field_36));
    Odrv4 I__4497 (
            .O(N__22771),
            .I(data_in_field_36));
    Odrv4 I__4496 (
            .O(N__22768),
            .I(data_in_field_36));
    LocalMux I__4495 (
            .O(N__22765),
            .I(data_in_field_36));
    LocalMux I__4494 (
            .O(N__22760),
            .I(data_in_field_36));
    InMux I__4493 (
            .O(N__22749),
            .I(N__22746));
    LocalMux I__4492 (
            .O(N__22746),
            .I(N__22743));
    Span4Mux_h I__4491 (
            .O(N__22743),
            .I(N__22740));
    Odrv4 I__4490 (
            .O(N__22740),
            .I(\c0.n1645 ));
    CascadeMux I__4489 (
            .O(N__22737),
            .I(N__22733));
    CascadeMux I__4488 (
            .O(N__22736),
            .I(N__22730));
    InMux I__4487 (
            .O(N__22733),
            .I(N__22725));
    InMux I__4486 (
            .O(N__22730),
            .I(N__22722));
    InMux I__4485 (
            .O(N__22729),
            .I(N__22719));
    InMux I__4484 (
            .O(N__22728),
            .I(N__22716));
    LocalMux I__4483 (
            .O(N__22725),
            .I(N__22710));
    LocalMux I__4482 (
            .O(N__22722),
            .I(N__22710));
    LocalMux I__4481 (
            .O(N__22719),
            .I(N__22707));
    LocalMux I__4480 (
            .O(N__22716),
            .I(N__22704));
    InMux I__4479 (
            .O(N__22715),
            .I(N__22701));
    Span4Mux_v I__4478 (
            .O(N__22710),
            .I(N__22698));
    Span4Mux_s2_v I__4477 (
            .O(N__22707),
            .I(N__22693));
    Span4Mux_h I__4476 (
            .O(N__22704),
            .I(N__22693));
    LocalMux I__4475 (
            .O(N__22701),
            .I(data_in_field_62));
    Odrv4 I__4474 (
            .O(N__22698),
            .I(data_in_field_62));
    Odrv4 I__4473 (
            .O(N__22693),
            .I(data_in_field_62));
    InMux I__4472 (
            .O(N__22686),
            .I(N__22682));
    InMux I__4471 (
            .O(N__22685),
            .I(N__22679));
    LocalMux I__4470 (
            .O(N__22682),
            .I(N__22676));
    LocalMux I__4469 (
            .O(N__22679),
            .I(N__22668));
    Span4Mux_h I__4468 (
            .O(N__22676),
            .I(N__22665));
    InMux I__4467 (
            .O(N__22675),
            .I(N__22662));
    InMux I__4466 (
            .O(N__22674),
            .I(N__22657));
    InMux I__4465 (
            .O(N__22673),
            .I(N__22657));
    InMux I__4464 (
            .O(N__22672),
            .I(N__22654));
    InMux I__4463 (
            .O(N__22671),
            .I(N__22651));
    Span4Mux_v I__4462 (
            .O(N__22668),
            .I(N__22648));
    Span4Mux_v I__4461 (
            .O(N__22665),
            .I(N__22643));
    LocalMux I__4460 (
            .O(N__22662),
            .I(N__22643));
    LocalMux I__4459 (
            .O(N__22657),
            .I(N__22640));
    LocalMux I__4458 (
            .O(N__22654),
            .I(N__22637));
    LocalMux I__4457 (
            .O(N__22651),
            .I(data_in_field_46));
    Odrv4 I__4456 (
            .O(N__22648),
            .I(data_in_field_46));
    Odrv4 I__4455 (
            .O(N__22643),
            .I(data_in_field_46));
    Odrv12 I__4454 (
            .O(N__22640),
            .I(data_in_field_46));
    Odrv4 I__4453 (
            .O(N__22637),
            .I(data_in_field_46));
    CascadeMux I__4452 (
            .O(N__22626),
            .I(\c0.n9632_cascade_ ));
    InMux I__4451 (
            .O(N__22623),
            .I(N__22620));
    LocalMux I__4450 (
            .O(N__22620),
            .I(N__22616));
    CascadeMux I__4449 (
            .O(N__22619),
            .I(N__22611));
    Span4Mux_v I__4448 (
            .O(N__22616),
            .I(N__22608));
    InMux I__4447 (
            .O(N__22615),
            .I(N__22605));
    InMux I__4446 (
            .O(N__22614),
            .I(N__22601));
    InMux I__4445 (
            .O(N__22611),
            .I(N__22598));
    Span4Mux_v I__4444 (
            .O(N__22608),
            .I(N__22595));
    LocalMux I__4443 (
            .O(N__22605),
            .I(N__22592));
    InMux I__4442 (
            .O(N__22604),
            .I(N__22589));
    LocalMux I__4441 (
            .O(N__22601),
            .I(N__22586));
    LocalMux I__4440 (
            .O(N__22598),
            .I(\c0.data_in_field_38 ));
    Odrv4 I__4439 (
            .O(N__22595),
            .I(\c0.data_in_field_38 ));
    Odrv4 I__4438 (
            .O(N__22592),
            .I(\c0.data_in_field_38 ));
    LocalMux I__4437 (
            .O(N__22589),
            .I(\c0.data_in_field_38 ));
    Odrv12 I__4436 (
            .O(N__22586),
            .I(\c0.data_in_field_38 ));
    CascadeMux I__4435 (
            .O(N__22575),
            .I(N__22571));
    InMux I__4434 (
            .O(N__22574),
            .I(N__22567));
    InMux I__4433 (
            .O(N__22571),
            .I(N__22564));
    InMux I__4432 (
            .O(N__22570),
            .I(N__22559));
    LocalMux I__4431 (
            .O(N__22567),
            .I(N__22554));
    LocalMux I__4430 (
            .O(N__22564),
            .I(N__22554));
    InMux I__4429 (
            .O(N__22563),
            .I(N__22549));
    InMux I__4428 (
            .O(N__22562),
            .I(N__22549));
    LocalMux I__4427 (
            .O(N__22559),
            .I(N__22546));
    Span12Mux_s4_v I__4426 (
            .O(N__22554),
            .I(N__22543));
    LocalMux I__4425 (
            .O(N__22549),
            .I(data_in_field_126));
    Odrv4 I__4424 (
            .O(N__22546),
            .I(data_in_field_126));
    Odrv12 I__4423 (
            .O(N__22543),
            .I(data_in_field_126));
    CascadeMux I__4422 (
            .O(N__22536),
            .I(\c0.n9620_cascade_ ));
    InMux I__4421 (
            .O(N__22533),
            .I(N__22528));
    InMux I__4420 (
            .O(N__22532),
            .I(N__22525));
    InMux I__4419 (
            .O(N__22531),
            .I(N__22520));
    LocalMux I__4418 (
            .O(N__22528),
            .I(N__22517));
    LocalMux I__4417 (
            .O(N__22525),
            .I(N__22513));
    InMux I__4416 (
            .O(N__22524),
            .I(N__22510));
    InMux I__4415 (
            .O(N__22523),
            .I(N__22507));
    LocalMux I__4414 (
            .O(N__22520),
            .I(N__22502));
    Span4Mux_s2_v I__4413 (
            .O(N__22517),
            .I(N__22502));
    InMux I__4412 (
            .O(N__22516),
            .I(N__22499));
    Span4Mux_v I__4411 (
            .O(N__22513),
            .I(N__22494));
    LocalMux I__4410 (
            .O(N__22510),
            .I(N__22494));
    LocalMux I__4409 (
            .O(N__22507),
            .I(N__22489));
    Span4Mux_v I__4408 (
            .O(N__22502),
            .I(N__22489));
    LocalMux I__4407 (
            .O(N__22499),
            .I(N__22484));
    Span4Mux_h I__4406 (
            .O(N__22494),
            .I(N__22484));
    Odrv4 I__4405 (
            .O(N__22489),
            .I(data_in_field_94));
    Odrv4 I__4404 (
            .O(N__22484),
            .I(data_in_field_94));
    CascadeMux I__4403 (
            .O(N__22479),
            .I(\c0.n9626_cascade_ ));
    InMux I__4402 (
            .O(N__22476),
            .I(N__22472));
    InMux I__4401 (
            .O(N__22475),
            .I(N__22469));
    LocalMux I__4400 (
            .O(N__22472),
            .I(N__22464));
    LocalMux I__4399 (
            .O(N__22469),
            .I(N__22460));
    InMux I__4398 (
            .O(N__22468),
            .I(N__22457));
    InMux I__4397 (
            .O(N__22467),
            .I(N__22454));
    Span4Mux_v I__4396 (
            .O(N__22464),
            .I(N__22451));
    InMux I__4395 (
            .O(N__22463),
            .I(N__22448));
    Span4Mux_h I__4394 (
            .O(N__22460),
            .I(N__22443));
    LocalMux I__4393 (
            .O(N__22457),
            .I(N__22443));
    LocalMux I__4392 (
            .O(N__22454),
            .I(N__22438));
    Span4Mux_v I__4391 (
            .O(N__22451),
            .I(N__22438));
    LocalMux I__4390 (
            .O(N__22448),
            .I(data_in_field_44));
    Odrv4 I__4389 (
            .O(N__22443),
            .I(data_in_field_44));
    Odrv4 I__4388 (
            .O(N__22438),
            .I(data_in_field_44));
    InMux I__4387 (
            .O(N__22431),
            .I(N__22428));
    LocalMux I__4386 (
            .O(N__22428),
            .I(N__22425));
    Odrv12 I__4385 (
            .O(N__22425),
            .I(\c0.n9572 ));
    CascadeMux I__4384 (
            .O(N__22422),
            .I(N__22419));
    InMux I__4383 (
            .O(N__22419),
            .I(N__22415));
    InMux I__4382 (
            .O(N__22418),
            .I(N__22412));
    LocalMux I__4381 (
            .O(N__22415),
            .I(N__22408));
    LocalMux I__4380 (
            .O(N__22412),
            .I(N__22404));
    InMux I__4379 (
            .O(N__22411),
            .I(N__22401));
    Span12Mux_s6_v I__4378 (
            .O(N__22408),
            .I(N__22398));
    InMux I__4377 (
            .O(N__22407),
            .I(N__22395));
    Span4Mux_s3_v I__4376 (
            .O(N__22404),
            .I(N__22392));
    LocalMux I__4375 (
            .O(N__22401),
            .I(data_in_field_77));
    Odrv12 I__4374 (
            .O(N__22398),
            .I(data_in_field_77));
    LocalMux I__4373 (
            .O(N__22395),
            .I(data_in_field_77));
    Odrv4 I__4372 (
            .O(N__22392),
            .I(data_in_field_77));
    InMux I__4371 (
            .O(N__22383),
            .I(N__22379));
    InMux I__4370 (
            .O(N__22382),
            .I(N__22376));
    LocalMux I__4369 (
            .O(N__22379),
            .I(N__22372));
    LocalMux I__4368 (
            .O(N__22376),
            .I(N__22369));
    InMux I__4367 (
            .O(N__22375),
            .I(N__22365));
    Span4Mux_v I__4366 (
            .O(N__22372),
            .I(N__22362));
    Span4Mux_h I__4365 (
            .O(N__22369),
            .I(N__22359));
    InMux I__4364 (
            .O(N__22368),
            .I(N__22355));
    LocalMux I__4363 (
            .O(N__22365),
            .I(N__22352));
    Span4Mux_h I__4362 (
            .O(N__22362),
            .I(N__22349));
    Span4Mux_h I__4361 (
            .O(N__22359),
            .I(N__22346));
    InMux I__4360 (
            .O(N__22358),
            .I(N__22343));
    LocalMux I__4359 (
            .O(N__22355),
            .I(data_in_field_49));
    Odrv12 I__4358 (
            .O(N__22352),
            .I(data_in_field_49));
    Odrv4 I__4357 (
            .O(N__22349),
            .I(data_in_field_49));
    Odrv4 I__4356 (
            .O(N__22346),
            .I(data_in_field_49));
    LocalMux I__4355 (
            .O(N__22343),
            .I(data_in_field_49));
    CascadeMux I__4354 (
            .O(N__22332),
            .I(\c0.n8887_cascade_ ));
    InMux I__4353 (
            .O(N__22329),
            .I(N__22323));
    InMux I__4352 (
            .O(N__22328),
            .I(N__22320));
    InMux I__4351 (
            .O(N__22327),
            .I(N__22317));
    InMux I__4350 (
            .O(N__22326),
            .I(N__22314));
    LocalMux I__4349 (
            .O(N__22323),
            .I(data_in_field_120));
    LocalMux I__4348 (
            .O(N__22320),
            .I(data_in_field_120));
    LocalMux I__4347 (
            .O(N__22317),
            .I(data_in_field_120));
    LocalMux I__4346 (
            .O(N__22314),
            .I(data_in_field_120));
    InMux I__4345 (
            .O(N__22305),
            .I(N__22301));
    InMux I__4344 (
            .O(N__22304),
            .I(N__22298));
    LocalMux I__4343 (
            .O(N__22301),
            .I(N__22295));
    LocalMux I__4342 (
            .O(N__22298),
            .I(N__22291));
    Span4Mux_v I__4341 (
            .O(N__22295),
            .I(N__22288));
    InMux I__4340 (
            .O(N__22294),
            .I(N__22285));
    Span4Mux_v I__4339 (
            .O(N__22291),
            .I(N__22279));
    Span4Mux_v I__4338 (
            .O(N__22288),
            .I(N__22279));
    LocalMux I__4337 (
            .O(N__22285),
            .I(N__22276));
    InMux I__4336 (
            .O(N__22284),
            .I(N__22273));
    Span4Mux_h I__4335 (
            .O(N__22279),
            .I(N__22270));
    Odrv4 I__4334 (
            .O(N__22276),
            .I(rand_data_30));
    LocalMux I__4333 (
            .O(N__22273),
            .I(rand_data_30));
    Odrv4 I__4332 (
            .O(N__22270),
            .I(rand_data_30));
    InMux I__4331 (
            .O(N__22263),
            .I(N__22256));
    InMux I__4330 (
            .O(N__22262),
            .I(N__22256));
    InMux I__4329 (
            .O(N__22261),
            .I(N__22253));
    LocalMux I__4328 (
            .O(N__22256),
            .I(N__22250));
    LocalMux I__4327 (
            .O(N__22253),
            .I(\c0.n8785 ));
    Odrv12 I__4326 (
            .O(N__22250),
            .I(\c0.n8785 ));
    InMux I__4325 (
            .O(N__22245),
            .I(N__22242));
    LocalMux I__4324 (
            .O(N__22242),
            .I(N__22239));
    Span4Mux_h I__4323 (
            .O(N__22239),
            .I(N__22235));
    InMux I__4322 (
            .O(N__22238),
            .I(N__22232));
    Odrv4 I__4321 (
            .O(N__22235),
            .I(\c0.n8887 ));
    LocalMux I__4320 (
            .O(N__22232),
            .I(\c0.n8887 ));
    CascadeMux I__4319 (
            .O(N__22227),
            .I(\c0.n4240_cascade_ ));
    InMux I__4318 (
            .O(N__22224),
            .I(N__22220));
    InMux I__4317 (
            .O(N__22223),
            .I(N__22217));
    LocalMux I__4316 (
            .O(N__22220),
            .I(N__22214));
    LocalMux I__4315 (
            .O(N__22217),
            .I(N__22209));
    Span4Mux_v I__4314 (
            .O(N__22214),
            .I(N__22209));
    Span4Mux_v I__4313 (
            .O(N__22209),
            .I(N__22204));
    InMux I__4312 (
            .O(N__22208),
            .I(N__22201));
    InMux I__4311 (
            .O(N__22207),
            .I(N__22196));
    Sp12to4 I__4310 (
            .O(N__22204),
            .I(N__22191));
    LocalMux I__4309 (
            .O(N__22201),
            .I(N__22191));
    InMux I__4308 (
            .O(N__22200),
            .I(N__22186));
    InMux I__4307 (
            .O(N__22199),
            .I(N__22186));
    LocalMux I__4306 (
            .O(N__22196),
            .I(\c0.data_in_field_13 ));
    Odrv12 I__4305 (
            .O(N__22191),
            .I(\c0.data_in_field_13 ));
    LocalMux I__4304 (
            .O(N__22186),
            .I(\c0.data_in_field_13 ));
    InMux I__4303 (
            .O(N__22179),
            .I(N__22176));
    LocalMux I__4302 (
            .O(N__22176),
            .I(N__22173));
    Span4Mux_s2_h I__4301 (
            .O(N__22173),
            .I(N__22170));
    Span4Mux_h I__4300 (
            .O(N__22170),
            .I(N__22167));
    Odrv4 I__4299 (
            .O(N__22167),
            .I(\c0.n44_adj_1609 ));
    InMux I__4298 (
            .O(N__22164),
            .I(N__22161));
    LocalMux I__4297 (
            .O(N__22161),
            .I(\c0.n4553 ));
    InMux I__4296 (
            .O(N__22158),
            .I(N__22152));
    InMux I__4295 (
            .O(N__22157),
            .I(N__22152));
    LocalMux I__4294 (
            .O(N__22152),
            .I(N__22148));
    InMux I__4293 (
            .O(N__22151),
            .I(N__22143));
    Span4Mux_v I__4292 (
            .O(N__22148),
            .I(N__22140));
    InMux I__4291 (
            .O(N__22147),
            .I(N__22135));
    InMux I__4290 (
            .O(N__22146),
            .I(N__22135));
    LocalMux I__4289 (
            .O(N__22143),
            .I(data_in_field_53));
    Odrv4 I__4288 (
            .O(N__22140),
            .I(data_in_field_53));
    LocalMux I__4287 (
            .O(N__22135),
            .I(data_in_field_53));
    CascadeMux I__4286 (
            .O(N__22128),
            .I(N__22125));
    InMux I__4285 (
            .O(N__22125),
            .I(N__22122));
    LocalMux I__4284 (
            .O(N__22122),
            .I(N__22119));
    Odrv12 I__4283 (
            .O(N__22119),
            .I(\c0.n8964 ));
    InMux I__4282 (
            .O(N__22116),
            .I(N__22113));
    LocalMux I__4281 (
            .O(N__22113),
            .I(N__22110));
    IoSpan4Mux I__4280 (
            .O(N__22110),
            .I(N__22107));
    IoSpan4Mux I__4279 (
            .O(N__22107),
            .I(N__22104));
    Odrv4 I__4278 (
            .O(N__22104),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__4277 (
            .O(N__22101),
            .I(N__22098));
    InMux I__4276 (
            .O(N__22098),
            .I(N__22094));
    InMux I__4275 (
            .O(N__22097),
            .I(N__22091));
    LocalMux I__4274 (
            .O(N__22094),
            .I(N__22088));
    LocalMux I__4273 (
            .O(N__22091),
            .I(N__22085));
    Span4Mux_v I__4272 (
            .O(N__22088),
            .I(N__22082));
    Span4Mux_v I__4271 (
            .O(N__22085),
            .I(N__22079));
    Span4Mux_h I__4270 (
            .O(N__22082),
            .I(N__22076));
    Span4Mux_h I__4269 (
            .O(N__22079),
            .I(N__22073));
    Odrv4 I__4268 (
            .O(N__22076),
            .I(\c0.n8942 ));
    Odrv4 I__4267 (
            .O(N__22073),
            .I(\c0.n8942 ));
    InMux I__4266 (
            .O(N__22068),
            .I(N__22065));
    LocalMux I__4265 (
            .O(N__22065),
            .I(N__22062));
    Span4Mux_s2_h I__4264 (
            .O(N__22062),
            .I(N__22059));
    Span4Mux_v I__4263 (
            .O(N__22059),
            .I(N__22053));
    InMux I__4262 (
            .O(N__22058),
            .I(N__22050));
    CascadeMux I__4261 (
            .O(N__22057),
            .I(N__22047));
    InMux I__4260 (
            .O(N__22056),
            .I(N__22044));
    Span4Mux_h I__4259 (
            .O(N__22053),
            .I(N__22039));
    LocalMux I__4258 (
            .O(N__22050),
            .I(N__22039));
    InMux I__4257 (
            .O(N__22047),
            .I(N__22036));
    LocalMux I__4256 (
            .O(N__22044),
            .I(N__22031));
    Span4Mux_s3_v I__4255 (
            .O(N__22039),
            .I(N__22031));
    LocalMux I__4254 (
            .O(N__22036),
            .I(N__22028));
    Odrv4 I__4253 (
            .O(N__22031),
            .I(data_in_field_57));
    Odrv12 I__4252 (
            .O(N__22028),
            .I(data_in_field_57));
    InMux I__4251 (
            .O(N__22023),
            .I(N__22019));
    InMux I__4250 (
            .O(N__22022),
            .I(N__22013));
    LocalMux I__4249 (
            .O(N__22019),
            .I(N__22010));
    InMux I__4248 (
            .O(N__22018),
            .I(N__22007));
    InMux I__4247 (
            .O(N__22017),
            .I(N__22004));
    InMux I__4246 (
            .O(N__22016),
            .I(N__22001));
    LocalMux I__4245 (
            .O(N__22013),
            .I(N__21997));
    Span4Mux_v I__4244 (
            .O(N__22010),
            .I(N__21994));
    LocalMux I__4243 (
            .O(N__22007),
            .I(N__21991));
    LocalMux I__4242 (
            .O(N__22004),
            .I(N__21986));
    LocalMux I__4241 (
            .O(N__22001),
            .I(N__21986));
    InMux I__4240 (
            .O(N__22000),
            .I(N__21983));
    Span4Mux_s2_v I__4239 (
            .O(N__21997),
            .I(N__21980));
    Span4Mux_h I__4238 (
            .O(N__21994),
            .I(N__21973));
    Span4Mux_s3_h I__4237 (
            .O(N__21991),
            .I(N__21973));
    Span4Mux_v I__4236 (
            .O(N__21986),
            .I(N__21973));
    LocalMux I__4235 (
            .O(N__21983),
            .I(data_in_field_93));
    Odrv4 I__4234 (
            .O(N__21980),
            .I(data_in_field_93));
    Odrv4 I__4233 (
            .O(N__21973),
            .I(data_in_field_93));
    CascadeMux I__4232 (
            .O(N__21966),
            .I(N__21963));
    InMux I__4231 (
            .O(N__21963),
            .I(N__21960));
    LocalMux I__4230 (
            .O(N__21960),
            .I(N__21957));
    Span4Mux_h I__4229 (
            .O(N__21957),
            .I(N__21954));
    Odrv4 I__4228 (
            .O(N__21954),
            .I(\c0.n4390 ));
    InMux I__4227 (
            .O(N__21951),
            .I(N__21946));
    InMux I__4226 (
            .O(N__21950),
            .I(N__21943));
    CascadeMux I__4225 (
            .O(N__21949),
            .I(N__21939));
    LocalMux I__4224 (
            .O(N__21946),
            .I(N__21936));
    LocalMux I__4223 (
            .O(N__21943),
            .I(N__21933));
    InMux I__4222 (
            .O(N__21942),
            .I(N__21930));
    InMux I__4221 (
            .O(N__21939),
            .I(N__21925));
    Span4Mux_s3_v I__4220 (
            .O(N__21936),
            .I(N__21922));
    Span4Mux_h I__4219 (
            .O(N__21933),
            .I(N__21917));
    LocalMux I__4218 (
            .O(N__21930),
            .I(N__21917));
    InMux I__4217 (
            .O(N__21929),
            .I(N__21914));
    InMux I__4216 (
            .O(N__21928),
            .I(N__21911));
    LocalMux I__4215 (
            .O(N__21925),
            .I(N__21908));
    Span4Mux_h I__4214 (
            .O(N__21922),
            .I(N__21903));
    Span4Mux_h I__4213 (
            .O(N__21917),
            .I(N__21903));
    LocalMux I__4212 (
            .O(N__21914),
            .I(data_in_field_87));
    LocalMux I__4211 (
            .O(N__21911),
            .I(data_in_field_87));
    Odrv12 I__4210 (
            .O(N__21908),
            .I(data_in_field_87));
    Odrv4 I__4209 (
            .O(N__21903),
            .I(data_in_field_87));
    CascadeMux I__4208 (
            .O(N__21894),
            .I(N__21888));
    InMux I__4207 (
            .O(N__21893),
            .I(N__21885));
    InMux I__4206 (
            .O(N__21892),
            .I(N__21882));
    InMux I__4205 (
            .O(N__21891),
            .I(N__21877));
    InMux I__4204 (
            .O(N__21888),
            .I(N__21874));
    LocalMux I__4203 (
            .O(N__21885),
            .I(N__21870));
    LocalMux I__4202 (
            .O(N__21882),
            .I(N__21867));
    InMux I__4201 (
            .O(N__21881),
            .I(N__21864));
    InMux I__4200 (
            .O(N__21880),
            .I(N__21861));
    LocalMux I__4199 (
            .O(N__21877),
            .I(N__21858));
    LocalMux I__4198 (
            .O(N__21874),
            .I(N__21855));
    InMux I__4197 (
            .O(N__21873),
            .I(N__21852));
    Span4Mux_h I__4196 (
            .O(N__21870),
            .I(N__21849));
    Span4Mux_v I__4195 (
            .O(N__21867),
            .I(N__21844));
    LocalMux I__4194 (
            .O(N__21864),
            .I(N__21844));
    LocalMux I__4193 (
            .O(N__21861),
            .I(N__21837));
    Span4Mux_s2_v I__4192 (
            .O(N__21858),
            .I(N__21837));
    Span4Mux_h I__4191 (
            .O(N__21855),
            .I(N__21837));
    LocalMux I__4190 (
            .O(N__21852),
            .I(data_in_field_91));
    Odrv4 I__4189 (
            .O(N__21849),
            .I(data_in_field_91));
    Odrv4 I__4188 (
            .O(N__21844),
            .I(data_in_field_91));
    Odrv4 I__4187 (
            .O(N__21837),
            .I(data_in_field_91));
    CascadeMux I__4186 (
            .O(N__21828),
            .I(N__21825));
    InMux I__4185 (
            .O(N__21825),
            .I(N__21822));
    LocalMux I__4184 (
            .O(N__21822),
            .I(N__21818));
    InMux I__4183 (
            .O(N__21821),
            .I(N__21815));
    Span4Mux_h I__4182 (
            .O(N__21818),
            .I(N__21812));
    LocalMux I__4181 (
            .O(N__21815),
            .I(\c0.n8909 ));
    Odrv4 I__4180 (
            .O(N__21812),
            .I(\c0.n8909 ));
    InMux I__4179 (
            .O(N__21807),
            .I(N__21804));
    LocalMux I__4178 (
            .O(N__21804),
            .I(N__21801));
    Span4Mux_h I__4177 (
            .O(N__21801),
            .I(N__21798));
    Odrv4 I__4176 (
            .O(N__21798),
            .I(\c0.n4197 ));
    InMux I__4175 (
            .O(N__21795),
            .I(N__21788));
    InMux I__4174 (
            .O(N__21794),
            .I(N__21788));
    CascadeMux I__4173 (
            .O(N__21793),
            .I(N__21784));
    LocalMux I__4172 (
            .O(N__21788),
            .I(N__21781));
    InMux I__4171 (
            .O(N__21787),
            .I(N__21778));
    InMux I__4170 (
            .O(N__21784),
            .I(N__21775));
    Span4Mux_v I__4169 (
            .O(N__21781),
            .I(N__21771));
    LocalMux I__4168 (
            .O(N__21778),
            .I(N__21766));
    LocalMux I__4167 (
            .O(N__21775),
            .I(N__21766));
    InMux I__4166 (
            .O(N__21774),
            .I(N__21763));
    Span4Mux_h I__4165 (
            .O(N__21771),
            .I(N__21758));
    Span4Mux_v I__4164 (
            .O(N__21766),
            .I(N__21758));
    LocalMux I__4163 (
            .O(N__21763),
            .I(data_in_field_60));
    Odrv4 I__4162 (
            .O(N__21758),
            .I(data_in_field_60));
    CascadeMux I__4161 (
            .O(N__21753),
            .I(\c0.n4197_cascade_ ));
    CascadeMux I__4160 (
            .O(N__21750),
            .I(N__21747));
    InMux I__4159 (
            .O(N__21747),
            .I(N__21744));
    LocalMux I__4158 (
            .O(N__21744),
            .I(N__21741));
    Span4Mux_h I__4157 (
            .O(N__21741),
            .I(N__21738));
    Odrv4 I__4156 (
            .O(N__21738),
            .I(\c0.n4399 ));
    CascadeMux I__4155 (
            .O(N__21735),
            .I(N__21732));
    InMux I__4154 (
            .O(N__21732),
            .I(N__21727));
    InMux I__4153 (
            .O(N__21731),
            .I(N__21722));
    InMux I__4152 (
            .O(N__21730),
            .I(N__21722));
    LocalMux I__4151 (
            .O(N__21727),
            .I(N__21719));
    LocalMux I__4150 (
            .O(N__21722),
            .I(N__21714));
    Span4Mux_h I__4149 (
            .O(N__21719),
            .I(N__21711));
    InMux I__4148 (
            .O(N__21718),
            .I(N__21708));
    InMux I__4147 (
            .O(N__21717),
            .I(N__21705));
    Span4Mux_h I__4146 (
            .O(N__21714),
            .I(N__21698));
    Span4Mux_v I__4145 (
            .O(N__21711),
            .I(N__21698));
    LocalMux I__4144 (
            .O(N__21708),
            .I(N__21698));
    LocalMux I__4143 (
            .O(N__21705),
            .I(data_in_field_61));
    Odrv4 I__4142 (
            .O(N__21698),
            .I(data_in_field_61));
    CascadeMux I__4141 (
            .O(N__21693),
            .I(\c0.n4399_cascade_ ));
    InMux I__4140 (
            .O(N__21690),
            .I(N__21687));
    LocalMux I__4139 (
            .O(N__21687),
            .I(N__21683));
    InMux I__4138 (
            .O(N__21686),
            .I(N__21680));
    Odrv12 I__4137 (
            .O(N__21683),
            .I(\c0.n4288 ));
    LocalMux I__4136 (
            .O(N__21680),
            .I(\c0.n4288 ));
    InMux I__4135 (
            .O(N__21675),
            .I(N__21672));
    LocalMux I__4134 (
            .O(N__21672),
            .I(\c0.n10 ));
    InMux I__4133 (
            .O(N__21669),
            .I(N__21666));
    LocalMux I__4132 (
            .O(N__21666),
            .I(N__21663));
    Span4Mux_v I__4131 (
            .O(N__21663),
            .I(N__21658));
    CascadeMux I__4130 (
            .O(N__21662),
            .I(N__21655));
    InMux I__4129 (
            .O(N__21661),
            .I(N__21651));
    Span4Mux_h I__4128 (
            .O(N__21658),
            .I(N__21647));
    InMux I__4127 (
            .O(N__21655),
            .I(N__21642));
    InMux I__4126 (
            .O(N__21654),
            .I(N__21642));
    LocalMux I__4125 (
            .O(N__21651),
            .I(N__21639));
    InMux I__4124 (
            .O(N__21650),
            .I(N__21636));
    Odrv4 I__4123 (
            .O(N__21647),
            .I(rand_data_9));
    LocalMux I__4122 (
            .O(N__21642),
            .I(rand_data_9));
    Odrv4 I__4121 (
            .O(N__21639),
            .I(rand_data_9));
    LocalMux I__4120 (
            .O(N__21636),
            .I(rand_data_9));
    InMux I__4119 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__4118 (
            .O(N__21624),
            .I(N__21619));
    InMux I__4117 (
            .O(N__21623),
            .I(N__21616));
    InMux I__4116 (
            .O(N__21622),
            .I(N__21613));
    Span4Mux_h I__4115 (
            .O(N__21619),
            .I(N__21608));
    LocalMux I__4114 (
            .O(N__21616),
            .I(N__21603));
    LocalMux I__4113 (
            .O(N__21613),
            .I(N__21603));
    InMux I__4112 (
            .O(N__21612),
            .I(N__21598));
    InMux I__4111 (
            .O(N__21611),
            .I(N__21598));
    Odrv4 I__4110 (
            .O(N__21608),
            .I(data_in_field_121));
    Odrv12 I__4109 (
            .O(N__21603),
            .I(data_in_field_121));
    LocalMux I__4108 (
            .O(N__21598),
            .I(data_in_field_121));
    InMux I__4107 (
            .O(N__21591),
            .I(N__21585));
    InMux I__4106 (
            .O(N__21590),
            .I(N__21585));
    LocalMux I__4105 (
            .O(N__21585),
            .I(N__21581));
    InMux I__4104 (
            .O(N__21584),
            .I(N__21578));
    Span12Mux_s4_v I__4103 (
            .O(N__21581),
            .I(N__21573));
    LocalMux I__4102 (
            .O(N__21578),
            .I(N__21570));
    InMux I__4101 (
            .O(N__21577),
            .I(N__21567));
    InMux I__4100 (
            .O(N__21576),
            .I(N__21564));
    Odrv12 I__4099 (
            .O(N__21573),
            .I(rand_data_15));
    Odrv4 I__4098 (
            .O(N__21570),
            .I(rand_data_15));
    LocalMux I__4097 (
            .O(N__21567),
            .I(rand_data_15));
    LocalMux I__4096 (
            .O(N__21564),
            .I(rand_data_15));
    InMux I__4095 (
            .O(N__21555),
            .I(N__21551));
    InMux I__4094 (
            .O(N__21554),
            .I(N__21546));
    LocalMux I__4093 (
            .O(N__21551),
            .I(N__21543));
    InMux I__4092 (
            .O(N__21550),
            .I(N__21538));
    InMux I__4091 (
            .O(N__21549),
            .I(N__21538));
    LocalMux I__4090 (
            .O(N__21546),
            .I(N__21532));
    Span4Mux_s1_v I__4089 (
            .O(N__21543),
            .I(N__21532));
    LocalMux I__4088 (
            .O(N__21538),
            .I(N__21529));
    InMux I__4087 (
            .O(N__21537),
            .I(N__21525));
    Span4Mux_v I__4086 (
            .O(N__21532),
            .I(N__21522));
    Span4Mux_h I__4085 (
            .O(N__21529),
            .I(N__21519));
    InMux I__4084 (
            .O(N__21528),
            .I(N__21516));
    LocalMux I__4083 (
            .O(N__21525),
            .I(data_in_field_143));
    Odrv4 I__4082 (
            .O(N__21522),
            .I(data_in_field_143));
    Odrv4 I__4081 (
            .O(N__21519),
            .I(data_in_field_143));
    LocalMux I__4080 (
            .O(N__21516),
            .I(data_in_field_143));
    InMux I__4079 (
            .O(N__21507),
            .I(N__21502));
    InMux I__4078 (
            .O(N__21506),
            .I(N__21499));
    InMux I__4077 (
            .O(N__21505),
            .I(N__21496));
    LocalMux I__4076 (
            .O(N__21502),
            .I(N__21493));
    LocalMux I__4075 (
            .O(N__21499),
            .I(N__21490));
    LocalMux I__4074 (
            .O(N__21496),
            .I(N__21487));
    Span4Mux_h I__4073 (
            .O(N__21493),
            .I(N__21483));
    Span4Mux_v I__4072 (
            .O(N__21490),
            .I(N__21478));
    Span4Mux_h I__4071 (
            .O(N__21487),
            .I(N__21478));
    InMux I__4070 (
            .O(N__21486),
            .I(N__21475));
    Span4Mux_h I__4069 (
            .O(N__21483),
            .I(N__21472));
    Odrv4 I__4068 (
            .O(N__21478),
            .I(rand_data_28));
    LocalMux I__4067 (
            .O(N__21475),
            .I(rand_data_28));
    Odrv4 I__4066 (
            .O(N__21472),
            .I(rand_data_28));
    InMux I__4065 (
            .O(N__21465),
            .I(N__21460));
    InMux I__4064 (
            .O(N__21464),
            .I(N__21455));
    InMux I__4063 (
            .O(N__21463),
            .I(N__21452));
    LocalMux I__4062 (
            .O(N__21460),
            .I(N__21449));
    InMux I__4061 (
            .O(N__21459),
            .I(N__21446));
    InMux I__4060 (
            .O(N__21458),
            .I(N__21443));
    LocalMux I__4059 (
            .O(N__21455),
            .I(rand_data_13));
    LocalMux I__4058 (
            .O(N__21452),
            .I(rand_data_13));
    Odrv4 I__4057 (
            .O(N__21449),
            .I(rand_data_13));
    LocalMux I__4056 (
            .O(N__21446),
            .I(rand_data_13));
    LocalMux I__4055 (
            .O(N__21443),
            .I(rand_data_13));
    InMux I__4054 (
            .O(N__21432),
            .I(N__21426));
    InMux I__4053 (
            .O(N__21431),
            .I(N__21423));
    InMux I__4052 (
            .O(N__21430),
            .I(N__21420));
    CascadeMux I__4051 (
            .O(N__21429),
            .I(N__21417));
    LocalMux I__4050 (
            .O(N__21426),
            .I(N__21414));
    LocalMux I__4049 (
            .O(N__21423),
            .I(N__21411));
    LocalMux I__4048 (
            .O(N__21420),
            .I(N__21406));
    InMux I__4047 (
            .O(N__21417),
            .I(N__21403));
    Span4Mux_v I__4046 (
            .O(N__21414),
            .I(N__21400));
    Span4Mux_v I__4045 (
            .O(N__21411),
            .I(N__21397));
    InMux I__4044 (
            .O(N__21410),
            .I(N__21394));
    InMux I__4043 (
            .O(N__21409),
            .I(N__21391));
    Span4Mux_h I__4042 (
            .O(N__21406),
            .I(N__21388));
    LocalMux I__4041 (
            .O(N__21403),
            .I(\c0.data_in_field_29 ));
    Odrv4 I__4040 (
            .O(N__21400),
            .I(\c0.data_in_field_29 ));
    Odrv4 I__4039 (
            .O(N__21397),
            .I(\c0.data_in_field_29 ));
    LocalMux I__4038 (
            .O(N__21394),
            .I(\c0.data_in_field_29 ));
    LocalMux I__4037 (
            .O(N__21391),
            .I(\c0.data_in_field_29 ));
    Odrv4 I__4036 (
            .O(N__21388),
            .I(\c0.data_in_field_29 ));
    CascadeMux I__4035 (
            .O(N__21375),
            .I(N__21371));
    InMux I__4034 (
            .O(N__21374),
            .I(N__21368));
    InMux I__4033 (
            .O(N__21371),
            .I(N__21364));
    LocalMux I__4032 (
            .O(N__21368),
            .I(N__21361));
    InMux I__4031 (
            .O(N__21367),
            .I(N__21358));
    LocalMux I__4030 (
            .O(N__21364),
            .I(N__21354));
    Span4Mux_v I__4029 (
            .O(N__21361),
            .I(N__21351));
    LocalMux I__4028 (
            .O(N__21358),
            .I(N__21348));
    InMux I__4027 (
            .O(N__21357),
            .I(N__21345));
    Span4Mux_s3_h I__4026 (
            .O(N__21354),
            .I(N__21342));
    Span4Mux_h I__4025 (
            .O(N__21351),
            .I(N__21337));
    Span4Mux_s3_h I__4024 (
            .O(N__21348),
            .I(N__21337));
    LocalMux I__4023 (
            .O(N__21345),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__4022 (
            .O(N__21342),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__4021 (
            .O(N__21337),
            .I(\c0.data_in_field_21 ));
    CascadeMux I__4020 (
            .O(N__21330),
            .I(\c0.n9608_cascade_ ));
    InMux I__4019 (
            .O(N__21327),
            .I(N__21323));
    CascadeMux I__4018 (
            .O(N__21326),
            .I(N__21319));
    LocalMux I__4017 (
            .O(N__21323),
            .I(N__21316));
    CascadeMux I__4016 (
            .O(N__21322),
            .I(N__21312));
    InMux I__4015 (
            .O(N__21319),
            .I(N__21309));
    Span4Mux_v I__4014 (
            .O(N__21316),
            .I(N__21306));
    InMux I__4013 (
            .O(N__21315),
            .I(N__21303));
    InMux I__4012 (
            .O(N__21312),
            .I(N__21300));
    LocalMux I__4011 (
            .O(N__21309),
            .I(\c0.data_in_field_5 ));
    Odrv4 I__4010 (
            .O(N__21306),
            .I(\c0.data_in_field_5 ));
    LocalMux I__4009 (
            .O(N__21303),
            .I(\c0.data_in_field_5 ));
    LocalMux I__4008 (
            .O(N__21300),
            .I(\c0.data_in_field_5 ));
    InMux I__4007 (
            .O(N__21291),
            .I(N__21288));
    LocalMux I__4006 (
            .O(N__21288),
            .I(N__21285));
    Span4Mux_s2_v I__4005 (
            .O(N__21285),
            .I(N__21282));
    Odrv4 I__4004 (
            .O(N__21282),
            .I(\c0.n9147 ));
    InMux I__4003 (
            .O(N__21279),
            .I(N__21275));
    InMux I__4002 (
            .O(N__21278),
            .I(N__21271));
    LocalMux I__4001 (
            .O(N__21275),
            .I(N__21268));
    InMux I__4000 (
            .O(N__21274),
            .I(N__21265));
    LocalMux I__3999 (
            .O(N__21271),
            .I(N__21262));
    Span4Mux_h I__3998 (
            .O(N__21268),
            .I(N__21259));
    LocalMux I__3997 (
            .O(N__21265),
            .I(N__21255));
    Span12Mux_v I__3996 (
            .O(N__21262),
            .I(N__21252));
    Span4Mux_h I__3995 (
            .O(N__21259),
            .I(N__21249));
    InMux I__3994 (
            .O(N__21258),
            .I(N__21246));
    Span12Mux_v I__3993 (
            .O(N__21255),
            .I(N__21243));
    Odrv12 I__3992 (
            .O(N__21252),
            .I(rand_data_29));
    Odrv4 I__3991 (
            .O(N__21249),
            .I(rand_data_29));
    LocalMux I__3990 (
            .O(N__21246),
            .I(rand_data_29));
    Odrv12 I__3989 (
            .O(N__21243),
            .I(rand_data_29));
    InMux I__3988 (
            .O(N__21234),
            .I(N__21229));
    InMux I__3987 (
            .O(N__21233),
            .I(N__21226));
    InMux I__3986 (
            .O(N__21232),
            .I(N__21222));
    LocalMux I__3985 (
            .O(N__21229),
            .I(N__21219));
    LocalMux I__3984 (
            .O(N__21226),
            .I(N__21215));
    InMux I__3983 (
            .O(N__21225),
            .I(N__21212));
    LocalMux I__3982 (
            .O(N__21222),
            .I(N__21209));
    Span4Mux_h I__3981 (
            .O(N__21219),
            .I(N__21206));
    InMux I__3980 (
            .O(N__21218),
            .I(N__21203));
    Span4Mux_h I__3979 (
            .O(N__21215),
            .I(N__21200));
    LocalMux I__3978 (
            .O(N__21212),
            .I(N__21197));
    Span4Mux_s2_v I__3977 (
            .O(N__21209),
            .I(N__21192));
    Span4Mux_v I__3976 (
            .O(N__21206),
            .I(N__21192));
    LocalMux I__3975 (
            .O(N__21203),
            .I(data_in_field_109));
    Odrv4 I__3974 (
            .O(N__21200),
            .I(data_in_field_109));
    Odrv4 I__3973 (
            .O(N__21197),
            .I(data_in_field_109));
    Odrv4 I__3972 (
            .O(N__21192),
            .I(data_in_field_109));
    InMux I__3971 (
            .O(N__21183),
            .I(N__21176));
    InMux I__3970 (
            .O(N__21182),
            .I(N__21173));
    InMux I__3969 (
            .O(N__21181),
            .I(N__21168));
    InMux I__3968 (
            .O(N__21180),
            .I(N__21168));
    InMux I__3967 (
            .O(N__21179),
            .I(N__21165));
    LocalMux I__3966 (
            .O(N__21176),
            .I(rand_data_4));
    LocalMux I__3965 (
            .O(N__21173),
            .I(rand_data_4));
    LocalMux I__3964 (
            .O(N__21168),
            .I(rand_data_4));
    LocalMux I__3963 (
            .O(N__21165),
            .I(rand_data_4));
    InMux I__3962 (
            .O(N__21156),
            .I(N__21150));
    InMux I__3961 (
            .O(N__21155),
            .I(N__21145));
    InMux I__3960 (
            .O(N__21154),
            .I(N__21145));
    InMux I__3959 (
            .O(N__21153),
            .I(N__21141));
    LocalMux I__3958 (
            .O(N__21150),
            .I(N__21136));
    LocalMux I__3957 (
            .O(N__21145),
            .I(N__21136));
    InMux I__3956 (
            .O(N__21144),
            .I(N__21133));
    LocalMux I__3955 (
            .O(N__21141),
            .I(rand_data_3));
    Odrv12 I__3954 (
            .O(N__21136),
            .I(rand_data_3));
    LocalMux I__3953 (
            .O(N__21133),
            .I(rand_data_3));
    CascadeMux I__3952 (
            .O(N__21126),
            .I(N__21122));
    InMux I__3951 (
            .O(N__21125),
            .I(N__21119));
    InMux I__3950 (
            .O(N__21122),
            .I(N__21116));
    LocalMux I__3949 (
            .O(N__21119),
            .I(N__21113));
    LocalMux I__3948 (
            .O(N__21116),
            .I(N__21108));
    Span4Mux_v I__3947 (
            .O(N__21113),
            .I(N__21108));
    Odrv4 I__3946 (
            .O(N__21108),
            .I(\c0.n8992 ));
    InMux I__3945 (
            .O(N__21105),
            .I(N__21102));
    LocalMux I__3944 (
            .O(N__21102),
            .I(N__21099));
    Span4Mux_s2_h I__3943 (
            .O(N__21099),
            .I(N__21096));
    Span4Mux_h I__3942 (
            .O(N__21096),
            .I(N__21093));
    Odrv4 I__3941 (
            .O(N__21093),
            .I(\c0.n21_adj_1624 ));
    InMux I__3940 (
            .O(N__21090),
            .I(N__21086));
    InMux I__3939 (
            .O(N__21089),
            .I(N__21082));
    LocalMux I__3938 (
            .O(N__21086),
            .I(N__21079));
    InMux I__3937 (
            .O(N__21085),
            .I(N__21076));
    LocalMux I__3936 (
            .O(N__21082),
            .I(N__21072));
    Span4Mux_v I__3935 (
            .O(N__21079),
            .I(N__21067));
    LocalMux I__3934 (
            .O(N__21076),
            .I(N__21067));
    InMux I__3933 (
            .O(N__21075),
            .I(N__21064));
    Span12Mux_v I__3932 (
            .O(N__21072),
            .I(N__21060));
    Span4Mux_s3_h I__3931 (
            .O(N__21067),
            .I(N__21055));
    LocalMux I__3930 (
            .O(N__21064),
            .I(N__21055));
    InMux I__3929 (
            .O(N__21063),
            .I(N__21052));
    Odrv12 I__3928 (
            .O(N__21060),
            .I(rand_data_7));
    Odrv4 I__3927 (
            .O(N__21055),
            .I(rand_data_7));
    LocalMux I__3926 (
            .O(N__21052),
            .I(rand_data_7));
    CascadeMux I__3925 (
            .O(N__21045),
            .I(N__21041));
    CascadeMux I__3924 (
            .O(N__21044),
            .I(N__21037));
    InMux I__3923 (
            .O(N__21041),
            .I(N__21034));
    InMux I__3922 (
            .O(N__21040),
            .I(N__21031));
    InMux I__3921 (
            .O(N__21037),
            .I(N__21028));
    LocalMux I__3920 (
            .O(N__21034),
            .I(N__21023));
    LocalMux I__3919 (
            .O(N__21031),
            .I(N__21023));
    LocalMux I__3918 (
            .O(N__21028),
            .I(N__21020));
    Span4Mux_v I__3917 (
            .O(N__21023),
            .I(N__21015));
    Span4Mux_v I__3916 (
            .O(N__21020),
            .I(N__21012));
    InMux I__3915 (
            .O(N__21019),
            .I(N__21009));
    InMux I__3914 (
            .O(N__21018),
            .I(N__21006));
    Odrv4 I__3913 (
            .O(N__21015),
            .I(rand_data_1));
    Odrv4 I__3912 (
            .O(N__21012),
            .I(rand_data_1));
    LocalMux I__3911 (
            .O(N__21009),
            .I(rand_data_1));
    LocalMux I__3910 (
            .O(N__21006),
            .I(rand_data_1));
    InMux I__3909 (
            .O(N__20997),
            .I(\c0.n8116 ));
    InMux I__3908 (
            .O(N__20994),
            .I(N__20990));
    InMux I__3907 (
            .O(N__20993),
            .I(N__20987));
    LocalMux I__3906 (
            .O(N__20990),
            .I(\c0.byte_transmit_counter2_5 ));
    LocalMux I__3905 (
            .O(N__20987),
            .I(\c0.byte_transmit_counter2_5 ));
    InMux I__3904 (
            .O(N__20982),
            .I(\c0.n8117 ));
    InMux I__3903 (
            .O(N__20979),
            .I(N__20975));
    InMux I__3902 (
            .O(N__20978),
            .I(N__20972));
    LocalMux I__3901 (
            .O(N__20975),
            .I(\c0.byte_transmit_counter2_6 ));
    LocalMux I__3900 (
            .O(N__20972),
            .I(\c0.byte_transmit_counter2_6 ));
    InMux I__3899 (
            .O(N__20967),
            .I(\c0.n8118 ));
    InMux I__3898 (
            .O(N__20964),
            .I(\c0.n8119 ));
    CascadeMux I__3897 (
            .O(N__20961),
            .I(N__20957));
    InMux I__3896 (
            .O(N__20960),
            .I(N__20954));
    InMux I__3895 (
            .O(N__20957),
            .I(N__20951));
    LocalMux I__3894 (
            .O(N__20954),
            .I(\c0.byte_transmit_counter2_7 ));
    LocalMux I__3893 (
            .O(N__20951),
            .I(\c0.byte_transmit_counter2_7 ));
    CEMux I__3892 (
            .O(N__20946),
            .I(N__20943));
    LocalMux I__3891 (
            .O(N__20943),
            .I(N__20940));
    Span4Mux_h I__3890 (
            .O(N__20940),
            .I(N__20937));
    Odrv4 I__3889 (
            .O(N__20937),
            .I(\c0.n4897 ));
    SRMux I__3888 (
            .O(N__20934),
            .I(N__20931));
    LocalMux I__3887 (
            .O(N__20931),
            .I(N__20928));
    Span4Mux_h I__3886 (
            .O(N__20928),
            .I(N__20925));
    Odrv4 I__3885 (
            .O(N__20925),
            .I(\c0.n5154 ));
    InMux I__3884 (
            .O(N__20922),
            .I(N__20917));
    InMux I__3883 (
            .O(N__20921),
            .I(N__20913));
    InMux I__3882 (
            .O(N__20920),
            .I(N__20910));
    LocalMux I__3881 (
            .O(N__20917),
            .I(N__20907));
    InMux I__3880 (
            .O(N__20916),
            .I(N__20904));
    LocalMux I__3879 (
            .O(N__20913),
            .I(N__20900));
    LocalMux I__3878 (
            .O(N__20910),
            .I(N__20897));
    Span4Mux_h I__3877 (
            .O(N__20907),
            .I(N__20892));
    LocalMux I__3876 (
            .O(N__20904),
            .I(N__20892));
    InMux I__3875 (
            .O(N__20903),
            .I(N__20889));
    Odrv4 I__3874 (
            .O(N__20900),
            .I(rand_data_8));
    Odrv12 I__3873 (
            .O(N__20897),
            .I(rand_data_8));
    Odrv4 I__3872 (
            .O(N__20892),
            .I(rand_data_8));
    LocalMux I__3871 (
            .O(N__20889),
            .I(rand_data_8));
    InMux I__3870 (
            .O(N__20880),
            .I(N__20876));
    InMux I__3869 (
            .O(N__20879),
            .I(N__20872));
    LocalMux I__3868 (
            .O(N__20876),
            .I(N__20869));
    InMux I__3867 (
            .O(N__20875),
            .I(N__20866));
    LocalMux I__3866 (
            .O(N__20872),
            .I(N__20863));
    Span4Mux_v I__3865 (
            .O(N__20869),
            .I(N__20858));
    LocalMux I__3864 (
            .O(N__20866),
            .I(N__20858));
    Span4Mux_h I__3863 (
            .O(N__20863),
            .I(N__20855));
    Span4Mux_v I__3862 (
            .O(N__20858),
            .I(N__20852));
    Span4Mux_v I__3861 (
            .O(N__20855),
            .I(N__20849));
    Span4Mux_h I__3860 (
            .O(N__20852),
            .I(N__20845));
    Span4Mux_v I__3859 (
            .O(N__20849),
            .I(N__20842));
    InMux I__3858 (
            .O(N__20848),
            .I(N__20839));
    Odrv4 I__3857 (
            .O(N__20845),
            .I(rand_data_22));
    Odrv4 I__3856 (
            .O(N__20842),
            .I(rand_data_22));
    LocalMux I__3855 (
            .O(N__20839),
            .I(rand_data_22));
    CascadeMux I__3854 (
            .O(N__20832),
            .I(\c0.n7194_cascade_ ));
    InMux I__3853 (
            .O(N__20829),
            .I(N__20826));
    LocalMux I__3852 (
            .O(N__20826),
            .I(N__20823));
    Span4Mux_h I__3851 (
            .O(N__20823),
            .I(N__20819));
    InMux I__3850 (
            .O(N__20822),
            .I(N__20816));
    Span4Mux_s3_h I__3849 (
            .O(N__20819),
            .I(N__20811));
    LocalMux I__3848 (
            .O(N__20816),
            .I(N__20811));
    Odrv4 I__3847 (
            .O(N__20811),
            .I(\c0.n8449 ));
    CEMux I__3846 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__3845 (
            .O(N__20805),
            .I(N__20802));
    Span4Mux_v I__3844 (
            .O(N__20802),
            .I(N__20799));
    Span4Mux_h I__3843 (
            .O(N__20799),
            .I(N__20796));
    Odrv4 I__3842 (
            .O(N__20796),
            .I(n4839));
    CascadeMux I__3841 (
            .O(N__20793),
            .I(n4839_cascade_));
    InMux I__3840 (
            .O(N__20790),
            .I(N__20786));
    InMux I__3839 (
            .O(N__20789),
            .I(N__20783));
    LocalMux I__3838 (
            .O(N__20786),
            .I(N__20780));
    LocalMux I__3837 (
            .O(N__20783),
            .I(N__20777));
    Span4Mux_h I__3836 (
            .O(N__20780),
            .I(N__20771));
    Span4Mux_h I__3835 (
            .O(N__20777),
            .I(N__20768));
    InMux I__3834 (
            .O(N__20776),
            .I(N__20765));
    InMux I__3833 (
            .O(N__20775),
            .I(N__20760));
    InMux I__3832 (
            .O(N__20774),
            .I(N__20760));
    Odrv4 I__3831 (
            .O(N__20771),
            .I(n31));
    Odrv4 I__3830 (
            .O(N__20768),
            .I(n31));
    LocalMux I__3829 (
            .O(N__20765),
            .I(n31));
    LocalMux I__3828 (
            .O(N__20760),
            .I(n31));
    InMux I__3827 (
            .O(N__20751),
            .I(N__20746));
    CascadeMux I__3826 (
            .O(N__20750),
            .I(N__20743));
    CascadeMux I__3825 (
            .O(N__20749),
            .I(N__20740));
    LocalMux I__3824 (
            .O(N__20746),
            .I(N__20736));
    InMux I__3823 (
            .O(N__20743),
            .I(N__20733));
    InMux I__3822 (
            .O(N__20740),
            .I(N__20730));
    InMux I__3821 (
            .O(N__20739),
            .I(N__20727));
    Span4Mux_v I__3820 (
            .O(N__20736),
            .I(N__20724));
    LocalMux I__3819 (
            .O(N__20733),
            .I(N__20719));
    LocalMux I__3818 (
            .O(N__20730),
            .I(N__20719));
    LocalMux I__3817 (
            .O(N__20727),
            .I(N__20711));
    Span4Mux_h I__3816 (
            .O(N__20724),
            .I(N__20711));
    Span4Mux_v I__3815 (
            .O(N__20719),
            .I(N__20711));
    InMux I__3814 (
            .O(N__20718),
            .I(N__20708));
    Span4Mux_v I__3813 (
            .O(N__20711),
            .I(N__20705));
    LocalMux I__3812 (
            .O(N__20708),
            .I(data_in_field_65));
    Odrv4 I__3811 (
            .O(N__20705),
            .I(data_in_field_65));
    CascadeMux I__3810 (
            .O(N__20700),
            .I(N__20697));
    InMux I__3809 (
            .O(N__20697),
            .I(N__20693));
    InMux I__3808 (
            .O(N__20696),
            .I(N__20690));
    LocalMux I__3807 (
            .O(N__20693),
            .I(\c0.tx2_transmit_N_1444 ));
    LocalMux I__3806 (
            .O(N__20690),
            .I(\c0.tx2_transmit_N_1444 ));
    InMux I__3805 (
            .O(N__20685),
            .I(\c0.n8113 ));
    InMux I__3804 (
            .O(N__20682),
            .I(\c0.n8114 ));
    InMux I__3803 (
            .O(N__20679),
            .I(\c0.n8115 ));
    InMux I__3802 (
            .O(N__20676),
            .I(N__20672));
    InMux I__3801 (
            .O(N__20675),
            .I(N__20668));
    LocalMux I__3800 (
            .O(N__20672),
            .I(N__20665));
    InMux I__3799 (
            .O(N__20671),
            .I(N__20661));
    LocalMux I__3798 (
            .O(N__20668),
            .I(N__20658));
    Span4Mux_v I__3797 (
            .O(N__20665),
            .I(N__20655));
    InMux I__3796 (
            .O(N__20664),
            .I(N__20652));
    LocalMux I__3795 (
            .O(N__20661),
            .I(rand_data_24));
    Odrv4 I__3794 (
            .O(N__20658),
            .I(rand_data_24));
    Odrv4 I__3793 (
            .O(N__20655),
            .I(rand_data_24));
    LocalMux I__3792 (
            .O(N__20652),
            .I(rand_data_24));
    InMux I__3791 (
            .O(N__20643),
            .I(N__20640));
    LocalMux I__3790 (
            .O(N__20640),
            .I(N__20637));
    Span4Mux_h I__3789 (
            .O(N__20637),
            .I(N__20634));
    Odrv4 I__3788 (
            .O(N__20634),
            .I(n1903));
    InMux I__3787 (
            .O(N__20631),
            .I(N__20626));
    InMux I__3786 (
            .O(N__20630),
            .I(N__20623));
    InMux I__3785 (
            .O(N__20629),
            .I(N__20620));
    LocalMux I__3784 (
            .O(N__20626),
            .I(N__20617));
    LocalMux I__3783 (
            .O(N__20623),
            .I(N__20614));
    LocalMux I__3782 (
            .O(N__20620),
            .I(N__20609));
    Span4Mux_v I__3781 (
            .O(N__20617),
            .I(N__20609));
    Span4Mux_s3_h I__3780 (
            .O(N__20614),
            .I(N__20606));
    Span4Mux_v I__3779 (
            .O(N__20609),
            .I(N__20601));
    Span4Mux_h I__3778 (
            .O(N__20606),
            .I(N__20598));
    InMux I__3777 (
            .O(N__20605),
            .I(N__20593));
    InMux I__3776 (
            .O(N__20604),
            .I(N__20593));
    Span4Mux_h I__3775 (
            .O(N__20601),
            .I(N__20590));
    Odrv4 I__3774 (
            .O(N__20598),
            .I(data_in_field_129));
    LocalMux I__3773 (
            .O(N__20593),
            .I(data_in_field_129));
    Odrv4 I__3772 (
            .O(N__20590),
            .I(data_in_field_129));
    CascadeMux I__3771 (
            .O(N__20583),
            .I(N__20580));
    InMux I__3770 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__3769 (
            .O(N__20577),
            .I(N__20574));
    Span4Mux_v I__3768 (
            .O(N__20574),
            .I(N__20571));
    Span4Mux_h I__3767 (
            .O(N__20571),
            .I(N__20568));
    Span4Mux_v I__3766 (
            .O(N__20568),
            .I(N__20565));
    Odrv4 I__3765 (
            .O(N__20565),
            .I(\c0.n8791 ));
    InMux I__3764 (
            .O(N__20562),
            .I(N__20558));
    CascadeMux I__3763 (
            .O(N__20561),
            .I(N__20555));
    LocalMux I__3762 (
            .O(N__20558),
            .I(N__20552));
    InMux I__3761 (
            .O(N__20555),
            .I(N__20549));
    Span4Mux_v I__3760 (
            .O(N__20552),
            .I(N__20546));
    LocalMux I__3759 (
            .O(N__20549),
            .I(N__20542));
    Span4Mux_h I__3758 (
            .O(N__20546),
            .I(N__20539));
    InMux I__3757 (
            .O(N__20545),
            .I(N__20536));
    Span4Mux_v I__3756 (
            .O(N__20542),
            .I(N__20533));
    Odrv4 I__3755 (
            .O(N__20539),
            .I(data_in_6_0));
    LocalMux I__3754 (
            .O(N__20536),
            .I(data_in_6_0));
    Odrv4 I__3753 (
            .O(N__20533),
            .I(data_in_6_0));
    InMux I__3752 (
            .O(N__20526),
            .I(N__20523));
    LocalMux I__3751 (
            .O(N__20523),
            .I(N__20520));
    Span4Mux_h I__3750 (
            .O(N__20520),
            .I(N__20515));
    InMux I__3749 (
            .O(N__20519),
            .I(N__20510));
    InMux I__3748 (
            .O(N__20518),
            .I(N__20510));
    Odrv4 I__3747 (
            .O(N__20515),
            .I(data_in_5_0));
    LocalMux I__3746 (
            .O(N__20510),
            .I(data_in_5_0));
    CascadeMux I__3745 (
            .O(N__20505),
            .I(\c0.n19_adj_1665_cascade_ ));
    InMux I__3744 (
            .O(N__20502),
            .I(N__20496));
    InMux I__3743 (
            .O(N__20501),
            .I(N__20496));
    LocalMux I__3742 (
            .O(N__20496),
            .I(N__20492));
    CascadeMux I__3741 (
            .O(N__20495),
            .I(N__20489));
    Span4Mux_h I__3740 (
            .O(N__20492),
            .I(N__20486));
    InMux I__3739 (
            .O(N__20489),
            .I(N__20483));
    Span4Mux_v I__3738 (
            .O(N__20486),
            .I(N__20480));
    LocalMux I__3737 (
            .O(N__20483),
            .I(tx2_active));
    Odrv4 I__3736 (
            .O(N__20480),
            .I(tx2_active));
    InMux I__3735 (
            .O(N__20475),
            .I(N__20468));
    InMux I__3734 (
            .O(N__20474),
            .I(N__20468));
    InMux I__3733 (
            .O(N__20473),
            .I(N__20465));
    LocalMux I__3732 (
            .O(N__20468),
            .I(N__20460));
    LocalMux I__3731 (
            .O(N__20465),
            .I(N__20460));
    Span4Mux_v I__3730 (
            .O(N__20460),
            .I(N__20457));
    Span4Mux_h I__3729 (
            .O(N__20457),
            .I(N__20453));
    CascadeMux I__3728 (
            .O(N__20456),
            .I(N__20450));
    Span4Mux_v I__3727 (
            .O(N__20453),
            .I(N__20446));
    InMux I__3726 (
            .O(N__20450),
            .I(N__20441));
    InMux I__3725 (
            .O(N__20449),
            .I(N__20441));
    Odrv4 I__3724 (
            .O(N__20446),
            .I(\c0.r_SM_Main_2_N_1483_0 ));
    LocalMux I__3723 (
            .O(N__20441),
            .I(\c0.r_SM_Main_2_N_1483_0 ));
    InMux I__3722 (
            .O(N__20436),
            .I(N__20433));
    LocalMux I__3721 (
            .O(N__20433),
            .I(\c0.n19_adj_1665 ));
    InMux I__3720 (
            .O(N__20430),
            .I(N__20426));
    InMux I__3719 (
            .O(N__20429),
            .I(N__20423));
    LocalMux I__3718 (
            .O(N__20426),
            .I(rx_data_6));
    LocalMux I__3717 (
            .O(N__20423),
            .I(rx_data_6));
    InMux I__3716 (
            .O(N__20418),
            .I(N__20415));
    LocalMux I__3715 (
            .O(N__20415),
            .I(N__20411));
    CascadeMux I__3714 (
            .O(N__20414),
            .I(N__20408));
    Span4Mux_h I__3713 (
            .O(N__20411),
            .I(N__20405));
    InMux I__3712 (
            .O(N__20408),
            .I(N__20402));
    Odrv4 I__3711 (
            .O(N__20405),
            .I(rx_data_4));
    LocalMux I__3710 (
            .O(N__20402),
            .I(rx_data_4));
    InMux I__3709 (
            .O(N__20397),
            .I(N__20391));
    InMux I__3708 (
            .O(N__20396),
            .I(N__20391));
    LocalMux I__3707 (
            .O(N__20391),
            .I(rx_data_7));
    InMux I__3706 (
            .O(N__20388),
            .I(N__20382));
    InMux I__3705 (
            .O(N__20387),
            .I(N__20382));
    LocalMux I__3704 (
            .O(N__20382),
            .I(data_in_20_7));
    InMux I__3703 (
            .O(N__20379),
            .I(N__20375));
    InMux I__3702 (
            .O(N__20378),
            .I(N__20372));
    LocalMux I__3701 (
            .O(N__20375),
            .I(data_in_19_7));
    LocalMux I__3700 (
            .O(N__20372),
            .I(data_in_19_7));
    InMux I__3699 (
            .O(N__20367),
            .I(N__20362));
    InMux I__3698 (
            .O(N__20366),
            .I(N__20357));
    InMux I__3697 (
            .O(N__20365),
            .I(N__20357));
    LocalMux I__3696 (
            .O(N__20362),
            .I(n4044));
    LocalMux I__3695 (
            .O(N__20357),
            .I(n4044));
    CascadeMux I__3694 (
            .O(N__20352),
            .I(N__20348));
    InMux I__3693 (
            .O(N__20351),
            .I(N__20345));
    InMux I__3692 (
            .O(N__20348),
            .I(N__20342));
    LocalMux I__3691 (
            .O(N__20345),
            .I(rx_data_5));
    LocalMux I__3690 (
            .O(N__20342),
            .I(rx_data_5));
    InMux I__3689 (
            .O(N__20337),
            .I(N__20331));
    InMux I__3688 (
            .O(N__20336),
            .I(N__20328));
    InMux I__3687 (
            .O(N__20335),
            .I(N__20323));
    InMux I__3686 (
            .O(N__20334),
            .I(N__20323));
    LocalMux I__3685 (
            .O(N__20331),
            .I(N__20320));
    LocalMux I__3684 (
            .O(N__20328),
            .I(N__20317));
    LocalMux I__3683 (
            .O(N__20323),
            .I(n4049));
    Odrv4 I__3682 (
            .O(N__20320),
            .I(n4049));
    Odrv4 I__3681 (
            .O(N__20317),
            .I(n4049));
    CascadeMux I__3680 (
            .O(N__20310),
            .I(N__20307));
    InMux I__3679 (
            .O(N__20307),
            .I(N__20304));
    LocalMux I__3678 (
            .O(N__20304),
            .I(N__20301));
    Span4Mux_s2_h I__3677 (
            .O(N__20301),
            .I(N__20298));
    Span4Mux_h I__3676 (
            .O(N__20298),
            .I(N__20295));
    Span4Mux_v I__3675 (
            .O(N__20295),
            .I(N__20292));
    Odrv4 I__3674 (
            .O(N__20292),
            .I(\c0.n9476 ));
    CascadeMux I__3673 (
            .O(N__20289),
            .I(N__20286));
    InMux I__3672 (
            .O(N__20286),
            .I(N__20283));
    LocalMux I__3671 (
            .O(N__20283),
            .I(N__20279));
    InMux I__3670 (
            .O(N__20282),
            .I(N__20276));
    Odrv4 I__3669 (
            .O(N__20279),
            .I(n4));
    LocalMux I__3668 (
            .O(N__20276),
            .I(n4));
    InMux I__3667 (
            .O(N__20271),
            .I(N__20267));
    InMux I__3666 (
            .O(N__20270),
            .I(N__20264));
    LocalMux I__3665 (
            .O(N__20267),
            .I(rx_data_3));
    LocalMux I__3664 (
            .O(N__20264),
            .I(rx_data_3));
    InMux I__3663 (
            .O(N__20259),
            .I(N__20255));
    InMux I__3662 (
            .O(N__20258),
            .I(N__20252));
    LocalMux I__3661 (
            .O(N__20255),
            .I(data_in_19_6));
    LocalMux I__3660 (
            .O(N__20252),
            .I(data_in_19_6));
    InMux I__3659 (
            .O(N__20247),
            .I(N__20243));
    CascadeMux I__3658 (
            .O(N__20246),
            .I(N__20240));
    LocalMux I__3657 (
            .O(N__20243),
            .I(N__20237));
    InMux I__3656 (
            .O(N__20240),
            .I(N__20234));
    Span4Mux_v I__3655 (
            .O(N__20237),
            .I(N__20231));
    LocalMux I__3654 (
            .O(N__20234),
            .I(rx_data_0));
    Odrv4 I__3653 (
            .O(N__20231),
            .I(rx_data_0));
    InMux I__3652 (
            .O(N__20226),
            .I(N__20223));
    LocalMux I__3651 (
            .O(N__20223),
            .I(N__20220));
    Span4Mux_h I__3650 (
            .O(N__20220),
            .I(N__20216));
    InMux I__3649 (
            .O(N__20219),
            .I(N__20213));
    Odrv4 I__3648 (
            .O(N__20216),
            .I(data_in_18_7));
    LocalMux I__3647 (
            .O(N__20213),
            .I(data_in_18_7));
    InMux I__3646 (
            .O(N__20208),
            .I(N__20202));
    InMux I__3645 (
            .O(N__20207),
            .I(N__20202));
    LocalMux I__3644 (
            .O(N__20202),
            .I(data_in_20_6));
    InMux I__3643 (
            .O(N__20199),
            .I(N__20196));
    LocalMux I__3642 (
            .O(N__20196),
            .I(n4_adj_1725));
    CascadeMux I__3641 (
            .O(N__20193),
            .I(n4_adj_1725_cascade_));
    InMux I__3640 (
            .O(N__20190),
            .I(N__20186));
    InMux I__3639 (
            .O(N__20189),
            .I(N__20183));
    LocalMux I__3638 (
            .O(N__20186),
            .I(rx_data_1));
    LocalMux I__3637 (
            .O(N__20183),
            .I(rx_data_1));
    CascadeMux I__3636 (
            .O(N__20178),
            .I(n4044_cascade_));
    InMux I__3635 (
            .O(N__20175),
            .I(N__20169));
    InMux I__3634 (
            .O(N__20174),
            .I(N__20169));
    LocalMux I__3633 (
            .O(N__20169),
            .I(data_in_16_5));
    InMux I__3632 (
            .O(N__20166),
            .I(N__20162));
    InMux I__3631 (
            .O(N__20165),
            .I(N__20159));
    LocalMux I__3630 (
            .O(N__20162),
            .I(data_in_18_5));
    LocalMux I__3629 (
            .O(N__20159),
            .I(data_in_18_5));
    InMux I__3628 (
            .O(N__20154),
            .I(N__20148));
    InMux I__3627 (
            .O(N__20153),
            .I(N__20148));
    LocalMux I__3626 (
            .O(N__20148),
            .I(data_in_17_5));
    InMux I__3625 (
            .O(N__20145),
            .I(N__20141));
    InMux I__3624 (
            .O(N__20144),
            .I(N__20138));
    LocalMux I__3623 (
            .O(N__20141),
            .I(data_in_18_6));
    LocalMux I__3622 (
            .O(N__20138),
            .I(data_in_18_6));
    InMux I__3621 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__3620 (
            .O(N__20130),
            .I(N__20127));
    Span4Mux_h I__3619 (
            .O(N__20127),
            .I(N__20123));
    InMux I__3618 (
            .O(N__20126),
            .I(N__20120));
    Odrv4 I__3617 (
            .O(N__20123),
            .I(data_in_18_1));
    LocalMux I__3616 (
            .O(N__20120),
            .I(data_in_18_1));
    InMux I__3615 (
            .O(N__20115),
            .I(N__20109));
    InMux I__3614 (
            .O(N__20114),
            .I(N__20109));
    LocalMux I__3613 (
            .O(N__20109),
            .I(data_in_19_1));
    InMux I__3612 (
            .O(N__20106),
            .I(N__20100));
    InMux I__3611 (
            .O(N__20105),
            .I(N__20100));
    LocalMux I__3610 (
            .O(N__20100),
            .I(data_in_20_1));
    CascadeMux I__3609 (
            .O(N__20097),
            .I(N__20094));
    InMux I__3608 (
            .O(N__20094),
            .I(N__20088));
    InMux I__3607 (
            .O(N__20093),
            .I(N__20088));
    LocalMux I__3606 (
            .O(N__20088),
            .I(rx_data_2));
    InMux I__3605 (
            .O(N__20085),
            .I(N__20082));
    LocalMux I__3604 (
            .O(N__20082),
            .I(N__20078));
    InMux I__3603 (
            .O(N__20081),
            .I(N__20075));
    Odrv4 I__3602 (
            .O(N__20078),
            .I(data_in_12_3));
    LocalMux I__3601 (
            .O(N__20075),
            .I(data_in_12_3));
    InMux I__3600 (
            .O(N__20070),
            .I(N__20067));
    LocalMux I__3599 (
            .O(N__20067),
            .I(N__20063));
    InMux I__3598 (
            .O(N__20066),
            .I(N__20060));
    Odrv4 I__3597 (
            .O(N__20063),
            .I(data_in_11_3));
    LocalMux I__3596 (
            .O(N__20060),
            .I(data_in_11_3));
    CascadeMux I__3595 (
            .O(N__20055),
            .I(\c0.n9590_cascade_ ));
    InMux I__3594 (
            .O(N__20052),
            .I(N__20049));
    LocalMux I__3593 (
            .O(N__20049),
            .I(\c0.n9153 ));
    CascadeMux I__3592 (
            .O(N__20046),
            .I(\c0.n9156_cascade_ ));
    CascadeMux I__3591 (
            .O(N__20043),
            .I(\c0.n9584_cascade_ ));
    InMux I__3590 (
            .O(N__20040),
            .I(N__20037));
    LocalMux I__3589 (
            .O(N__20037),
            .I(N__20034));
    Span12Mux_s3_v I__3588 (
            .O(N__20034),
            .I(N__20031));
    Odrv12 I__3587 (
            .O(N__20031),
            .I(\c0.n9150 ));
    InMux I__3586 (
            .O(N__20028),
            .I(N__20025));
    LocalMux I__3585 (
            .O(N__20025),
            .I(N__20022));
    Span4Mux_v I__3584 (
            .O(N__20022),
            .I(N__20019));
    Span4Mux_h I__3583 (
            .O(N__20019),
            .I(N__20016));
    Odrv4 I__3582 (
            .O(N__20016),
            .I(\c0.n22_adj_1678 ));
    CascadeMux I__3581 (
            .O(N__20013),
            .I(\c0.n9587_cascade_ ));
    InMux I__3580 (
            .O(N__20010),
            .I(N__20007));
    LocalMux I__3579 (
            .O(N__20007),
            .I(N__20004));
    Odrv4 I__3578 (
            .O(N__20004),
            .I(\c0.tx2.r_Tx_Data_5 ));
    InMux I__3577 (
            .O(N__20001),
            .I(N__19998));
    LocalMux I__3576 (
            .O(N__19998),
            .I(N__19995));
    Span4Mux_v I__3575 (
            .O(N__19995),
            .I(N__19991));
    InMux I__3574 (
            .O(N__19994),
            .I(N__19988));
    Odrv4 I__3573 (
            .O(N__19991),
            .I(data_in_10_5));
    LocalMux I__3572 (
            .O(N__19988),
            .I(data_in_10_5));
    InMux I__3571 (
            .O(N__19983),
            .I(N__19977));
    InMux I__3570 (
            .O(N__19982),
            .I(N__19977));
    LocalMux I__3569 (
            .O(N__19977),
            .I(data_in_11_5));
    InMux I__3568 (
            .O(N__19974),
            .I(N__19970));
    InMux I__3567 (
            .O(N__19973),
            .I(N__19967));
    LocalMux I__3566 (
            .O(N__19970),
            .I(data_in_13_5));
    LocalMux I__3565 (
            .O(N__19967),
            .I(data_in_13_5));
    InMux I__3564 (
            .O(N__19962),
            .I(N__19956));
    InMux I__3563 (
            .O(N__19961),
            .I(N__19956));
    LocalMux I__3562 (
            .O(N__19956),
            .I(data_in_12_5));
    InMux I__3561 (
            .O(N__19953),
            .I(N__19949));
    InMux I__3560 (
            .O(N__19952),
            .I(N__19946));
    LocalMux I__3559 (
            .O(N__19949),
            .I(data_in_14_5));
    LocalMux I__3558 (
            .O(N__19946),
            .I(data_in_14_5));
    InMux I__3557 (
            .O(N__19941),
            .I(N__19935));
    InMux I__3556 (
            .O(N__19940),
            .I(N__19935));
    LocalMux I__3555 (
            .O(N__19935),
            .I(data_in_15_5));
    InMux I__3554 (
            .O(N__19932),
            .I(N__19929));
    LocalMux I__3553 (
            .O(N__19929),
            .I(N__19924));
    InMux I__3552 (
            .O(N__19928),
            .I(N__19921));
    InMux I__3551 (
            .O(N__19927),
            .I(N__19917));
    Span4Mux_v I__3550 (
            .O(N__19924),
            .I(N__19914));
    LocalMux I__3549 (
            .O(N__19921),
            .I(N__19911));
    InMux I__3548 (
            .O(N__19920),
            .I(N__19907));
    LocalMux I__3547 (
            .O(N__19917),
            .I(N__19902));
    Span4Mux_h I__3546 (
            .O(N__19914),
            .I(N__19902));
    Span4Mux_s2_v I__3545 (
            .O(N__19911),
            .I(N__19899));
    InMux I__3544 (
            .O(N__19910),
            .I(N__19896));
    LocalMux I__3543 (
            .O(N__19907),
            .I(data_in_field_141));
    Odrv4 I__3542 (
            .O(N__19902),
            .I(data_in_field_141));
    Odrv4 I__3541 (
            .O(N__19899),
            .I(data_in_field_141));
    LocalMux I__3540 (
            .O(N__19896),
            .I(data_in_field_141));
    InMux I__3539 (
            .O(N__19887),
            .I(N__19883));
    InMux I__3538 (
            .O(N__19886),
            .I(N__19879));
    LocalMux I__3537 (
            .O(N__19883),
            .I(N__19876));
    InMux I__3536 (
            .O(N__19882),
            .I(N__19872));
    LocalMux I__3535 (
            .O(N__19879),
            .I(N__19867));
    Span12Mux_v I__3534 (
            .O(N__19876),
            .I(N__19867));
    InMux I__3533 (
            .O(N__19875),
            .I(N__19864));
    LocalMux I__3532 (
            .O(N__19872),
            .I(rand_data_21));
    Odrv12 I__3531 (
            .O(N__19867),
            .I(rand_data_21));
    LocalMux I__3530 (
            .O(N__19864),
            .I(rand_data_21));
    InMux I__3529 (
            .O(N__19857),
            .I(N__19853));
    InMux I__3528 (
            .O(N__19856),
            .I(N__19849));
    LocalMux I__3527 (
            .O(N__19853),
            .I(N__19846));
    InMux I__3526 (
            .O(N__19852),
            .I(N__19843));
    LocalMux I__3525 (
            .O(N__19849),
            .I(N__19840));
    Span4Mux_h I__3524 (
            .O(N__19846),
            .I(N__19836));
    LocalMux I__3523 (
            .O(N__19843),
            .I(N__19833));
    Span12Mux_v I__3522 (
            .O(N__19840),
            .I(N__19830));
    InMux I__3521 (
            .O(N__19839),
            .I(N__19827));
    Odrv4 I__3520 (
            .O(N__19836),
            .I(rand_data_17));
    Odrv12 I__3519 (
            .O(N__19833),
            .I(rand_data_17));
    Odrv12 I__3518 (
            .O(N__19830),
            .I(rand_data_17));
    LocalMux I__3517 (
            .O(N__19827),
            .I(rand_data_17));
    CascadeMux I__3516 (
            .O(N__19818),
            .I(N__19814));
    InMux I__3515 (
            .O(N__19817),
            .I(N__19811));
    InMux I__3514 (
            .O(N__19814),
            .I(N__19808));
    LocalMux I__3513 (
            .O(N__19811),
            .I(N__19805));
    LocalMux I__3512 (
            .O(N__19808),
            .I(N__19802));
    Span4Mux_v I__3511 (
            .O(N__19805),
            .I(N__19795));
    Span4Mux_s2_h I__3510 (
            .O(N__19802),
            .I(N__19795));
    InMux I__3509 (
            .O(N__19801),
            .I(N__19790));
    InMux I__3508 (
            .O(N__19800),
            .I(N__19790));
    Span4Mux_h I__3507 (
            .O(N__19795),
            .I(N__19787));
    LocalMux I__3506 (
            .O(N__19790),
            .I(data_in_field_113));
    Odrv4 I__3505 (
            .O(N__19787),
            .I(data_in_field_113));
    CascadeMux I__3504 (
            .O(N__19782),
            .I(N__19778));
    InMux I__3503 (
            .O(N__19781),
            .I(N__19775));
    InMux I__3502 (
            .O(N__19778),
            .I(N__19772));
    LocalMux I__3501 (
            .O(N__19775),
            .I(N__19766));
    LocalMux I__3500 (
            .O(N__19772),
            .I(N__19763));
    InMux I__3499 (
            .O(N__19771),
            .I(N__19760));
    InMux I__3498 (
            .O(N__19770),
            .I(N__19757));
    InMux I__3497 (
            .O(N__19769),
            .I(N__19754));
    Sp12to4 I__3496 (
            .O(N__19766),
            .I(N__19747));
    Sp12to4 I__3495 (
            .O(N__19763),
            .I(N__19747));
    LocalMux I__3494 (
            .O(N__19760),
            .I(N__19747));
    LocalMux I__3493 (
            .O(N__19757),
            .I(N__19744));
    LocalMux I__3492 (
            .O(N__19754),
            .I(data_in_field_149));
    Odrv12 I__3491 (
            .O(N__19747),
            .I(data_in_field_149));
    Odrv12 I__3490 (
            .O(N__19744),
            .I(data_in_field_149));
    CascadeMux I__3489 (
            .O(N__19737),
            .I(N__19734));
    InMux I__3488 (
            .O(N__19734),
            .I(N__19731));
    LocalMux I__3487 (
            .O(N__19731),
            .I(N__19728));
    Span4Mux_v I__3486 (
            .O(N__19728),
            .I(N__19725));
    Odrv4 I__3485 (
            .O(N__19725),
            .I(\c0.n1893_adj_1635 ));
    InMux I__3484 (
            .O(N__19722),
            .I(N__19719));
    LocalMux I__3483 (
            .O(N__19719),
            .I(N__19716));
    Span4Mux_h I__3482 (
            .O(N__19716),
            .I(N__19711));
    InMux I__3481 (
            .O(N__19715),
            .I(N__19708));
    InMux I__3480 (
            .O(N__19714),
            .I(N__19705));
    Sp12to4 I__3479 (
            .O(N__19711),
            .I(N__19699));
    LocalMux I__3478 (
            .O(N__19708),
            .I(N__19699));
    LocalMux I__3477 (
            .O(N__19705),
            .I(N__19696));
    InMux I__3476 (
            .O(N__19704),
            .I(N__19693));
    Odrv12 I__3475 (
            .O(N__19699),
            .I(rand_data_23));
    Odrv12 I__3474 (
            .O(N__19696),
            .I(rand_data_23));
    LocalMux I__3473 (
            .O(N__19693),
            .I(rand_data_23));
    InMux I__3472 (
            .O(N__19686),
            .I(N__19681));
    InMux I__3471 (
            .O(N__19685),
            .I(N__19678));
    InMux I__3470 (
            .O(N__19684),
            .I(N__19673));
    LocalMux I__3469 (
            .O(N__19681),
            .I(N__19670));
    LocalMux I__3468 (
            .O(N__19678),
            .I(N__19667));
    InMux I__3467 (
            .O(N__19677),
            .I(N__19664));
    InMux I__3466 (
            .O(N__19676),
            .I(N__19661));
    LocalMux I__3465 (
            .O(N__19673),
            .I(N__19658));
    Span4Mux_h I__3464 (
            .O(N__19670),
            .I(N__19655));
    Span4Mux_s1_v I__3463 (
            .O(N__19667),
            .I(N__19650));
    LocalMux I__3462 (
            .O(N__19664),
            .I(N__19650));
    LocalMux I__3461 (
            .O(N__19661),
            .I(N__19645));
    Span4Mux_v I__3460 (
            .O(N__19658),
            .I(N__19645));
    Odrv4 I__3459 (
            .O(N__19655),
            .I(data_in_field_85));
    Odrv4 I__3458 (
            .O(N__19650),
            .I(data_in_field_85));
    Odrv4 I__3457 (
            .O(N__19645),
            .I(data_in_field_85));
    CascadeMux I__3456 (
            .O(N__19638),
            .I(\c0.n9596_cascade_ ));
    InMux I__3455 (
            .O(N__19635),
            .I(N__19632));
    LocalMux I__3454 (
            .O(N__19632),
            .I(N__19628));
    InMux I__3453 (
            .O(N__19631),
            .I(N__19624));
    Span4Mux_h I__3452 (
            .O(N__19628),
            .I(N__19621));
    InMux I__3451 (
            .O(N__19627),
            .I(N__19618));
    LocalMux I__3450 (
            .O(N__19624),
            .I(data_in_field_117));
    Odrv4 I__3449 (
            .O(N__19621),
            .I(data_in_field_117));
    LocalMux I__3448 (
            .O(N__19618),
            .I(data_in_field_117));
    CascadeMux I__3447 (
            .O(N__19611),
            .I(N__19607));
    InMux I__3446 (
            .O(N__19610),
            .I(N__19602));
    InMux I__3445 (
            .O(N__19607),
            .I(N__19602));
    LocalMux I__3444 (
            .O(N__19602),
            .I(N__19598));
    InMux I__3443 (
            .O(N__19601),
            .I(N__19595));
    Span4Mux_v I__3442 (
            .O(N__19598),
            .I(N__19592));
    LocalMux I__3441 (
            .O(N__19595),
            .I(N__19589));
    Span4Mux_s2_v I__3440 (
            .O(N__19592),
            .I(N__19585));
    Span12Mux_v I__3439 (
            .O(N__19589),
            .I(N__19582));
    InMux I__3438 (
            .O(N__19588),
            .I(N__19579));
    Odrv4 I__3437 (
            .O(N__19585),
            .I(rand_data_25));
    Odrv12 I__3436 (
            .O(N__19582),
            .I(rand_data_25));
    LocalMux I__3435 (
            .O(N__19579),
            .I(rand_data_25));
    InMux I__3434 (
            .O(N__19572),
            .I(n8179));
    InMux I__3433 (
            .O(N__19569),
            .I(n8180));
    InMux I__3432 (
            .O(N__19566),
            .I(N__19562));
    InMux I__3431 (
            .O(N__19565),
            .I(N__19559));
    LocalMux I__3430 (
            .O(N__19562),
            .I(N__19556));
    LocalMux I__3429 (
            .O(N__19559),
            .I(N__19553));
    Span4Mux_v I__3428 (
            .O(N__19556),
            .I(N__19549));
    Span4Mux_v I__3427 (
            .O(N__19553),
            .I(N__19546));
    InMux I__3426 (
            .O(N__19552),
            .I(N__19543));
    Sp12to4 I__3425 (
            .O(N__19549),
            .I(N__19540));
    Span4Mux_h I__3424 (
            .O(N__19546),
            .I(N__19534));
    LocalMux I__3423 (
            .O(N__19543),
            .I(N__19534));
    Span12Mux_s5_h I__3422 (
            .O(N__19540),
            .I(N__19531));
    InMux I__3421 (
            .O(N__19539),
            .I(N__19528));
    Odrv4 I__3420 (
            .O(N__19534),
            .I(rand_data_27));
    Odrv12 I__3419 (
            .O(N__19531),
            .I(rand_data_27));
    LocalMux I__3418 (
            .O(N__19528),
            .I(rand_data_27));
    InMux I__3417 (
            .O(N__19521),
            .I(n8181));
    InMux I__3416 (
            .O(N__19518),
            .I(n8182));
    InMux I__3415 (
            .O(N__19515),
            .I(n8183));
    InMux I__3414 (
            .O(N__19512),
            .I(n8184));
    InMux I__3413 (
            .O(N__19509),
            .I(n8185));
    InMux I__3412 (
            .O(N__19506),
            .I(N__19503));
    LocalMux I__3411 (
            .O(N__19503),
            .I(N__19497));
    InMux I__3410 (
            .O(N__19502),
            .I(N__19494));
    InMux I__3409 (
            .O(N__19501),
            .I(N__19489));
    InMux I__3408 (
            .O(N__19500),
            .I(N__19489));
    Span4Mux_v I__3407 (
            .O(N__19497),
            .I(N__19486));
    LocalMux I__3406 (
            .O(N__19494),
            .I(rand_data_31));
    LocalMux I__3405 (
            .O(N__19489),
            .I(rand_data_31));
    Odrv4 I__3404 (
            .O(N__19486),
            .I(rand_data_31));
    InMux I__3403 (
            .O(N__19479),
            .I(N__19476));
    LocalMux I__3402 (
            .O(N__19476),
            .I(N__19470));
    InMux I__3401 (
            .O(N__19475),
            .I(N__19467));
    InMux I__3400 (
            .O(N__19474),
            .I(N__19462));
    InMux I__3399 (
            .O(N__19473),
            .I(N__19462));
    Span4Mux_s2_v I__3398 (
            .O(N__19470),
            .I(N__19459));
    LocalMux I__3397 (
            .O(N__19467),
            .I(data_in_field_104));
    LocalMux I__3396 (
            .O(N__19462),
            .I(data_in_field_104));
    Odrv4 I__3395 (
            .O(N__19459),
            .I(data_in_field_104));
    CascadeMux I__3394 (
            .O(N__19452),
            .I(\c0.n9734_cascade_ ));
    InMux I__3393 (
            .O(N__19449),
            .I(bfn_6_29_0_));
    InMux I__3392 (
            .O(N__19446),
            .I(n8171));
    InMux I__3391 (
            .O(N__19443),
            .I(n8172));
    InMux I__3390 (
            .O(N__19440),
            .I(N__19435));
    InMux I__3389 (
            .O(N__19439),
            .I(N__19432));
    InMux I__3388 (
            .O(N__19438),
            .I(N__19429));
    LocalMux I__3387 (
            .O(N__19435),
            .I(N__19424));
    LocalMux I__3386 (
            .O(N__19432),
            .I(N__19424));
    LocalMux I__3385 (
            .O(N__19429),
            .I(N__19421));
    Span4Mux_h I__3384 (
            .O(N__19424),
            .I(N__19417));
    Span12Mux_s5_h I__3383 (
            .O(N__19421),
            .I(N__19414));
    InMux I__3382 (
            .O(N__19420),
            .I(N__19411));
    Odrv4 I__3381 (
            .O(N__19417),
            .I(rand_data_19));
    Odrv12 I__3380 (
            .O(N__19414),
            .I(rand_data_19));
    LocalMux I__3379 (
            .O(N__19411),
            .I(rand_data_19));
    InMux I__3378 (
            .O(N__19404),
            .I(n8173));
    InMux I__3377 (
            .O(N__19401),
            .I(n8174));
    InMux I__3376 (
            .O(N__19398),
            .I(n8175));
    InMux I__3375 (
            .O(N__19395),
            .I(n8176));
    InMux I__3374 (
            .O(N__19392),
            .I(n8177));
    InMux I__3373 (
            .O(N__19389),
            .I(bfn_6_30_0_));
    InMux I__3372 (
            .O(N__19386),
            .I(n8161));
    InMux I__3371 (
            .O(N__19383),
            .I(bfn_6_28_0_));
    InMux I__3370 (
            .O(N__19380),
            .I(n8163));
    InMux I__3369 (
            .O(N__19377),
            .I(n8164));
    InMux I__3368 (
            .O(N__19374),
            .I(n8165));
    InMux I__3367 (
            .O(N__19371),
            .I(n8166));
    InMux I__3366 (
            .O(N__19368),
            .I(n8167));
    InMux I__3365 (
            .O(N__19365),
            .I(N__19362));
    LocalMux I__3364 (
            .O(N__19362),
            .I(N__19358));
    InMux I__3363 (
            .O(N__19361),
            .I(N__19355));
    Sp12to4 I__3362 (
            .O(N__19358),
            .I(N__19347));
    LocalMux I__3361 (
            .O(N__19355),
            .I(N__19347));
    InMux I__3360 (
            .O(N__19354),
            .I(N__19344));
    InMux I__3359 (
            .O(N__19353),
            .I(N__19341));
    InMux I__3358 (
            .O(N__19352),
            .I(N__19338));
    Odrv12 I__3357 (
            .O(N__19347),
            .I(rand_data_14));
    LocalMux I__3356 (
            .O(N__19344),
            .I(rand_data_14));
    LocalMux I__3355 (
            .O(N__19341),
            .I(rand_data_14));
    LocalMux I__3354 (
            .O(N__19338),
            .I(rand_data_14));
    InMux I__3353 (
            .O(N__19329),
            .I(n8168));
    InMux I__3352 (
            .O(N__19326),
            .I(n8169));
    CascadeMux I__3351 (
            .O(N__19323),
            .I(\c0.n4897_cascade_ ));
    InMux I__3350 (
            .O(N__19320),
            .I(bfn_6_27_0_));
    InMux I__3349 (
            .O(N__19317),
            .I(n8155));
    InMux I__3348 (
            .O(N__19314),
            .I(n8156));
    InMux I__3347 (
            .O(N__19311),
            .I(n8157));
    InMux I__3346 (
            .O(N__19308),
            .I(n8158));
    InMux I__3345 (
            .O(N__19305),
            .I(N__19300));
    InMux I__3344 (
            .O(N__19304),
            .I(N__19296));
    InMux I__3343 (
            .O(N__19303),
            .I(N__19293));
    LocalMux I__3342 (
            .O(N__19300),
            .I(N__19290));
    InMux I__3341 (
            .O(N__19299),
            .I(N__19287));
    LocalMux I__3340 (
            .O(N__19296),
            .I(N__19284));
    LocalMux I__3339 (
            .O(N__19293),
            .I(N__19281));
    Span4Mux_v I__3338 (
            .O(N__19290),
            .I(N__19278));
    LocalMux I__3337 (
            .O(N__19287),
            .I(N__19273));
    Sp12to4 I__3336 (
            .O(N__19284),
            .I(N__19273));
    Span12Mux_s4_h I__3335 (
            .O(N__19281),
            .I(N__19265));
    Sp12to4 I__3334 (
            .O(N__19278),
            .I(N__19265));
    Span12Mux_s5_v I__3333 (
            .O(N__19273),
            .I(N__19265));
    InMux I__3332 (
            .O(N__19272),
            .I(N__19262));
    Odrv12 I__3331 (
            .O(N__19265),
            .I(rand_data_5));
    LocalMux I__3330 (
            .O(N__19262),
            .I(rand_data_5));
    InMux I__3329 (
            .O(N__19257),
            .I(n8159));
    InMux I__3328 (
            .O(N__19254),
            .I(n8160));
    InMux I__3327 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__3326 (
            .O(N__19248),
            .I(n9091));
    CascadeMux I__3325 (
            .O(N__19245),
            .I(n9092_cascade_));
    IoInMux I__3324 (
            .O(N__19242),
            .I(N__19239));
    LocalMux I__3323 (
            .O(N__19239),
            .I(N__19236));
    Span4Mux_s2_v I__3322 (
            .O(N__19236),
            .I(N__19233));
    Span4Mux_v I__3321 (
            .O(N__19233),
            .I(N__19230));
    Odrv4 I__3320 (
            .O(N__19230),
            .I(LED_c));
    SRMux I__3319 (
            .O(N__19227),
            .I(N__19224));
    LocalMux I__3318 (
            .O(N__19224),
            .I(N__19221));
    Span12Mux_v I__3317 (
            .O(N__19221),
            .I(N__19218));
    Odrv12 I__3316 (
            .O(N__19218),
            .I(n8761));
    CascadeMux I__3315 (
            .O(N__19215),
            .I(N__19210));
    InMux I__3314 (
            .O(N__19214),
            .I(N__19207));
    InMux I__3313 (
            .O(N__19213),
            .I(N__19203));
    InMux I__3312 (
            .O(N__19210),
            .I(N__19200));
    LocalMux I__3311 (
            .O(N__19207),
            .I(N__19197));
    InMux I__3310 (
            .O(N__19206),
            .I(N__19194));
    LocalMux I__3309 (
            .O(N__19203),
            .I(data_in_field_48));
    LocalMux I__3308 (
            .O(N__19200),
            .I(data_in_field_48));
    Odrv4 I__3307 (
            .O(N__19197),
            .I(data_in_field_48));
    LocalMux I__3306 (
            .O(N__19194),
            .I(data_in_field_48));
    InMux I__3305 (
            .O(N__19185),
            .I(N__19182));
    LocalMux I__3304 (
            .O(N__19182),
            .I(N__19176));
    InMux I__3303 (
            .O(N__19181),
            .I(N__19173));
    InMux I__3302 (
            .O(N__19180),
            .I(N__19168));
    InMux I__3301 (
            .O(N__19179),
            .I(N__19168));
    Span4Mux_h I__3300 (
            .O(N__19176),
            .I(N__19165));
    LocalMux I__3299 (
            .O(N__19173),
            .I(data_in_1_4));
    LocalMux I__3298 (
            .O(N__19168),
            .I(data_in_1_4));
    Odrv4 I__3297 (
            .O(N__19165),
            .I(data_in_1_4));
    CascadeMux I__3296 (
            .O(N__19158),
            .I(N__19155));
    InMux I__3295 (
            .O(N__19155),
            .I(N__19143));
    InMux I__3294 (
            .O(N__19154),
            .I(N__19138));
    InMux I__3293 (
            .O(N__19153),
            .I(N__19138));
    CascadeMux I__3292 (
            .O(N__19152),
            .I(N__19135));
    CascadeMux I__3291 (
            .O(N__19151),
            .I(N__19121));
    InMux I__3290 (
            .O(N__19150),
            .I(N__19114));
    InMux I__3289 (
            .O(N__19149),
            .I(N__19109));
    InMux I__3288 (
            .O(N__19148),
            .I(N__19105));
    InMux I__3287 (
            .O(N__19147),
            .I(N__19102));
    InMux I__3286 (
            .O(N__19146),
            .I(N__19099));
    LocalMux I__3285 (
            .O(N__19143),
            .I(N__19096));
    LocalMux I__3284 (
            .O(N__19138),
            .I(N__19093));
    InMux I__3283 (
            .O(N__19135),
            .I(N__19090));
    CascadeMux I__3282 (
            .O(N__19134),
            .I(N__19081));
    CascadeMux I__3281 (
            .O(N__19133),
            .I(N__19078));
    CascadeMux I__3280 (
            .O(N__19132),
            .I(N__19075));
    CascadeMux I__3279 (
            .O(N__19131),
            .I(N__19071));
    CascadeMux I__3278 (
            .O(N__19130),
            .I(N__19068));
    CascadeMux I__3277 (
            .O(N__19129),
            .I(N__19050));
    CascadeMux I__3276 (
            .O(N__19128),
            .I(N__19047));
    CascadeMux I__3275 (
            .O(N__19127),
            .I(N__19042));
    InMux I__3274 (
            .O(N__19126),
            .I(N__19036));
    InMux I__3273 (
            .O(N__19125),
            .I(N__19027));
    InMux I__3272 (
            .O(N__19124),
            .I(N__19027));
    InMux I__3271 (
            .O(N__19121),
            .I(N__19027));
    InMux I__3270 (
            .O(N__19120),
            .I(N__19027));
    InMux I__3269 (
            .O(N__19119),
            .I(N__19020));
    InMux I__3268 (
            .O(N__19118),
            .I(N__19020));
    InMux I__3267 (
            .O(N__19117),
            .I(N__19020));
    LocalMux I__3266 (
            .O(N__19114),
            .I(N__19017));
    InMux I__3265 (
            .O(N__19113),
            .I(N__19012));
    InMux I__3264 (
            .O(N__19112),
            .I(N__19012));
    LocalMux I__3263 (
            .O(N__19109),
            .I(N__19009));
    InMux I__3262 (
            .O(N__19108),
            .I(N__19006));
    LocalMux I__3261 (
            .O(N__19105),
            .I(N__19003));
    LocalMux I__3260 (
            .O(N__19102),
            .I(N__18992));
    LocalMux I__3259 (
            .O(N__19099),
            .I(N__18992));
    Span4Mux_v I__3258 (
            .O(N__19096),
            .I(N__18992));
    Span4Mux_s1_h I__3257 (
            .O(N__19093),
            .I(N__18992));
    LocalMux I__3256 (
            .O(N__19090),
            .I(N__18992));
    InMux I__3255 (
            .O(N__19089),
            .I(N__18987));
    InMux I__3254 (
            .O(N__19088),
            .I(N__18987));
    InMux I__3253 (
            .O(N__19087),
            .I(N__18982));
    InMux I__3252 (
            .O(N__19086),
            .I(N__18982));
    InMux I__3251 (
            .O(N__19085),
            .I(N__18971));
    InMux I__3250 (
            .O(N__19084),
            .I(N__18971));
    InMux I__3249 (
            .O(N__19081),
            .I(N__18971));
    InMux I__3248 (
            .O(N__19078),
            .I(N__18971));
    InMux I__3247 (
            .O(N__19075),
            .I(N__18971));
    InMux I__3246 (
            .O(N__19074),
            .I(N__18964));
    InMux I__3245 (
            .O(N__19071),
            .I(N__18964));
    InMux I__3244 (
            .O(N__19068),
            .I(N__18964));
    InMux I__3243 (
            .O(N__19067),
            .I(N__18959));
    InMux I__3242 (
            .O(N__19066),
            .I(N__18959));
    InMux I__3241 (
            .O(N__19065),
            .I(N__18956));
    InMux I__3240 (
            .O(N__19064),
            .I(N__18949));
    InMux I__3239 (
            .O(N__19063),
            .I(N__18949));
    InMux I__3238 (
            .O(N__19062),
            .I(N__18949));
    InMux I__3237 (
            .O(N__19061),
            .I(N__18934));
    InMux I__3236 (
            .O(N__19060),
            .I(N__18934));
    InMux I__3235 (
            .O(N__19059),
            .I(N__18934));
    InMux I__3234 (
            .O(N__19058),
            .I(N__18934));
    InMux I__3233 (
            .O(N__19057),
            .I(N__18934));
    InMux I__3232 (
            .O(N__19056),
            .I(N__18934));
    InMux I__3231 (
            .O(N__19055),
            .I(N__18934));
    InMux I__3230 (
            .O(N__19054),
            .I(N__18923));
    InMux I__3229 (
            .O(N__19053),
            .I(N__18923));
    InMux I__3228 (
            .O(N__19050),
            .I(N__18923));
    InMux I__3227 (
            .O(N__19047),
            .I(N__18923));
    InMux I__3226 (
            .O(N__19046),
            .I(N__18923));
    InMux I__3225 (
            .O(N__19045),
            .I(N__18912));
    InMux I__3224 (
            .O(N__19042),
            .I(N__18912));
    InMux I__3223 (
            .O(N__19041),
            .I(N__18912));
    InMux I__3222 (
            .O(N__19040),
            .I(N__18912));
    InMux I__3221 (
            .O(N__19039),
            .I(N__18912));
    LocalMux I__3220 (
            .O(N__19036),
            .I(N__18907));
    LocalMux I__3219 (
            .O(N__19027),
            .I(N__18907));
    LocalMux I__3218 (
            .O(N__19020),
            .I(N__18904));
    Span12Mux_s3_h I__3217 (
            .O(N__19017),
            .I(N__18901));
    LocalMux I__3216 (
            .O(N__19012),
            .I(N__18896));
    Span4Mux_v I__3215 (
            .O(N__19009),
            .I(N__18896));
    LocalMux I__3214 (
            .O(N__19006),
            .I(N__18889));
    Span4Mux_v I__3213 (
            .O(N__19003),
            .I(N__18889));
    Span4Mux_v I__3212 (
            .O(N__18992),
            .I(N__18889));
    LocalMux I__3211 (
            .O(N__18987),
            .I(n9069));
    LocalMux I__3210 (
            .O(N__18982),
            .I(n9069));
    LocalMux I__3209 (
            .O(N__18971),
            .I(n9069));
    LocalMux I__3208 (
            .O(N__18964),
            .I(n9069));
    LocalMux I__3207 (
            .O(N__18959),
            .I(n9069));
    LocalMux I__3206 (
            .O(N__18956),
            .I(n9069));
    LocalMux I__3205 (
            .O(N__18949),
            .I(n9069));
    LocalMux I__3204 (
            .O(N__18934),
            .I(n9069));
    LocalMux I__3203 (
            .O(N__18923),
            .I(n9069));
    LocalMux I__3202 (
            .O(N__18912),
            .I(n9069));
    Odrv4 I__3201 (
            .O(N__18907),
            .I(n9069));
    Odrv4 I__3200 (
            .O(N__18904),
            .I(n9069));
    Odrv12 I__3199 (
            .O(N__18901),
            .I(n9069));
    Odrv4 I__3198 (
            .O(N__18896),
            .I(n9069));
    Odrv4 I__3197 (
            .O(N__18889),
            .I(n9069));
    InMux I__3196 (
            .O(N__18858),
            .I(N__18854));
    CascadeMux I__3195 (
            .O(N__18857),
            .I(N__18851));
    LocalMux I__3194 (
            .O(N__18854),
            .I(N__18846));
    InMux I__3193 (
            .O(N__18851),
            .I(N__18843));
    InMux I__3192 (
            .O(N__18850),
            .I(N__18840));
    InMux I__3191 (
            .O(N__18849),
            .I(N__18837));
    Span4Mux_h I__3190 (
            .O(N__18846),
            .I(N__18834));
    LocalMux I__3189 (
            .O(N__18843),
            .I(N__18831));
    LocalMux I__3188 (
            .O(N__18840),
            .I(data_in_field_45));
    LocalMux I__3187 (
            .O(N__18837),
            .I(data_in_field_45));
    Odrv4 I__3186 (
            .O(N__18834),
            .I(data_in_field_45));
    Odrv12 I__3185 (
            .O(N__18831),
            .I(data_in_field_45));
    CascadeMux I__3184 (
            .O(N__18822),
            .I(N__18819));
    InMux I__3183 (
            .O(N__18819),
            .I(N__18816));
    LocalMux I__3182 (
            .O(N__18816),
            .I(\c0.n9602 ));
    InMux I__3181 (
            .O(N__18813),
            .I(N__18809));
    CascadeMux I__3180 (
            .O(N__18812),
            .I(N__18806));
    LocalMux I__3179 (
            .O(N__18809),
            .I(N__18803));
    InMux I__3178 (
            .O(N__18806),
            .I(N__18798));
    Span4Mux_h I__3177 (
            .O(N__18803),
            .I(N__18795));
    InMux I__3176 (
            .O(N__18802),
            .I(N__18792));
    InMux I__3175 (
            .O(N__18801),
            .I(N__18789));
    LocalMux I__3174 (
            .O(N__18798),
            .I(\c0.data_in_field_12 ));
    Odrv4 I__3173 (
            .O(N__18795),
            .I(\c0.data_in_field_12 ));
    LocalMux I__3172 (
            .O(N__18792),
            .I(\c0.data_in_field_12 ));
    LocalMux I__3171 (
            .O(N__18789),
            .I(\c0.data_in_field_12 ));
    InMux I__3170 (
            .O(N__18780),
            .I(N__18777));
    LocalMux I__3169 (
            .O(N__18777),
            .I(N__18774));
    Span4Mux_v I__3168 (
            .O(N__18774),
            .I(N__18770));
    InMux I__3167 (
            .O(N__18773),
            .I(N__18767));
    Sp12to4 I__3166 (
            .O(N__18770),
            .I(N__18762));
    LocalMux I__3165 (
            .O(N__18767),
            .I(N__18762));
    Odrv12 I__3164 (
            .O(N__18762),
            .I(\c0.n9019 ));
    InMux I__3163 (
            .O(N__18759),
            .I(N__18754));
    InMux I__3162 (
            .O(N__18758),
            .I(N__18751));
    InMux I__3161 (
            .O(N__18757),
            .I(N__18748));
    LocalMux I__3160 (
            .O(N__18754),
            .I(N__18745));
    LocalMux I__3159 (
            .O(N__18751),
            .I(N__18740));
    LocalMux I__3158 (
            .O(N__18748),
            .I(N__18737));
    Span4Mux_h I__3157 (
            .O(N__18745),
            .I(N__18734));
    InMux I__3156 (
            .O(N__18744),
            .I(N__18729));
    InMux I__3155 (
            .O(N__18743),
            .I(N__18729));
    Odrv4 I__3154 (
            .O(N__18740),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__3153 (
            .O(N__18737),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__3152 (
            .O(N__18734),
            .I(\c0.data_in_field_28 ));
    LocalMux I__3151 (
            .O(N__18729),
            .I(\c0.data_in_field_28 ));
    CascadeMux I__3150 (
            .O(N__18720),
            .I(\c0.n9746_cascade_ ));
    InMux I__3149 (
            .O(N__18717),
            .I(N__18712));
    InMux I__3148 (
            .O(N__18716),
            .I(N__18708));
    InMux I__3147 (
            .O(N__18715),
            .I(N__18704));
    LocalMux I__3146 (
            .O(N__18712),
            .I(N__18701));
    InMux I__3145 (
            .O(N__18711),
            .I(N__18698));
    LocalMux I__3144 (
            .O(N__18708),
            .I(N__18695));
    InMux I__3143 (
            .O(N__18707),
            .I(N__18692));
    LocalMux I__3142 (
            .O(N__18704),
            .I(\c0.data_in_field_32 ));
    Odrv4 I__3141 (
            .O(N__18701),
            .I(\c0.data_in_field_32 ));
    LocalMux I__3140 (
            .O(N__18698),
            .I(\c0.data_in_field_32 ));
    Odrv4 I__3139 (
            .O(N__18695),
            .I(\c0.data_in_field_32 ));
    LocalMux I__3138 (
            .O(N__18692),
            .I(\c0.data_in_field_32 ));
    InMux I__3137 (
            .O(N__18681),
            .I(N__18678));
    LocalMux I__3136 (
            .O(N__18678),
            .I(N__18672));
    InMux I__3135 (
            .O(N__18677),
            .I(N__18669));
    InMux I__3134 (
            .O(N__18676),
            .I(N__18665));
    InMux I__3133 (
            .O(N__18675),
            .I(N__18662));
    Span4Mux_h I__3132 (
            .O(N__18672),
            .I(N__18659));
    LocalMux I__3131 (
            .O(N__18669),
            .I(N__18656));
    InMux I__3130 (
            .O(N__18668),
            .I(N__18653));
    LocalMux I__3129 (
            .O(N__18665),
            .I(data_in_field_42));
    LocalMux I__3128 (
            .O(N__18662),
            .I(data_in_field_42));
    Odrv4 I__3127 (
            .O(N__18659),
            .I(data_in_field_42));
    Odrv4 I__3126 (
            .O(N__18656),
            .I(data_in_field_42));
    LocalMux I__3125 (
            .O(N__18653),
            .I(data_in_field_42));
    InMux I__3124 (
            .O(N__18642),
            .I(N__18637));
    InMux I__3123 (
            .O(N__18641),
            .I(N__18631));
    InMux I__3122 (
            .O(N__18640),
            .I(N__18628));
    LocalMux I__3121 (
            .O(N__18637),
            .I(N__18625));
    InMux I__3120 (
            .O(N__18636),
            .I(N__18622));
    InMux I__3119 (
            .O(N__18635),
            .I(N__18617));
    InMux I__3118 (
            .O(N__18634),
            .I(N__18617));
    LocalMux I__3117 (
            .O(N__18631),
            .I(data_in_field_40));
    LocalMux I__3116 (
            .O(N__18628),
            .I(data_in_field_40));
    Odrv4 I__3115 (
            .O(N__18625),
            .I(data_in_field_40));
    LocalMux I__3114 (
            .O(N__18622),
            .I(data_in_field_40));
    LocalMux I__3113 (
            .O(N__18617),
            .I(data_in_field_40));
    InMux I__3112 (
            .O(N__18606),
            .I(N__18603));
    LocalMux I__3111 (
            .O(N__18603),
            .I(N__18598));
    InMux I__3110 (
            .O(N__18602),
            .I(N__18593));
    InMux I__3109 (
            .O(N__18601),
            .I(N__18593));
    Span4Mux_h I__3108 (
            .O(N__18598),
            .I(N__18590));
    LocalMux I__3107 (
            .O(N__18593),
            .I(N__18587));
    Odrv4 I__3106 (
            .O(N__18590),
            .I(\c0.n4208 ));
    Odrv12 I__3105 (
            .O(N__18587),
            .I(\c0.n4208 ));
    InMux I__3104 (
            .O(N__18582),
            .I(N__18579));
    LocalMux I__3103 (
            .O(N__18579),
            .I(N__18574));
    InMux I__3102 (
            .O(N__18578),
            .I(N__18570));
    InMux I__3101 (
            .O(N__18577),
            .I(N__18567));
    Span4Mux_v I__3100 (
            .O(N__18574),
            .I(N__18564));
    InMux I__3099 (
            .O(N__18573),
            .I(N__18561));
    LocalMux I__3098 (
            .O(N__18570),
            .I(data_in_3_4));
    LocalMux I__3097 (
            .O(N__18567),
            .I(data_in_3_4));
    Odrv4 I__3096 (
            .O(N__18564),
            .I(data_in_3_4));
    LocalMux I__3095 (
            .O(N__18561),
            .I(data_in_3_4));
    InMux I__3094 (
            .O(N__18552),
            .I(N__18548));
    InMux I__3093 (
            .O(N__18551),
            .I(N__18545));
    LocalMux I__3092 (
            .O(N__18548),
            .I(N__18540));
    LocalMux I__3091 (
            .O(N__18545),
            .I(N__18537));
    InMux I__3090 (
            .O(N__18544),
            .I(N__18534));
    InMux I__3089 (
            .O(N__18543),
            .I(N__18531));
    Span4Mux_h I__3088 (
            .O(N__18540),
            .I(N__18528));
    Odrv4 I__3087 (
            .O(N__18537),
            .I(data_in_3_2));
    LocalMux I__3086 (
            .O(N__18534),
            .I(data_in_3_2));
    LocalMux I__3085 (
            .O(N__18531),
            .I(data_in_3_2));
    Odrv4 I__3084 (
            .O(N__18528),
            .I(data_in_3_2));
    CascadeMux I__3083 (
            .O(N__18519),
            .I(N__18516));
    InMux I__3082 (
            .O(N__18516),
            .I(N__18512));
    InMux I__3081 (
            .O(N__18515),
            .I(N__18509));
    LocalMux I__3080 (
            .O(N__18512),
            .I(N__18504));
    LocalMux I__3079 (
            .O(N__18509),
            .I(N__18501));
    InMux I__3078 (
            .O(N__18508),
            .I(N__18496));
    InMux I__3077 (
            .O(N__18507),
            .I(N__18496));
    Span4Mux_h I__3076 (
            .O(N__18504),
            .I(N__18493));
    Span4Mux_h I__3075 (
            .O(N__18501),
            .I(N__18490));
    LocalMux I__3074 (
            .O(N__18496),
            .I(data_in_2_4));
    Odrv4 I__3073 (
            .O(N__18493),
            .I(data_in_2_4));
    Odrv4 I__3072 (
            .O(N__18490),
            .I(data_in_2_4));
    InMux I__3071 (
            .O(N__18483),
            .I(N__18479));
    InMux I__3070 (
            .O(N__18482),
            .I(N__18476));
    LocalMux I__3069 (
            .O(N__18479),
            .I(data_in_17_0));
    LocalMux I__3068 (
            .O(N__18476),
            .I(data_in_17_0));
    InMux I__3067 (
            .O(N__18471),
            .I(N__18467));
    InMux I__3066 (
            .O(N__18470),
            .I(N__18464));
    LocalMux I__3065 (
            .O(N__18467),
            .I(N__18459));
    LocalMux I__3064 (
            .O(N__18464),
            .I(N__18459));
    Span4Mux_h I__3063 (
            .O(N__18459),
            .I(N__18456));
    Span4Mux_v I__3062 (
            .O(N__18456),
            .I(N__18453));
    Odrv4 I__3061 (
            .O(N__18453),
            .I(\c0.n8960 ));
    InMux I__3060 (
            .O(N__18450),
            .I(N__18446));
    InMux I__3059 (
            .O(N__18449),
            .I(N__18443));
    LocalMux I__3058 (
            .O(N__18446),
            .I(N__18440));
    LocalMux I__3057 (
            .O(N__18443),
            .I(N__18436));
    Span4Mux_h I__3056 (
            .O(N__18440),
            .I(N__18433));
    InMux I__3055 (
            .O(N__18439),
            .I(N__18430));
    Span4Mux_h I__3054 (
            .O(N__18436),
            .I(N__18427));
    Odrv4 I__3053 (
            .O(N__18433),
            .I(data_in_0_4));
    LocalMux I__3052 (
            .O(N__18430),
            .I(data_in_0_4));
    Odrv4 I__3051 (
            .O(N__18427),
            .I(data_in_0_4));
    InMux I__3050 (
            .O(N__18420),
            .I(N__18417));
    LocalMux I__3049 (
            .O(N__18417),
            .I(N__18414));
    Odrv4 I__3048 (
            .O(N__18414),
            .I(n1890));
    InMux I__3047 (
            .O(N__18411),
            .I(N__18408));
    LocalMux I__3046 (
            .O(N__18408),
            .I(N__18405));
    Span4Mux_v I__3045 (
            .O(N__18405),
            .I(N__18401));
    InMux I__3044 (
            .O(N__18404),
            .I(N__18398));
    Odrv4 I__3043 (
            .O(N__18401),
            .I(data_in_14_0));
    LocalMux I__3042 (
            .O(N__18398),
            .I(data_in_14_0));
    InMux I__3041 (
            .O(N__18393),
            .I(N__18387));
    InMux I__3040 (
            .O(N__18392),
            .I(N__18387));
    LocalMux I__3039 (
            .O(N__18387),
            .I(data_in_15_0));
    InMux I__3038 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__3037 (
            .O(N__18381),
            .I(N__18376));
    InMux I__3036 (
            .O(N__18380),
            .I(N__18370));
    InMux I__3035 (
            .O(N__18379),
            .I(N__18370));
    Span4Mux_h I__3034 (
            .O(N__18376),
            .I(N__18367));
    InMux I__3033 (
            .O(N__18375),
            .I(N__18364));
    LocalMux I__3032 (
            .O(N__18370),
            .I(N__18361));
    Odrv4 I__3031 (
            .O(N__18367),
            .I(data_in_2_2));
    LocalMux I__3030 (
            .O(N__18364),
            .I(data_in_2_2));
    Odrv12 I__3029 (
            .O(N__18361),
            .I(data_in_2_2));
    InMux I__3028 (
            .O(N__18354),
            .I(N__18348));
    InMux I__3027 (
            .O(N__18353),
            .I(N__18348));
    LocalMux I__3026 (
            .O(N__18348),
            .I(data_in_16_0));
    CascadeMux I__3025 (
            .O(N__18345),
            .I(N__18342));
    InMux I__3024 (
            .O(N__18342),
            .I(N__18336));
    InMux I__3023 (
            .O(N__18341),
            .I(N__18336));
    LocalMux I__3022 (
            .O(N__18336),
            .I(data_in_20_0));
    InMux I__3021 (
            .O(N__18333),
            .I(N__18330));
    LocalMux I__3020 (
            .O(N__18330),
            .I(N__18327));
    Odrv4 I__3019 (
            .O(N__18327),
            .I(n1898));
    InMux I__3018 (
            .O(N__18324),
            .I(N__18320));
    InMux I__3017 (
            .O(N__18323),
            .I(N__18317));
    LocalMux I__3016 (
            .O(N__18320),
            .I(data_in_20_5));
    LocalMux I__3015 (
            .O(N__18317),
            .I(data_in_20_5));
    InMux I__3014 (
            .O(N__18312),
            .I(N__18303));
    InMux I__3013 (
            .O(N__18311),
            .I(N__18303));
    InMux I__3012 (
            .O(N__18310),
            .I(N__18303));
    LocalMux I__3011 (
            .O(N__18303),
            .I(data_in_5_5));
    CascadeMux I__3010 (
            .O(N__18300),
            .I(N__18297));
    InMux I__3009 (
            .O(N__18297),
            .I(N__18294));
    LocalMux I__3008 (
            .O(N__18294),
            .I(N__18291));
    Span4Mux_h I__3007 (
            .O(N__18291),
            .I(N__18286));
    InMux I__3006 (
            .O(N__18290),
            .I(N__18283));
    InMux I__3005 (
            .O(N__18289),
            .I(N__18280));
    Span4Mux_h I__3004 (
            .O(N__18286),
            .I(N__18277));
    LocalMux I__3003 (
            .O(N__18283),
            .I(data_in_4_5));
    LocalMux I__3002 (
            .O(N__18280),
            .I(data_in_4_5));
    Odrv4 I__3001 (
            .O(N__18277),
            .I(data_in_4_5));
    InMux I__3000 (
            .O(N__18270),
            .I(N__18261));
    InMux I__2999 (
            .O(N__18269),
            .I(N__18261));
    InMux I__2998 (
            .O(N__18268),
            .I(N__18261));
    LocalMux I__2997 (
            .O(N__18261),
            .I(data_in_6_5));
    InMux I__2996 (
            .O(N__18258),
            .I(N__18252));
    InMux I__2995 (
            .O(N__18257),
            .I(N__18252));
    LocalMux I__2994 (
            .O(N__18252),
            .I(data_in_7_5));
    InMux I__2993 (
            .O(N__18249),
            .I(N__18243));
    InMux I__2992 (
            .O(N__18248),
            .I(N__18243));
    LocalMux I__2991 (
            .O(N__18243),
            .I(data_in_8_5));
    InMux I__2990 (
            .O(N__18240),
            .I(N__18234));
    InMux I__2989 (
            .O(N__18239),
            .I(N__18234));
    LocalMux I__2988 (
            .O(N__18234),
            .I(data_in_9_5));
    InMux I__2987 (
            .O(N__18231),
            .I(N__18227));
    InMux I__2986 (
            .O(N__18230),
            .I(N__18224));
    LocalMux I__2985 (
            .O(N__18227),
            .I(data_in_16_3));
    LocalMux I__2984 (
            .O(N__18224),
            .I(data_in_16_3));
    InMux I__2983 (
            .O(N__18219),
            .I(N__18213));
    InMux I__2982 (
            .O(N__18218),
            .I(N__18213));
    LocalMux I__2981 (
            .O(N__18213),
            .I(data_in_15_3));
    InMux I__2980 (
            .O(N__18210),
            .I(N__18206));
    InMux I__2979 (
            .O(N__18209),
            .I(N__18203));
    LocalMux I__2978 (
            .O(N__18206),
            .I(data_in_17_3));
    LocalMux I__2977 (
            .O(N__18203),
            .I(data_in_17_3));
    InMux I__2976 (
            .O(N__18198),
            .I(N__18194));
    InMux I__2975 (
            .O(N__18197),
            .I(N__18191));
    LocalMux I__2974 (
            .O(N__18194),
            .I(data_in_18_3));
    LocalMux I__2973 (
            .O(N__18191),
            .I(data_in_18_3));
    InMux I__2972 (
            .O(N__18186),
            .I(N__18180));
    InMux I__2971 (
            .O(N__18185),
            .I(N__18180));
    LocalMux I__2970 (
            .O(N__18180),
            .I(data_in_19_3));
    InMux I__2969 (
            .O(N__18177),
            .I(N__18171));
    InMux I__2968 (
            .O(N__18176),
            .I(N__18171));
    LocalMux I__2967 (
            .O(N__18171),
            .I(data_in_20_3));
    InMux I__2966 (
            .O(N__18168),
            .I(N__18162));
    InMux I__2965 (
            .O(N__18167),
            .I(N__18162));
    LocalMux I__2964 (
            .O(N__18162),
            .I(data_in_19_5));
    InMux I__2963 (
            .O(N__18159),
            .I(N__18156));
    LocalMux I__2962 (
            .O(N__18156),
            .I(N__18152));
    InMux I__2961 (
            .O(N__18155),
            .I(N__18149));
    Odrv4 I__2960 (
            .O(N__18152),
            .I(data_in_17_6));
    LocalMux I__2959 (
            .O(N__18149),
            .I(data_in_17_6));
    InMux I__2958 (
            .O(N__18144),
            .I(N__18141));
    LocalMux I__2957 (
            .O(N__18141),
            .I(N__18137));
    InMux I__2956 (
            .O(N__18140),
            .I(N__18134));
    Odrv4 I__2955 (
            .O(N__18137),
            .I(data_in_10_3));
    LocalMux I__2954 (
            .O(N__18134),
            .I(data_in_10_3));
    InMux I__2953 (
            .O(N__18129),
            .I(N__18126));
    LocalMux I__2952 (
            .O(N__18126),
            .I(N__18122));
    InMux I__2951 (
            .O(N__18125),
            .I(N__18119));
    Odrv4 I__2950 (
            .O(N__18122),
            .I(data_in_9_3));
    LocalMux I__2949 (
            .O(N__18119),
            .I(data_in_9_3));
    CascadeMux I__2948 (
            .O(N__18114),
            .I(\c0.n3056_cascade_ ));
    InMux I__2947 (
            .O(N__18111),
            .I(N__18108));
    LocalMux I__2946 (
            .O(N__18108),
            .I(N__18105));
    Span4Mux_h I__2945 (
            .O(N__18105),
            .I(N__18102));
    Odrv4 I__2944 (
            .O(N__18102),
            .I(\c0.n22_adj_1676 ));
    InMux I__2943 (
            .O(N__18099),
            .I(N__18096));
    LocalMux I__2942 (
            .O(N__18096),
            .I(\c0.n38_adj_1616 ));
    CascadeMux I__2941 (
            .O(N__18093),
            .I(N__18090));
    InMux I__2940 (
            .O(N__18090),
            .I(N__18087));
    LocalMux I__2939 (
            .O(N__18087),
            .I(N__18084));
    Odrv4 I__2938 (
            .O(N__18084),
            .I(\c0.n36 ));
    InMux I__2937 (
            .O(N__18081),
            .I(N__18078));
    LocalMux I__2936 (
            .O(N__18078),
            .I(\c0.n37 ));
    CascadeMux I__2935 (
            .O(N__18075),
            .I(N__18072));
    InMux I__2934 (
            .O(N__18072),
            .I(N__18069));
    LocalMux I__2933 (
            .O(N__18069),
            .I(\c0.data_in_frame_19_7 ));
    InMux I__2932 (
            .O(N__18066),
            .I(N__18063));
    LocalMux I__2931 (
            .O(N__18063),
            .I(N__18058));
    InMux I__2930 (
            .O(N__18062),
            .I(N__18052));
    InMux I__2929 (
            .O(N__18061),
            .I(N__18052));
    Span4Mux_s2_v I__2928 (
            .O(N__18058),
            .I(N__18049));
    InMux I__2927 (
            .O(N__18057),
            .I(N__18046));
    LocalMux I__2926 (
            .O(N__18052),
            .I(data_in_field_135));
    Odrv4 I__2925 (
            .O(N__18049),
            .I(data_in_field_135));
    LocalMux I__2924 (
            .O(N__18046),
            .I(data_in_field_135));
    CascadeMux I__2923 (
            .O(N__18039),
            .I(\c0.n9662_cascade_ ));
    InMux I__2922 (
            .O(N__18036),
            .I(N__18033));
    LocalMux I__2921 (
            .O(N__18033),
            .I(\c0.n9665 ));
    InMux I__2920 (
            .O(N__18030),
            .I(N__18024));
    InMux I__2919 (
            .O(N__18029),
            .I(N__18024));
    LocalMux I__2918 (
            .O(N__18024),
            .I(data_in_13_3));
    InMux I__2917 (
            .O(N__18021),
            .I(N__18015));
    InMux I__2916 (
            .O(N__18020),
            .I(N__18015));
    LocalMux I__2915 (
            .O(N__18015),
            .I(data_in_14_3));
    CascadeMux I__2914 (
            .O(N__18012),
            .I(\c0.n6_adj_1604_cascade_ ));
    InMux I__2913 (
            .O(N__18009),
            .I(N__18006));
    LocalMux I__2912 (
            .O(N__18006),
            .I(N__18003));
    Span4Mux_h I__2911 (
            .O(N__18003),
            .I(N__18000));
    Odrv4 I__2910 (
            .O(N__18000),
            .I(\c0.n8983 ));
    InMux I__2909 (
            .O(N__17997),
            .I(N__17994));
    LocalMux I__2908 (
            .O(N__17994),
            .I(N__17991));
    Span12Mux_s5_v I__2907 (
            .O(N__17991),
            .I(N__17988));
    Odrv12 I__2906 (
            .O(N__17988),
            .I(\c0.n8948 ));
    InMux I__2905 (
            .O(N__17985),
            .I(N__17982));
    LocalMux I__2904 (
            .O(N__17982),
            .I(N__17979));
    Odrv4 I__2903 (
            .O(N__17979),
            .I(\c0.n8945 ));
    CascadeMux I__2902 (
            .O(N__17976),
            .I(\c0.n8983_cascade_ ));
    InMux I__2901 (
            .O(N__17973),
            .I(N__17970));
    LocalMux I__2900 (
            .O(N__17970),
            .I(N__17967));
    Span12Mux_s3_v I__2899 (
            .O(N__17967),
            .I(N__17963));
    InMux I__2898 (
            .O(N__17966),
            .I(N__17960));
    Odrv12 I__2897 (
            .O(N__17963),
            .I(\c0.n9004 ));
    LocalMux I__2896 (
            .O(N__17960),
            .I(\c0.n9004 ));
    CascadeMux I__2895 (
            .O(N__17955),
            .I(N__17951));
    InMux I__2894 (
            .O(N__17954),
            .I(N__17948));
    InMux I__2893 (
            .O(N__17951),
            .I(N__17945));
    LocalMux I__2892 (
            .O(N__17948),
            .I(N__17939));
    LocalMux I__2891 (
            .O(N__17945),
            .I(N__17936));
    InMux I__2890 (
            .O(N__17944),
            .I(N__17933));
    InMux I__2889 (
            .O(N__17943),
            .I(N__17928));
    InMux I__2888 (
            .O(N__17942),
            .I(N__17928));
    Span12Mux_h I__2887 (
            .O(N__17939),
            .I(N__17925));
    Span4Mux_s2_h I__2886 (
            .O(N__17936),
            .I(N__17922));
    LocalMux I__2885 (
            .O(N__17933),
            .I(data_in_field_89));
    LocalMux I__2884 (
            .O(N__17928),
            .I(data_in_field_89));
    Odrv12 I__2883 (
            .O(N__17925),
            .I(data_in_field_89));
    Odrv4 I__2882 (
            .O(N__17922),
            .I(data_in_field_89));
    InMux I__2881 (
            .O(N__17913),
            .I(N__17909));
    InMux I__2880 (
            .O(N__17912),
            .I(N__17906));
    LocalMux I__2879 (
            .O(N__17909),
            .I(N__17903));
    LocalMux I__2878 (
            .O(N__17906),
            .I(\c0.n4203 ));
    Odrv4 I__2877 (
            .O(N__17903),
            .I(\c0.n4203 ));
    InMux I__2876 (
            .O(N__17898),
            .I(N__17895));
    LocalMux I__2875 (
            .O(N__17895),
            .I(N__17892));
    Span4Mux_s2_v I__2874 (
            .O(N__17892),
            .I(N__17889));
    Odrv4 I__2873 (
            .O(N__17889),
            .I(\c0.n8890 ));
    InMux I__2872 (
            .O(N__17886),
            .I(N__17882));
    InMux I__2871 (
            .O(N__17885),
            .I(N__17879));
    LocalMux I__2870 (
            .O(N__17882),
            .I(\c0.n8874 ));
    LocalMux I__2869 (
            .O(N__17879),
            .I(\c0.n8874 ));
    InMux I__2868 (
            .O(N__17874),
            .I(N__17871));
    LocalMux I__2867 (
            .O(N__17871),
            .I(N__17868));
    Span4Mux_s2_v I__2866 (
            .O(N__17868),
            .I(N__17865));
    Odrv4 I__2865 (
            .O(N__17865),
            .I(\c0.n24_adj_1607 ));
    InMux I__2864 (
            .O(N__17862),
            .I(N__17859));
    LocalMux I__2863 (
            .O(N__17859),
            .I(\c0.n23 ));
    CascadeMux I__2862 (
            .O(N__17856),
            .I(\c0.n25_cascade_ ));
    InMux I__2861 (
            .O(N__17853),
            .I(N__17850));
    LocalMux I__2860 (
            .O(N__17850),
            .I(\c0.n26_adj_1606 ));
    InMux I__2859 (
            .O(N__17847),
            .I(N__17844));
    LocalMux I__2858 (
            .O(N__17844),
            .I(N__17841));
    Span4Mux_v I__2857 (
            .O(N__17841),
            .I(N__17838));
    Span4Mux_h I__2856 (
            .O(N__17838),
            .I(N__17835));
    Odrv4 I__2855 (
            .O(N__17835),
            .I(\c0.data_in_frame_20_3 ));
    InMux I__2854 (
            .O(N__17832),
            .I(N__17829));
    LocalMux I__2853 (
            .O(N__17829),
            .I(N__17825));
    InMux I__2852 (
            .O(N__17828),
            .I(N__17822));
    Span4Mux_v I__2851 (
            .O(N__17825),
            .I(N__17819));
    LocalMux I__2850 (
            .O(N__17822),
            .I(N__17816));
    Span4Mux_h I__2849 (
            .O(N__17819),
            .I(N__17811));
    Span4Mux_s1_v I__2848 (
            .O(N__17816),
            .I(N__17811));
    Span4Mux_v I__2847 (
            .O(N__17811),
            .I(N__17808));
    Odrv4 I__2846 (
            .O(N__17808),
            .I(\c0.n8974 ));
    CascadeMux I__2845 (
            .O(N__17805),
            .I(N__17802));
    InMux I__2844 (
            .O(N__17802),
            .I(N__17799));
    LocalMux I__2843 (
            .O(N__17799),
            .I(N__17796));
    Span4Mux_s2_v I__2842 (
            .O(N__17796),
            .I(N__17793));
    Odrv4 I__2841 (
            .O(N__17793),
            .I(\c0.n22_adj_1617 ));
    InMux I__2840 (
            .O(N__17790),
            .I(N__17787));
    LocalMux I__2839 (
            .O(N__17787),
            .I(N__17784));
    Span4Mux_s3_v I__2838 (
            .O(N__17784),
            .I(N__17781));
    Odrv4 I__2837 (
            .O(N__17781),
            .I(\c0.n8933 ));
    InMux I__2836 (
            .O(N__17778),
            .I(N__17775));
    LocalMux I__2835 (
            .O(N__17775),
            .I(N__17772));
    Span4Mux_s2_v I__2834 (
            .O(N__17772),
            .I(N__17769));
    Span4Mux_v I__2833 (
            .O(N__17769),
            .I(N__17766));
    Odrv4 I__2832 (
            .O(N__17766),
            .I(\c0.data_in_frame_20_7 ));
    InMux I__2831 (
            .O(N__17763),
            .I(N__17757));
    InMux I__2830 (
            .O(N__17762),
            .I(N__17757));
    LocalMux I__2829 (
            .O(N__17757),
            .I(N__17752));
    InMux I__2828 (
            .O(N__17756),
            .I(N__17749));
    InMux I__2827 (
            .O(N__17755),
            .I(N__17746));
    Span4Mux_v I__2826 (
            .O(N__17752),
            .I(N__17741));
    LocalMux I__2825 (
            .O(N__17749),
            .I(N__17741));
    LocalMux I__2824 (
            .O(N__17746),
            .I(data_in_field_111));
    Odrv4 I__2823 (
            .O(N__17741),
            .I(data_in_field_111));
    CascadeMux I__2822 (
            .O(N__17736),
            .I(\c0.n4525_cascade_ ));
    InMux I__2821 (
            .O(N__17733),
            .I(N__17729));
    InMux I__2820 (
            .O(N__17732),
            .I(N__17725));
    LocalMux I__2819 (
            .O(N__17729),
            .I(N__17722));
    InMux I__2818 (
            .O(N__17728),
            .I(N__17719));
    LocalMux I__2817 (
            .O(N__17725),
            .I(N__17714));
    Span4Mux_h I__2816 (
            .O(N__17722),
            .I(N__17714));
    LocalMux I__2815 (
            .O(N__17719),
            .I(data_in_field_107));
    Odrv4 I__2814 (
            .O(N__17714),
            .I(data_in_field_107));
    InMux I__2813 (
            .O(N__17709),
            .I(N__17706));
    LocalMux I__2812 (
            .O(N__17706),
            .I(N__17700));
    InMux I__2811 (
            .O(N__17705),
            .I(N__17697));
    InMux I__2810 (
            .O(N__17704),
            .I(N__17692));
    InMux I__2809 (
            .O(N__17703),
            .I(N__17692));
    Span4Mux_h I__2808 (
            .O(N__17700),
            .I(N__17687));
    LocalMux I__2807 (
            .O(N__17697),
            .I(N__17687));
    LocalMux I__2806 (
            .O(N__17692),
            .I(data_in_field_137));
    Odrv4 I__2805 (
            .O(N__17687),
            .I(data_in_field_137));
    CascadeMux I__2804 (
            .O(N__17682),
            .I(\c0.n8874_cascade_ ));
    InMux I__2803 (
            .O(N__17679),
            .I(N__17675));
    InMux I__2802 (
            .O(N__17678),
            .I(N__17672));
    LocalMux I__2801 (
            .O(N__17675),
            .I(N__17668));
    LocalMux I__2800 (
            .O(N__17672),
            .I(N__17665));
    InMux I__2799 (
            .O(N__17671),
            .I(N__17661));
    Span4Mux_v I__2798 (
            .O(N__17668),
            .I(N__17658));
    Span4Mux_v I__2797 (
            .O(N__17665),
            .I(N__17655));
    InMux I__2796 (
            .O(N__17664),
            .I(N__17652));
    LocalMux I__2795 (
            .O(N__17661),
            .I(data_in_field_55));
    Odrv4 I__2794 (
            .O(N__17658),
            .I(data_in_field_55));
    Odrv4 I__2793 (
            .O(N__17655),
            .I(data_in_field_55));
    LocalMux I__2792 (
            .O(N__17652),
            .I(data_in_field_55));
    InMux I__2791 (
            .O(N__17643),
            .I(N__17640));
    LocalMux I__2790 (
            .O(N__17640),
            .I(\c0.n6_adj_1636 ));
    CascadeMux I__2789 (
            .O(N__17637),
            .I(N__17633));
    CascadeMux I__2788 (
            .O(N__17636),
            .I(N__17630));
    InMux I__2787 (
            .O(N__17633),
            .I(N__17627));
    InMux I__2786 (
            .O(N__17630),
            .I(N__17624));
    LocalMux I__2785 (
            .O(N__17627),
            .I(N__17621));
    LocalMux I__2784 (
            .O(N__17624),
            .I(N__17618));
    Span4Mux_h I__2783 (
            .O(N__17621),
            .I(N__17615));
    Span12Mux_v I__2782 (
            .O(N__17618),
            .I(N__17612));
    Span4Mux_h I__2781 (
            .O(N__17615),
            .I(N__17609));
    Odrv12 I__2780 (
            .O(N__17612),
            .I(\c0.n8989 ));
    Odrv4 I__2779 (
            .O(N__17609),
            .I(\c0.n8989 ));
    InMux I__2778 (
            .O(N__17604),
            .I(N__17599));
    CascadeMux I__2777 (
            .O(N__17603),
            .I(N__17596));
    InMux I__2776 (
            .O(N__17602),
            .I(N__17590));
    LocalMux I__2775 (
            .O(N__17599),
            .I(N__17586));
    InMux I__2774 (
            .O(N__17596),
            .I(N__17583));
    InMux I__2773 (
            .O(N__17595),
            .I(N__17580));
    InMux I__2772 (
            .O(N__17594),
            .I(N__17577));
    InMux I__2771 (
            .O(N__17593),
            .I(N__17574));
    LocalMux I__2770 (
            .O(N__17590),
            .I(N__17571));
    InMux I__2769 (
            .O(N__17589),
            .I(N__17568));
    Span4Mux_s2_v I__2768 (
            .O(N__17586),
            .I(N__17563));
    LocalMux I__2767 (
            .O(N__17583),
            .I(N__17563));
    LocalMux I__2766 (
            .O(N__17580),
            .I(data_in_field_63));
    LocalMux I__2765 (
            .O(N__17577),
            .I(data_in_field_63));
    LocalMux I__2764 (
            .O(N__17574),
            .I(data_in_field_63));
    Odrv12 I__2763 (
            .O(N__17571),
            .I(data_in_field_63));
    LocalMux I__2762 (
            .O(N__17568),
            .I(data_in_field_63));
    Odrv4 I__2761 (
            .O(N__17563),
            .I(data_in_field_63));
    CascadeMux I__2760 (
            .O(N__17550),
            .I(N__17546));
    CascadeMux I__2759 (
            .O(N__17549),
            .I(N__17543));
    InMux I__2758 (
            .O(N__17546),
            .I(N__17537));
    InMux I__2757 (
            .O(N__17543),
            .I(N__17534));
    InMux I__2756 (
            .O(N__17542),
            .I(N__17527));
    InMux I__2755 (
            .O(N__17541),
            .I(N__17527));
    InMux I__2754 (
            .O(N__17540),
            .I(N__17527));
    LocalMux I__2753 (
            .O(N__17537),
            .I(N__17524));
    LocalMux I__2752 (
            .O(N__17534),
            .I(N__17521));
    LocalMux I__2751 (
            .O(N__17527),
            .I(N__17514));
    Span4Mux_h I__2750 (
            .O(N__17524),
            .I(N__17514));
    Span4Mux_s3_h I__2749 (
            .O(N__17521),
            .I(N__17514));
    Odrv4 I__2748 (
            .O(N__17514),
            .I(data_in_field_59));
    InMux I__2747 (
            .O(N__17511),
            .I(N__17507));
    InMux I__2746 (
            .O(N__17510),
            .I(N__17504));
    LocalMux I__2745 (
            .O(N__17507),
            .I(N__17498));
    LocalMux I__2744 (
            .O(N__17504),
            .I(N__17495));
    InMux I__2743 (
            .O(N__17503),
            .I(N__17490));
    InMux I__2742 (
            .O(N__17502),
            .I(N__17490));
    InMux I__2741 (
            .O(N__17501),
            .I(N__17487));
    Span4Mux_v I__2740 (
            .O(N__17498),
            .I(N__17484));
    Span4Mux_v I__2739 (
            .O(N__17495),
            .I(N__17479));
    LocalMux I__2738 (
            .O(N__17490),
            .I(N__17479));
    LocalMux I__2737 (
            .O(N__17487),
            .I(data_in_field_51));
    Odrv4 I__2736 (
            .O(N__17484),
            .I(data_in_field_51));
    Odrv4 I__2735 (
            .O(N__17479),
            .I(data_in_field_51));
    InMux I__2734 (
            .O(N__17472),
            .I(N__17469));
    LocalMux I__2733 (
            .O(N__17469),
            .I(N__17465));
    InMux I__2732 (
            .O(N__17468),
            .I(N__17462));
    Span4Mux_v I__2731 (
            .O(N__17465),
            .I(N__17457));
    LocalMux I__2730 (
            .O(N__17462),
            .I(N__17457));
    Span4Mux_h I__2729 (
            .O(N__17457),
            .I(N__17454));
    Odrv4 I__2728 (
            .O(N__17454),
            .I(\c0.n4302 ));
    CascadeMux I__2727 (
            .O(N__17451),
            .I(N__17447));
    InMux I__2726 (
            .O(N__17450),
            .I(N__17443));
    InMux I__2725 (
            .O(N__17447),
            .I(N__17440));
    InMux I__2724 (
            .O(N__17446),
            .I(N__17437));
    LocalMux I__2723 (
            .O(N__17443),
            .I(N__17432));
    LocalMux I__2722 (
            .O(N__17440),
            .I(N__17429));
    LocalMux I__2721 (
            .O(N__17437),
            .I(N__17426));
    InMux I__2720 (
            .O(N__17436),
            .I(N__17423));
    InMux I__2719 (
            .O(N__17435),
            .I(N__17420));
    Span4Mux_v I__2718 (
            .O(N__17432),
            .I(N__17413));
    Span4Mux_s3_v I__2717 (
            .O(N__17429),
            .I(N__17413));
    Span4Mux_s3_v I__2716 (
            .O(N__17426),
            .I(N__17413));
    LocalMux I__2715 (
            .O(N__17423),
            .I(data_in_field_79));
    LocalMux I__2714 (
            .O(N__17420),
            .I(data_in_field_79));
    Odrv4 I__2713 (
            .O(N__17413),
            .I(data_in_field_79));
    InMux I__2712 (
            .O(N__17406),
            .I(N__17403));
    LocalMux I__2711 (
            .O(N__17403),
            .I(N__17399));
    CascadeMux I__2710 (
            .O(N__17402),
            .I(N__17395));
    Span4Mux_v I__2709 (
            .O(N__17399),
            .I(N__17390));
    InMux I__2708 (
            .O(N__17398),
            .I(N__17387));
    InMux I__2707 (
            .O(N__17395),
            .I(N__17384));
    InMux I__2706 (
            .O(N__17394),
            .I(N__17381));
    InMux I__2705 (
            .O(N__17393),
            .I(N__17378));
    Span4Mux_h I__2704 (
            .O(N__17390),
            .I(N__17375));
    LocalMux I__2703 (
            .O(N__17387),
            .I(N__17372));
    LocalMux I__2702 (
            .O(N__17384),
            .I(N__17369));
    LocalMux I__2701 (
            .O(N__17381),
            .I(data_in_field_139));
    LocalMux I__2700 (
            .O(N__17378),
            .I(data_in_field_139));
    Odrv4 I__2699 (
            .O(N__17375),
            .I(data_in_field_139));
    Odrv12 I__2698 (
            .O(N__17372),
            .I(data_in_field_139));
    Odrv12 I__2697 (
            .O(N__17369),
            .I(data_in_field_139));
    InMux I__2696 (
            .O(N__17358),
            .I(N__17354));
    InMux I__2695 (
            .O(N__17357),
            .I(N__17351));
    LocalMux I__2694 (
            .O(N__17354),
            .I(N__17348));
    LocalMux I__2693 (
            .O(N__17351),
            .I(N__17343));
    Span4Mux_h I__2692 (
            .O(N__17348),
            .I(N__17343));
    Odrv4 I__2691 (
            .O(N__17343),
            .I(\c0.n8825 ));
    InMux I__2690 (
            .O(N__17340),
            .I(N__17337));
    LocalMux I__2689 (
            .O(N__17337),
            .I(N__17334));
    Odrv12 I__2688 (
            .O(N__17334),
            .I(\c0.n6_adj_1654 ));
    InMux I__2687 (
            .O(N__17331),
            .I(N__17328));
    LocalMux I__2686 (
            .O(N__17328),
            .I(\c0.n4253 ));
    CascadeMux I__2685 (
            .O(N__17325),
            .I(N__17322));
    InMux I__2684 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__2683 (
            .O(N__17319),
            .I(N__17316));
    Odrv12 I__2682 (
            .O(N__17316),
            .I(\c0.n4151 ));
    InMux I__2681 (
            .O(N__17313),
            .I(N__17306));
    InMux I__2680 (
            .O(N__17312),
            .I(N__17306));
    InMux I__2679 (
            .O(N__17311),
            .I(N__17301));
    LocalMux I__2678 (
            .O(N__17306),
            .I(N__17298));
    InMux I__2677 (
            .O(N__17305),
            .I(N__17295));
    InMux I__2676 (
            .O(N__17304),
            .I(N__17292));
    LocalMux I__2675 (
            .O(N__17301),
            .I(N__17289));
    Span4Mux_h I__2674 (
            .O(N__17298),
            .I(N__17286));
    LocalMux I__2673 (
            .O(N__17295),
            .I(N__17283));
    LocalMux I__2672 (
            .O(N__17292),
            .I(\c0.data_in_field_17 ));
    Odrv12 I__2671 (
            .O(N__17289),
            .I(\c0.data_in_field_17 ));
    Odrv4 I__2670 (
            .O(N__17286),
            .I(\c0.data_in_field_17 ));
    Odrv12 I__2669 (
            .O(N__17283),
            .I(\c0.data_in_field_17 ));
    InMux I__2668 (
            .O(N__17274),
            .I(N__17271));
    LocalMux I__2667 (
            .O(N__17271),
            .I(N__17268));
    Odrv12 I__2666 (
            .O(N__17268),
            .I(\c0.n45 ));
    CascadeMux I__2665 (
            .O(N__17265),
            .I(N__17262));
    InMux I__2664 (
            .O(N__17262),
            .I(N__17258));
    InMux I__2663 (
            .O(N__17261),
            .I(N__17255));
    LocalMux I__2662 (
            .O(N__17258),
            .I(N__17251));
    LocalMux I__2661 (
            .O(N__17255),
            .I(N__17248));
    InMux I__2660 (
            .O(N__17254),
            .I(N__17245));
    Span4Mux_v I__2659 (
            .O(N__17251),
            .I(N__17242));
    Odrv4 I__2658 (
            .O(N__17248),
            .I(\c0.n4183 ));
    LocalMux I__2657 (
            .O(N__17245),
            .I(\c0.n4183 ));
    Odrv4 I__2656 (
            .O(N__17242),
            .I(\c0.n4183 ));
    InMux I__2655 (
            .O(N__17235),
            .I(N__17232));
    LocalMux I__2654 (
            .O(N__17232),
            .I(N__17229));
    Span4Mux_h I__2653 (
            .O(N__17229),
            .I(N__17225));
    InMux I__2652 (
            .O(N__17228),
            .I(N__17222));
    Odrv4 I__2651 (
            .O(N__17225),
            .I(\c0.n8864 ));
    LocalMux I__2650 (
            .O(N__17222),
            .I(\c0.n8864 ));
    CascadeMux I__2649 (
            .O(N__17217),
            .I(N__17214));
    InMux I__2648 (
            .O(N__17214),
            .I(N__17211));
    LocalMux I__2647 (
            .O(N__17211),
            .I(N__17208));
    Odrv12 I__2646 (
            .O(N__17208),
            .I(\c0.n8843 ));
    InMux I__2645 (
            .O(N__17205),
            .I(N__17201));
    InMux I__2644 (
            .O(N__17204),
            .I(N__17198));
    LocalMux I__2643 (
            .O(N__17201),
            .I(N__17195));
    LocalMux I__2642 (
            .O(N__17198),
            .I(\c0.n8930 ));
    Odrv12 I__2641 (
            .O(N__17195),
            .I(\c0.n8930 ));
    InMux I__2640 (
            .O(N__17190),
            .I(N__17187));
    LocalMux I__2639 (
            .O(N__17187),
            .I(N__17184));
    Span4Mux_h I__2638 (
            .O(N__17184),
            .I(N__17181));
    Odrv4 I__2637 (
            .O(N__17181),
            .I(\c0.n20 ));
    CascadeMux I__2636 (
            .O(N__17178),
            .I(\c0.n21_cascade_ ));
    InMux I__2635 (
            .O(N__17175),
            .I(N__17172));
    LocalMux I__2634 (
            .O(N__17172),
            .I(N__17169));
    Span4Mux_v I__2633 (
            .O(N__17169),
            .I(N__17166));
    Odrv4 I__2632 (
            .O(N__17166),
            .I(\c0.n19 ));
    InMux I__2631 (
            .O(N__17163),
            .I(N__17160));
    LocalMux I__2630 (
            .O(N__17160),
            .I(\c0.n18 ));
    CascadeMux I__2629 (
            .O(N__17157),
            .I(\c0.n8421_cascade_ ));
    InMux I__2628 (
            .O(N__17154),
            .I(N__17150));
    InMux I__2627 (
            .O(N__17153),
            .I(N__17147));
    LocalMux I__2626 (
            .O(N__17150),
            .I(N__17144));
    LocalMux I__2625 (
            .O(N__17147),
            .I(N__17141));
    Odrv4 I__2624 (
            .O(N__17144),
            .I(\c0.tx2_transmit_N_1334 ));
    Odrv4 I__2623 (
            .O(N__17141),
            .I(\c0.tx2_transmit_N_1334 ));
    InMux I__2622 (
            .O(N__17136),
            .I(N__17133));
    LocalMux I__2621 (
            .O(N__17133),
            .I(\c0.n24_adj_1605 ));
    InMux I__2620 (
            .O(N__17130),
            .I(N__17127));
    LocalMux I__2619 (
            .O(N__17127),
            .I(N__17121));
    InMux I__2618 (
            .O(N__17126),
            .I(N__17118));
    InMux I__2617 (
            .O(N__17125),
            .I(N__17113));
    InMux I__2616 (
            .O(N__17124),
            .I(N__17113));
    Span12Mux_s5_v I__2615 (
            .O(N__17121),
            .I(N__17110));
    LocalMux I__2614 (
            .O(N__17118),
            .I(data_in_field_75));
    LocalMux I__2613 (
            .O(N__17113),
            .I(data_in_field_75));
    Odrv12 I__2612 (
            .O(N__17110),
            .I(data_in_field_75));
    InMux I__2611 (
            .O(N__17103),
            .I(N__17100));
    LocalMux I__2610 (
            .O(N__17100),
            .I(N__17094));
    InMux I__2609 (
            .O(N__17099),
            .I(N__17089));
    InMux I__2608 (
            .O(N__17098),
            .I(N__17089));
    InMux I__2607 (
            .O(N__17097),
            .I(N__17086));
    Span4Mux_v I__2606 (
            .O(N__17094),
            .I(N__17083));
    LocalMux I__2605 (
            .O(N__17089),
            .I(N__17080));
    LocalMux I__2604 (
            .O(N__17086),
            .I(data_in_field_67));
    Odrv4 I__2603 (
            .O(N__17083),
            .I(data_in_field_67));
    Odrv12 I__2602 (
            .O(N__17080),
            .I(data_in_field_67));
    CascadeMux I__2601 (
            .O(N__17073),
            .I(\c0.n9506_cascade_ ));
    InMux I__2600 (
            .O(N__17070),
            .I(N__17064));
    InMux I__2599 (
            .O(N__17069),
            .I(N__17061));
    InMux I__2598 (
            .O(N__17068),
            .I(N__17058));
    InMux I__2597 (
            .O(N__17067),
            .I(N__17054));
    LocalMux I__2596 (
            .O(N__17064),
            .I(N__17051));
    LocalMux I__2595 (
            .O(N__17061),
            .I(N__17046));
    LocalMux I__2594 (
            .O(N__17058),
            .I(N__17046));
    InMux I__2593 (
            .O(N__17057),
            .I(N__17043));
    LocalMux I__2592 (
            .O(N__17054),
            .I(\c0.data_in_field_34 ));
    Odrv4 I__2591 (
            .O(N__17051),
            .I(\c0.data_in_field_34 ));
    Odrv4 I__2590 (
            .O(N__17046),
            .I(\c0.data_in_field_34 ));
    LocalMux I__2589 (
            .O(N__17043),
            .I(\c0.data_in_field_34 ));
    CascadeMux I__2588 (
            .O(N__17034),
            .I(\c0.n4_adj_1592_cascade_ ));
    InMux I__2587 (
            .O(N__17031),
            .I(N__17028));
    LocalMux I__2586 (
            .O(N__17028),
            .I(N__17025));
    Span4Mux_h I__2585 (
            .O(N__17025),
            .I(N__17022));
    Odrv4 I__2584 (
            .O(N__17022),
            .I(\c0.n4324 ));
    InMux I__2583 (
            .O(N__17019),
            .I(N__17016));
    LocalMux I__2582 (
            .O(N__17016),
            .I(\c0.n21_adj_1599 ));
    InMux I__2581 (
            .O(N__17013),
            .I(N__17010));
    LocalMux I__2580 (
            .O(N__17010),
            .I(N__17007));
    Span4Mux_v I__2579 (
            .O(N__17007),
            .I(N__17003));
    InMux I__2578 (
            .O(N__17006),
            .I(N__17000));
    Odrv4 I__2577 (
            .O(N__17003),
            .I(\c0.n4200 ));
    LocalMux I__2576 (
            .O(N__17000),
            .I(\c0.n4200 ));
    CascadeMux I__2575 (
            .O(N__16995),
            .I(N__16992));
    InMux I__2574 (
            .O(N__16992),
            .I(N__16989));
    LocalMux I__2573 (
            .O(N__16989),
            .I(\c0.n28 ));
    InMux I__2572 (
            .O(N__16986),
            .I(N__16983));
    LocalMux I__2571 (
            .O(N__16983),
            .I(\c0.n23_adj_1608 ));
    InMux I__2570 (
            .O(N__16980),
            .I(N__16977));
    LocalMux I__2569 (
            .O(N__16977),
            .I(N__16974));
    Span4Mux_h I__2568 (
            .O(N__16974),
            .I(N__16968));
    InMux I__2567 (
            .O(N__16973),
            .I(N__16963));
    InMux I__2566 (
            .O(N__16972),
            .I(N__16963));
    InMux I__2565 (
            .O(N__16971),
            .I(N__16960));
    Odrv4 I__2564 (
            .O(N__16968),
            .I(data_in_1_7));
    LocalMux I__2563 (
            .O(N__16963),
            .I(data_in_1_7));
    LocalMux I__2562 (
            .O(N__16960),
            .I(data_in_1_7));
    InMux I__2561 (
            .O(N__16953),
            .I(N__16950));
    LocalMux I__2560 (
            .O(N__16950),
            .I(N__16947));
    Span4Mux_v I__2559 (
            .O(N__16947),
            .I(N__16942));
    InMux I__2558 (
            .O(N__16946),
            .I(N__16937));
    InMux I__2557 (
            .O(N__16945),
            .I(N__16937));
    Odrv4 I__2556 (
            .O(N__16942),
            .I(\c0.data_in_field_15 ));
    LocalMux I__2555 (
            .O(N__16937),
            .I(\c0.data_in_field_15 ));
    CascadeMux I__2554 (
            .O(N__16932),
            .I(n1895_cascade_));
    InMux I__2553 (
            .O(N__16929),
            .I(N__16926));
    LocalMux I__2552 (
            .O(N__16926),
            .I(N__16923));
    Odrv4 I__2551 (
            .O(N__16923),
            .I(n1889));
    InMux I__2550 (
            .O(N__16920),
            .I(N__16917));
    LocalMux I__2549 (
            .O(N__16917),
            .I(N__16914));
    Span4Mux_h I__2548 (
            .O(N__16914),
            .I(N__16911));
    Odrv4 I__2547 (
            .O(N__16911),
            .I(n1897));
    InMux I__2546 (
            .O(N__16908),
            .I(N__16904));
    InMux I__2545 (
            .O(N__16907),
            .I(N__16901));
    LocalMux I__2544 (
            .O(N__16904),
            .I(N__16897));
    LocalMux I__2543 (
            .O(N__16901),
            .I(N__16894));
    InMux I__2542 (
            .O(N__16900),
            .I(N__16891));
    Odrv12 I__2541 (
            .O(N__16897),
            .I(data_in_4_4));
    Odrv4 I__2540 (
            .O(N__16894),
            .I(data_in_4_4));
    LocalMux I__2539 (
            .O(N__16891),
            .I(data_in_4_4));
    CascadeMux I__2538 (
            .O(N__16884),
            .I(N__16880));
    InMux I__2537 (
            .O(N__16883),
            .I(N__16875));
    InMux I__2536 (
            .O(N__16880),
            .I(N__16872));
    CascadeMux I__2535 (
            .O(N__16879),
            .I(N__16869));
    InMux I__2534 (
            .O(N__16878),
            .I(N__16866));
    LocalMux I__2533 (
            .O(N__16875),
            .I(N__16863));
    LocalMux I__2532 (
            .O(N__16872),
            .I(N__16860));
    InMux I__2531 (
            .O(N__16869),
            .I(N__16857));
    LocalMux I__2530 (
            .O(N__16866),
            .I(data_in_2_0));
    Odrv4 I__2529 (
            .O(N__16863),
            .I(data_in_2_0));
    Odrv12 I__2528 (
            .O(N__16860),
            .I(data_in_2_0));
    LocalMux I__2527 (
            .O(N__16857),
            .I(data_in_2_0));
    InMux I__2526 (
            .O(N__16848),
            .I(N__16843));
    InMux I__2525 (
            .O(N__16847),
            .I(N__16840));
    InMux I__2524 (
            .O(N__16846),
            .I(N__16836));
    LocalMux I__2523 (
            .O(N__16843),
            .I(N__16833));
    LocalMux I__2522 (
            .O(N__16840),
            .I(N__16830));
    InMux I__2521 (
            .O(N__16839),
            .I(N__16827));
    LocalMux I__2520 (
            .O(N__16836),
            .I(\c0.data_in_field_26 ));
    Odrv4 I__2519 (
            .O(N__16833),
            .I(\c0.data_in_field_26 ));
    Odrv4 I__2518 (
            .O(N__16830),
            .I(\c0.data_in_field_26 ));
    LocalMux I__2517 (
            .O(N__16827),
            .I(\c0.data_in_field_26 ));
    CascadeMux I__2516 (
            .O(N__16818),
            .I(N__16813));
    CascadeMux I__2515 (
            .O(N__16817),
            .I(N__16810));
    InMux I__2514 (
            .O(N__16816),
            .I(N__16807));
    InMux I__2513 (
            .O(N__16813),
            .I(N__16802));
    InMux I__2512 (
            .O(N__16810),
            .I(N__16799));
    LocalMux I__2511 (
            .O(N__16807),
            .I(N__16796));
    InMux I__2510 (
            .O(N__16806),
            .I(N__16793));
    InMux I__2509 (
            .O(N__16805),
            .I(N__16790));
    LocalMux I__2508 (
            .O(N__16802),
            .I(\c0.data_in_field_18 ));
    LocalMux I__2507 (
            .O(N__16799),
            .I(\c0.data_in_field_18 ));
    Odrv4 I__2506 (
            .O(N__16796),
            .I(\c0.data_in_field_18 ));
    LocalMux I__2505 (
            .O(N__16793),
            .I(\c0.data_in_field_18 ));
    LocalMux I__2504 (
            .O(N__16790),
            .I(\c0.data_in_field_18 ));
    CascadeMux I__2503 (
            .O(N__16779),
            .I(N__16776));
    InMux I__2502 (
            .O(N__16776),
            .I(N__16773));
    LocalMux I__2501 (
            .O(N__16773),
            .I(N__16770));
    Span12Mux_s4_h I__2500 (
            .O(N__16770),
            .I(N__16767));
    Odrv12 I__2499 (
            .O(N__16767),
            .I(\c0.n9512 ));
    InMux I__2498 (
            .O(N__16764),
            .I(N__16761));
    LocalMux I__2497 (
            .O(N__16761),
            .I(N__16757));
    InMux I__2496 (
            .O(N__16760),
            .I(N__16754));
    Span4Mux_v I__2495 (
            .O(N__16757),
            .I(N__16751));
    LocalMux I__2494 (
            .O(N__16754),
            .I(N__16746));
    Span4Mux_h I__2493 (
            .O(N__16751),
            .I(N__16743));
    InMux I__2492 (
            .O(N__16750),
            .I(N__16738));
    InMux I__2491 (
            .O(N__16749),
            .I(N__16738));
    Span4Mux_h I__2490 (
            .O(N__16746),
            .I(N__16735));
    Odrv4 I__2489 (
            .O(N__16743),
            .I(data_in_2_1));
    LocalMux I__2488 (
            .O(N__16738),
            .I(data_in_2_1));
    Odrv4 I__2487 (
            .O(N__16735),
            .I(data_in_2_1));
    InMux I__2486 (
            .O(N__16728),
            .I(N__16725));
    LocalMux I__2485 (
            .O(N__16725),
            .I(N__16722));
    Span4Mux_h I__2484 (
            .O(N__16722),
            .I(N__16719));
    Odrv4 I__2483 (
            .O(N__16719),
            .I(\c0.n4492 ));
    InMux I__2482 (
            .O(N__16716),
            .I(N__16713));
    LocalMux I__2481 (
            .O(N__16713),
            .I(N__16709));
    InMux I__2480 (
            .O(N__16712),
            .I(N__16706));
    Span4Mux_h I__2479 (
            .O(N__16709),
            .I(N__16703));
    LocalMux I__2478 (
            .O(N__16706),
            .I(\c0.n24 ));
    Odrv4 I__2477 (
            .O(N__16703),
            .I(\c0.n24 ));
    InMux I__2476 (
            .O(N__16698),
            .I(N__16694));
    InMux I__2475 (
            .O(N__16697),
            .I(N__16691));
    LocalMux I__2474 (
            .O(N__16694),
            .I(\c0.n8902 ));
    LocalMux I__2473 (
            .O(N__16691),
            .I(\c0.n8902 ));
    CascadeMux I__2472 (
            .O(N__16686),
            .I(\c0.n4492_cascade_ ));
    CascadeMux I__2471 (
            .O(N__16683),
            .I(\c0.n8948_cascade_ ));
    InMux I__2470 (
            .O(N__16680),
            .I(N__16677));
    LocalMux I__2469 (
            .O(N__16677),
            .I(N__16673));
    InMux I__2468 (
            .O(N__16676),
            .I(N__16670));
    Span4Mux_v I__2467 (
            .O(N__16673),
            .I(N__16667));
    LocalMux I__2466 (
            .O(N__16670),
            .I(N__16664));
    Odrv4 I__2465 (
            .O(N__16667),
            .I(\c0.n8858 ));
    Odrv12 I__2464 (
            .O(N__16664),
            .I(\c0.n8858 ));
    CascadeMux I__2463 (
            .O(N__16659),
            .I(N__16656));
    InMux I__2462 (
            .O(N__16656),
            .I(N__16653));
    LocalMux I__2461 (
            .O(N__16653),
            .I(\c0.n19_adj_1602 ));
    InMux I__2460 (
            .O(N__16650),
            .I(N__16647));
    LocalMux I__2459 (
            .O(N__16647),
            .I(N__16643));
    InMux I__2458 (
            .O(N__16646),
            .I(N__16639));
    Span4Mux_h I__2457 (
            .O(N__16643),
            .I(N__16636));
    InMux I__2456 (
            .O(N__16642),
            .I(N__16633));
    LocalMux I__2455 (
            .O(N__16639),
            .I(data_in_0_1));
    Odrv4 I__2454 (
            .O(N__16636),
            .I(data_in_0_1));
    LocalMux I__2453 (
            .O(N__16633),
            .I(data_in_0_1));
    InMux I__2452 (
            .O(N__16626),
            .I(N__16623));
    LocalMux I__2451 (
            .O(N__16623),
            .I(N__16620));
    Span4Mux_h I__2450 (
            .O(N__16620),
            .I(N__16617));
    Span4Mux_h I__2449 (
            .O(N__16617),
            .I(N__16611));
    InMux I__2448 (
            .O(N__16616),
            .I(N__16608));
    InMux I__2447 (
            .O(N__16615),
            .I(N__16603));
    InMux I__2446 (
            .O(N__16614),
            .I(N__16603));
    Odrv4 I__2445 (
            .O(N__16611),
            .I(\c0.data_in_field_1 ));
    LocalMux I__2444 (
            .O(N__16608),
            .I(\c0.data_in_field_1 ));
    LocalMux I__2443 (
            .O(N__16603),
            .I(\c0.data_in_field_1 ));
    InMux I__2442 (
            .O(N__16596),
            .I(N__16587));
    InMux I__2441 (
            .O(N__16595),
            .I(N__16587));
    InMux I__2440 (
            .O(N__16594),
            .I(N__16587));
    LocalMux I__2439 (
            .O(N__16587),
            .I(data_in_6_6));
    InMux I__2438 (
            .O(N__16584),
            .I(N__16581));
    LocalMux I__2437 (
            .O(N__16581),
            .I(N__16577));
    InMux I__2436 (
            .O(N__16580),
            .I(N__16574));
    Span4Mux_h I__2435 (
            .O(N__16577),
            .I(N__16571));
    LocalMux I__2434 (
            .O(N__16574),
            .I(data_in_8_6));
    Odrv4 I__2433 (
            .O(N__16571),
            .I(data_in_8_6));
    CascadeMux I__2432 (
            .O(N__16566),
            .I(N__16563));
    InMux I__2431 (
            .O(N__16563),
            .I(N__16557));
    InMux I__2430 (
            .O(N__16562),
            .I(N__16557));
    LocalMux I__2429 (
            .O(N__16557),
            .I(data_in_7_6));
    InMux I__2428 (
            .O(N__16554),
            .I(N__16551));
    LocalMux I__2427 (
            .O(N__16551),
            .I(N__16548));
    Span4Mux_h I__2426 (
            .O(N__16548),
            .I(N__16545));
    Span4Mux_v I__2425 (
            .O(N__16545),
            .I(N__16539));
    InMux I__2424 (
            .O(N__16544),
            .I(N__16534));
    InMux I__2423 (
            .O(N__16543),
            .I(N__16534));
    InMux I__2422 (
            .O(N__16542),
            .I(N__16531));
    Odrv4 I__2421 (
            .O(N__16539),
            .I(data_in_3_5));
    LocalMux I__2420 (
            .O(N__16534),
            .I(data_in_3_5));
    LocalMux I__2419 (
            .O(N__16531),
            .I(data_in_3_5));
    CascadeMux I__2418 (
            .O(N__16524),
            .I(N__16521));
    InMux I__2417 (
            .O(N__16521),
            .I(N__16515));
    InMux I__2416 (
            .O(N__16520),
            .I(N__16508));
    InMux I__2415 (
            .O(N__16519),
            .I(N__16508));
    InMux I__2414 (
            .O(N__16518),
            .I(N__16508));
    LocalMux I__2413 (
            .O(N__16515),
            .I(data_in_3_6));
    LocalMux I__2412 (
            .O(N__16508),
            .I(data_in_3_6));
    CascadeMux I__2411 (
            .O(N__16503),
            .I(\c0.n8843_cascade_ ));
    InMux I__2410 (
            .O(N__16500),
            .I(N__16497));
    LocalMux I__2409 (
            .O(N__16497),
            .I(N__16493));
    InMux I__2408 (
            .O(N__16496),
            .I(N__16490));
    Span4Mux_v I__2407 (
            .O(N__16493),
            .I(N__16484));
    LocalMux I__2406 (
            .O(N__16490),
            .I(N__16481));
    InMux I__2405 (
            .O(N__16489),
            .I(N__16478));
    InMux I__2404 (
            .O(N__16488),
            .I(N__16473));
    InMux I__2403 (
            .O(N__16487),
            .I(N__16473));
    Odrv4 I__2402 (
            .O(N__16484),
            .I(\c0.data_in_field_31 ));
    Odrv4 I__2401 (
            .O(N__16481),
            .I(\c0.data_in_field_31 ));
    LocalMux I__2400 (
            .O(N__16478),
            .I(\c0.data_in_field_31 ));
    LocalMux I__2399 (
            .O(N__16473),
            .I(\c0.data_in_field_31 ));
    CascadeMux I__2398 (
            .O(N__16464),
            .I(\c0.n4151_cascade_ ));
    InMux I__2397 (
            .O(N__16461),
            .I(N__16451));
    InMux I__2396 (
            .O(N__16460),
            .I(N__16451));
    InMux I__2395 (
            .O(N__16459),
            .I(N__16451));
    InMux I__2394 (
            .O(N__16458),
            .I(N__16448));
    LocalMux I__2393 (
            .O(N__16451),
            .I(\c0.data_in_field_30 ));
    LocalMux I__2392 (
            .O(N__16448),
            .I(\c0.data_in_field_30 ));
    InMux I__2391 (
            .O(N__16443),
            .I(N__16440));
    LocalMux I__2390 (
            .O(N__16440),
            .I(N__16436));
    InMux I__2389 (
            .O(N__16439),
            .I(N__16431));
    Span4Mux_h I__2388 (
            .O(N__16436),
            .I(N__16428));
    InMux I__2387 (
            .O(N__16435),
            .I(N__16425));
    InMux I__2386 (
            .O(N__16434),
            .I(N__16422));
    LocalMux I__2385 (
            .O(N__16431),
            .I(\c0.data_in_field_22 ));
    Odrv4 I__2384 (
            .O(N__16428),
            .I(\c0.data_in_field_22 ));
    LocalMux I__2383 (
            .O(N__16425),
            .I(\c0.data_in_field_22 ));
    LocalMux I__2382 (
            .O(N__16422),
            .I(\c0.data_in_field_22 ));
    CascadeMux I__2381 (
            .O(N__16413),
            .I(N__16408));
    InMux I__2380 (
            .O(N__16412),
            .I(N__16405));
    CascadeMux I__2379 (
            .O(N__16411),
            .I(N__16401));
    InMux I__2378 (
            .O(N__16408),
            .I(N__16398));
    LocalMux I__2377 (
            .O(N__16405),
            .I(N__16395));
    InMux I__2376 (
            .O(N__16404),
            .I(N__16390));
    InMux I__2375 (
            .O(N__16401),
            .I(N__16390));
    LocalMux I__2374 (
            .O(N__16398),
            .I(\c0.data_in_field_14 ));
    Odrv4 I__2373 (
            .O(N__16395),
            .I(\c0.data_in_field_14 ));
    LocalMux I__2372 (
            .O(N__16390),
            .I(\c0.data_in_field_14 ));
    CascadeMux I__2371 (
            .O(N__16383),
            .I(\c0.n9638_cascade_ ));
    InMux I__2370 (
            .O(N__16380),
            .I(N__16375));
    InMux I__2369 (
            .O(N__16379),
            .I(N__16372));
    CascadeMux I__2368 (
            .O(N__16378),
            .I(N__16368));
    LocalMux I__2367 (
            .O(N__16375),
            .I(N__16365));
    LocalMux I__2366 (
            .O(N__16372),
            .I(N__16362));
    InMux I__2365 (
            .O(N__16371),
            .I(N__16359));
    InMux I__2364 (
            .O(N__16368),
            .I(N__16355));
    Span4Mux_h I__2363 (
            .O(N__16365),
            .I(N__16352));
    Span4Mux_v I__2362 (
            .O(N__16362),
            .I(N__16347));
    LocalMux I__2361 (
            .O(N__16359),
            .I(N__16347));
    InMux I__2360 (
            .O(N__16358),
            .I(N__16344));
    LocalMux I__2359 (
            .O(N__16355),
            .I(\c0.data_in_field_6 ));
    Odrv4 I__2358 (
            .O(N__16352),
            .I(\c0.data_in_field_6 ));
    Odrv4 I__2357 (
            .O(N__16347),
            .I(\c0.data_in_field_6 ));
    LocalMux I__2356 (
            .O(N__16344),
            .I(\c0.data_in_field_6 ));
    InMux I__2355 (
            .O(N__16335),
            .I(N__16332));
    LocalMux I__2354 (
            .O(N__16332),
            .I(N__16329));
    Span4Mux_v I__2353 (
            .O(N__16329),
            .I(N__16325));
    InMux I__2352 (
            .O(N__16328),
            .I(N__16322));
    Odrv4 I__2351 (
            .O(N__16325),
            .I(data_in_15_4));
    LocalMux I__2350 (
            .O(N__16322),
            .I(data_in_15_4));
    InMux I__2349 (
            .O(N__16317),
            .I(N__16313));
    InMux I__2348 (
            .O(N__16316),
            .I(N__16310));
    LocalMux I__2347 (
            .O(N__16313),
            .I(data_in_17_4));
    LocalMux I__2346 (
            .O(N__16310),
            .I(data_in_17_4));
    InMux I__2345 (
            .O(N__16305),
            .I(N__16299));
    InMux I__2344 (
            .O(N__16304),
            .I(N__16299));
    LocalMux I__2343 (
            .O(N__16299),
            .I(data_in_16_4));
    InMux I__2342 (
            .O(N__16296),
            .I(N__16290));
    InMux I__2341 (
            .O(N__16295),
            .I(N__16290));
    LocalMux I__2340 (
            .O(N__16290),
            .I(data_in_17_7));
    InMux I__2339 (
            .O(N__16287),
            .I(N__16283));
    InMux I__2338 (
            .O(N__16286),
            .I(N__16280));
    LocalMux I__2337 (
            .O(N__16283),
            .I(data_in_19_4));
    LocalMux I__2336 (
            .O(N__16280),
            .I(data_in_19_4));
    InMux I__2335 (
            .O(N__16275),
            .I(N__16271));
    InMux I__2334 (
            .O(N__16274),
            .I(N__16268));
    LocalMux I__2333 (
            .O(N__16271),
            .I(data_in_18_4));
    LocalMux I__2332 (
            .O(N__16268),
            .I(data_in_18_4));
    CascadeMux I__2331 (
            .O(N__16263),
            .I(N__16259));
    InMux I__2330 (
            .O(N__16262),
            .I(N__16256));
    InMux I__2329 (
            .O(N__16259),
            .I(N__16251));
    LocalMux I__2328 (
            .O(N__16256),
            .I(N__16248));
    CascadeMux I__2327 (
            .O(N__16255),
            .I(N__16245));
    InMux I__2326 (
            .O(N__16254),
            .I(N__16242));
    LocalMux I__2325 (
            .O(N__16251),
            .I(N__16239));
    Span4Mux_h I__2324 (
            .O(N__16248),
            .I(N__16236));
    InMux I__2323 (
            .O(N__16245),
            .I(N__16233));
    LocalMux I__2322 (
            .O(N__16242),
            .I(data_in_2_5));
    Odrv4 I__2321 (
            .O(N__16239),
            .I(data_in_2_5));
    Odrv4 I__2320 (
            .O(N__16236),
            .I(data_in_2_5));
    LocalMux I__2319 (
            .O(N__16233),
            .I(data_in_2_5));
    InMux I__2318 (
            .O(N__16224),
            .I(N__16221));
    LocalMux I__2317 (
            .O(N__16221),
            .I(N__16216));
    InMux I__2316 (
            .O(N__16220),
            .I(N__16211));
    InMux I__2315 (
            .O(N__16219),
            .I(N__16211));
    Span4Mux_h I__2314 (
            .O(N__16216),
            .I(N__16208));
    LocalMux I__2313 (
            .O(N__16211),
            .I(data_in_5_6));
    Odrv4 I__2312 (
            .O(N__16208),
            .I(data_in_5_6));
    InMux I__2311 (
            .O(N__16203),
            .I(N__16200));
    LocalMux I__2310 (
            .O(N__16200),
            .I(N__16197));
    Span4Mux_v I__2309 (
            .O(N__16197),
            .I(N__16192));
    InMux I__2308 (
            .O(N__16196),
            .I(N__16189));
    InMux I__2307 (
            .O(N__16195),
            .I(N__16186));
    Odrv4 I__2306 (
            .O(N__16192),
            .I(data_in_4_6));
    LocalMux I__2305 (
            .O(N__16189),
            .I(data_in_4_6));
    LocalMux I__2304 (
            .O(N__16186),
            .I(data_in_4_6));
    InMux I__2303 (
            .O(N__16179),
            .I(N__16174));
    InMux I__2302 (
            .O(N__16178),
            .I(N__16166));
    InMux I__2301 (
            .O(N__16177),
            .I(N__16166));
    LocalMux I__2300 (
            .O(N__16174),
            .I(N__16163));
    InMux I__2299 (
            .O(N__16173),
            .I(N__16158));
    InMux I__2298 (
            .O(N__16172),
            .I(N__16158));
    InMux I__2297 (
            .O(N__16171),
            .I(N__16155));
    LocalMux I__2296 (
            .O(N__16166),
            .I(r_Bit_Index_0_adj_1743));
    Odrv4 I__2295 (
            .O(N__16163),
            .I(r_Bit_Index_0_adj_1743));
    LocalMux I__2294 (
            .O(N__16158),
            .I(r_Bit_Index_0_adj_1743));
    LocalMux I__2293 (
            .O(N__16155),
            .I(r_Bit_Index_0_adj_1743));
    InMux I__2292 (
            .O(N__16146),
            .I(N__16139));
    InMux I__2291 (
            .O(N__16145),
            .I(N__16139));
    InMux I__2290 (
            .O(N__16144),
            .I(N__16136));
    LocalMux I__2289 (
            .O(N__16139),
            .I(N__16133));
    LocalMux I__2288 (
            .O(N__16136),
            .I(n9075));
    Odrv4 I__2287 (
            .O(N__16133),
            .I(n9075));
    InMux I__2286 (
            .O(N__16128),
            .I(N__16122));
    InMux I__2285 (
            .O(N__16127),
            .I(N__16122));
    LocalMux I__2284 (
            .O(N__16122),
            .I(N__16118));
    InMux I__2283 (
            .O(N__16121),
            .I(N__16115));
    Odrv4 I__2282 (
            .O(N__16118),
            .I(n5346));
    LocalMux I__2281 (
            .O(N__16115),
            .I(n5346));
    InMux I__2280 (
            .O(N__16110),
            .I(N__16104));
    CascadeMux I__2279 (
            .O(N__16109),
            .I(N__16099));
    CascadeMux I__2278 (
            .O(N__16108),
            .I(N__16096));
    CascadeMux I__2277 (
            .O(N__16107),
            .I(N__16092));
    LocalMux I__2276 (
            .O(N__16104),
            .I(N__16089));
    InMux I__2275 (
            .O(N__16103),
            .I(N__16082));
    InMux I__2274 (
            .O(N__16102),
            .I(N__16082));
    InMux I__2273 (
            .O(N__16099),
            .I(N__16082));
    InMux I__2272 (
            .O(N__16096),
            .I(N__16075));
    InMux I__2271 (
            .O(N__16095),
            .I(N__16075));
    InMux I__2270 (
            .O(N__16092),
            .I(N__16075));
    Odrv4 I__2269 (
            .O(N__16089),
            .I(r_Bit_Index_1_adj_1742));
    LocalMux I__2268 (
            .O(N__16082),
            .I(r_Bit_Index_1_adj_1742));
    LocalMux I__2267 (
            .O(N__16075),
            .I(r_Bit_Index_1_adj_1742));
    InMux I__2266 (
            .O(N__16068),
            .I(N__16065));
    LocalMux I__2265 (
            .O(N__16065),
            .I(N__16062));
    Span4Mux_v I__2264 (
            .O(N__16062),
            .I(N__16058));
    InMux I__2263 (
            .O(N__16061),
            .I(N__16055));
    Odrv4 I__2262 (
            .O(N__16058),
            .I(data_in_15_1));
    LocalMux I__2261 (
            .O(N__16055),
            .I(data_in_15_1));
    InMux I__2260 (
            .O(N__16050),
            .I(N__16046));
    InMux I__2259 (
            .O(N__16049),
            .I(N__16043));
    LocalMux I__2258 (
            .O(N__16046),
            .I(N__16040));
    LocalMux I__2257 (
            .O(N__16043),
            .I(N__16037));
    Span4Mux_v I__2256 (
            .O(N__16040),
            .I(N__16033));
    Span4Mux_h I__2255 (
            .O(N__16037),
            .I(N__16030));
    InMux I__2254 (
            .O(N__16036),
            .I(N__16027));
    Span4Mux_v I__2253 (
            .O(N__16033),
            .I(N__16024));
    Odrv4 I__2252 (
            .O(N__16030),
            .I(data_in_5_4));
    LocalMux I__2251 (
            .O(N__16027),
            .I(data_in_5_4));
    Odrv4 I__2250 (
            .O(N__16024),
            .I(data_in_5_4));
    InMux I__2249 (
            .O(N__16017),
            .I(N__16013));
    InMux I__2248 (
            .O(N__16016),
            .I(N__16010));
    LocalMux I__2247 (
            .O(N__16013),
            .I(data_in_17_1));
    LocalMux I__2246 (
            .O(N__16010),
            .I(data_in_17_1));
    InMux I__2245 (
            .O(N__16005),
            .I(N__16001));
    InMux I__2244 (
            .O(N__16004),
            .I(N__15998));
    LocalMux I__2243 (
            .O(N__16001),
            .I(data_in_16_1));
    LocalMux I__2242 (
            .O(N__15998),
            .I(data_in_16_1));
    InMux I__2241 (
            .O(N__15993),
            .I(N__15989));
    InMux I__2240 (
            .O(N__15992),
            .I(N__15986));
    LocalMux I__2239 (
            .O(N__15989),
            .I(data_in_14_7));
    LocalMux I__2238 (
            .O(N__15986),
            .I(data_in_14_7));
    InMux I__2237 (
            .O(N__15981),
            .I(N__15975));
    InMux I__2236 (
            .O(N__15980),
            .I(N__15975));
    LocalMux I__2235 (
            .O(N__15975),
            .I(data_in_15_7));
    InMux I__2234 (
            .O(N__15972),
            .I(N__15966));
    InMux I__2233 (
            .O(N__15971),
            .I(N__15966));
    LocalMux I__2232 (
            .O(N__15966),
            .I(data_in_16_7));
    InMux I__2231 (
            .O(N__15963),
            .I(N__15960));
    LocalMux I__2230 (
            .O(N__15960),
            .I(\c0.n24_adj_1615 ));
    InMux I__2229 (
            .O(N__15957),
            .I(N__15954));
    LocalMux I__2228 (
            .O(N__15954),
            .I(\c0.n34 ));
    InMux I__2227 (
            .O(N__15951),
            .I(N__15947));
    CascadeMux I__2226 (
            .O(N__15950),
            .I(N__15944));
    LocalMux I__2225 (
            .O(N__15947),
            .I(N__15934));
    InMux I__2224 (
            .O(N__15944),
            .I(N__15925));
    InMux I__2223 (
            .O(N__15943),
            .I(N__15925));
    InMux I__2222 (
            .O(N__15942),
            .I(N__15925));
    InMux I__2221 (
            .O(N__15941),
            .I(N__15925));
    InMux I__2220 (
            .O(N__15940),
            .I(N__15922));
    InMux I__2219 (
            .O(N__15939),
            .I(N__15915));
    InMux I__2218 (
            .O(N__15938),
            .I(N__15915));
    InMux I__2217 (
            .O(N__15937),
            .I(N__15915));
    Odrv12 I__2216 (
            .O(N__15934),
            .I(r_SM_Main_1_adj_1739));
    LocalMux I__2215 (
            .O(N__15925),
            .I(r_SM_Main_1_adj_1739));
    LocalMux I__2214 (
            .O(N__15922),
            .I(r_SM_Main_1_adj_1739));
    LocalMux I__2213 (
            .O(N__15915),
            .I(r_SM_Main_1_adj_1739));
    InMux I__2212 (
            .O(N__15906),
            .I(N__15903));
    LocalMux I__2211 (
            .O(N__15903),
            .I(n8747));
    InMux I__2210 (
            .O(N__15900),
            .I(N__15897));
    LocalMux I__2209 (
            .O(N__15897),
            .I(\c0.tx2.r_Tx_Data_7 ));
    CascadeMux I__2208 (
            .O(N__15894),
            .I(\c0.tx2.n9716_cascade_ ));
    InMux I__2207 (
            .O(N__15891),
            .I(N__15888));
    LocalMux I__2206 (
            .O(N__15888),
            .I(\c0.tx2.n9719 ));
    CascadeMux I__2205 (
            .O(N__15885),
            .I(n4691_cascade_));
    CascadeMux I__2204 (
            .O(N__15882),
            .I(\c0.n4574_cascade_ ));
    InMux I__2203 (
            .O(N__15879),
            .I(N__15873));
    InMux I__2202 (
            .O(N__15878),
            .I(N__15873));
    LocalMux I__2201 (
            .O(N__15873),
            .I(N__15866));
    InMux I__2200 (
            .O(N__15872),
            .I(N__15861));
    InMux I__2199 (
            .O(N__15871),
            .I(N__15861));
    InMux I__2198 (
            .O(N__15870),
            .I(N__15858));
    InMux I__2197 (
            .O(N__15869),
            .I(N__15855));
    Odrv4 I__2196 (
            .O(N__15866),
            .I(data_in_field_81));
    LocalMux I__2195 (
            .O(N__15861),
            .I(data_in_field_81));
    LocalMux I__2194 (
            .O(N__15858),
            .I(data_in_field_81));
    LocalMux I__2193 (
            .O(N__15855),
            .I(data_in_field_81));
    InMux I__2192 (
            .O(N__15846),
            .I(N__15842));
    InMux I__2191 (
            .O(N__15845),
            .I(N__15838));
    LocalMux I__2190 (
            .O(N__15842),
            .I(N__15834));
    InMux I__2189 (
            .O(N__15841),
            .I(N__15831));
    LocalMux I__2188 (
            .O(N__15838),
            .I(N__15828));
    InMux I__2187 (
            .O(N__15837),
            .I(N__15823));
    Span12Mux_h I__2186 (
            .O(N__15834),
            .I(N__15818));
    LocalMux I__2185 (
            .O(N__15831),
            .I(N__15818));
    Span4Mux_s2_h I__2184 (
            .O(N__15828),
            .I(N__15815));
    InMux I__2183 (
            .O(N__15827),
            .I(N__15810));
    InMux I__2182 (
            .O(N__15826),
            .I(N__15810));
    LocalMux I__2181 (
            .O(N__15823),
            .I(data_in_field_47));
    Odrv12 I__2180 (
            .O(N__15818),
            .I(data_in_field_47));
    Odrv4 I__2179 (
            .O(N__15815),
            .I(data_in_field_47));
    LocalMux I__2178 (
            .O(N__15810),
            .I(data_in_field_47));
    InMux I__2177 (
            .O(N__15801),
            .I(N__15798));
    LocalMux I__2176 (
            .O(N__15798),
            .I(\c0.n4333 ));
    CascadeMux I__2175 (
            .O(N__15795),
            .I(\c0.n4333_cascade_ ));
    InMux I__2174 (
            .O(N__15792),
            .I(N__15789));
    LocalMux I__2173 (
            .O(N__15789),
            .I(n3_adj_1749));
    IoInMux I__2172 (
            .O(N__15786),
            .I(N__15783));
    LocalMux I__2171 (
            .O(N__15783),
            .I(N__15779));
    InMux I__2170 (
            .O(N__15782),
            .I(N__15776));
    IoSpan4Mux I__2169 (
            .O(N__15779),
            .I(N__15773));
    LocalMux I__2168 (
            .O(N__15776),
            .I(N__15770));
    Span4Mux_s3_h I__2167 (
            .O(N__15773),
            .I(N__15764));
    Span4Mux_s3_h I__2166 (
            .O(N__15770),
            .I(N__15764));
    InMux I__2165 (
            .O(N__15769),
            .I(N__15761));
    Odrv4 I__2164 (
            .O(N__15764),
            .I(tx2_o));
    LocalMux I__2163 (
            .O(N__15761),
            .I(tx2_o));
    CascadeMux I__2162 (
            .O(N__15756),
            .I(\c0.n8788_cascade_ ));
    InMux I__2161 (
            .O(N__15753),
            .I(N__15750));
    LocalMux I__2160 (
            .O(N__15750),
            .I(\c0.n14_adj_1648 ));
    CascadeMux I__2159 (
            .O(N__15747),
            .I(N__15744));
    InMux I__2158 (
            .O(N__15744),
            .I(N__15741));
    LocalMux I__2157 (
            .O(N__15741),
            .I(N__15737));
    InMux I__2156 (
            .O(N__15740),
            .I(N__15734));
    Odrv4 I__2155 (
            .O(N__15737),
            .I(\c0.n8936 ));
    LocalMux I__2154 (
            .O(N__15734),
            .I(\c0.n8936 ));
    CascadeMux I__2153 (
            .O(N__15729),
            .I(\c0.n24_adj_1600_cascade_ ));
    InMux I__2152 (
            .O(N__15726),
            .I(N__15723));
    LocalMux I__2151 (
            .O(N__15723),
            .I(\c0.n18_adj_1603 ));
    InMux I__2150 (
            .O(N__15720),
            .I(N__15716));
    InMux I__2149 (
            .O(N__15719),
            .I(N__15713));
    LocalMux I__2148 (
            .O(N__15716),
            .I(N__15710));
    LocalMux I__2147 (
            .O(N__15713),
            .I(N__15707));
    Odrv4 I__2146 (
            .O(N__15710),
            .I(\c0.n4107 ));
    Odrv12 I__2145 (
            .O(N__15707),
            .I(\c0.n4107 ));
    CascadeMux I__2144 (
            .O(N__15702),
            .I(\c0.tx2_transmit_N_1334_cascade_ ));
    InMux I__2143 (
            .O(N__15699),
            .I(N__15696));
    LocalMux I__2142 (
            .O(N__15696),
            .I(N__15693));
    Odrv4 I__2141 (
            .O(N__15693),
            .I(\c0.n8980 ));
    CascadeMux I__2140 (
            .O(N__15690),
            .I(\c0.n22_adj_1601_cascade_ ));
    InMux I__2139 (
            .O(N__15687),
            .I(N__15684));
    LocalMux I__2138 (
            .O(N__15684),
            .I(\c0.n26 ));
    InMux I__2137 (
            .O(N__15681),
            .I(N__15678));
    LocalMux I__2136 (
            .O(N__15678),
            .I(N__15675));
    Span4Mux_h I__2135 (
            .O(N__15675),
            .I(N__15672));
    Odrv4 I__2134 (
            .O(N__15672),
            .I(\c0.n16 ));
    InMux I__2133 (
            .O(N__15669),
            .I(N__15663));
    InMux I__2132 (
            .O(N__15668),
            .I(N__15660));
    InMux I__2131 (
            .O(N__15667),
            .I(N__15655));
    InMux I__2130 (
            .O(N__15666),
            .I(N__15655));
    LocalMux I__2129 (
            .O(N__15663),
            .I(N__15652));
    LocalMux I__2128 (
            .O(N__15660),
            .I(data_in_field_115));
    LocalMux I__2127 (
            .O(N__15655),
            .I(data_in_field_115));
    Odrv12 I__2126 (
            .O(N__15652),
            .I(data_in_field_115));
    InMux I__2125 (
            .O(N__15645),
            .I(N__15642));
    LocalMux I__2124 (
            .O(N__15642),
            .I(\c0.n4452 ));
    CascadeMux I__2123 (
            .O(N__15639),
            .I(\c0.n4253_cascade_ ));
    InMux I__2122 (
            .O(N__15636),
            .I(N__15632));
    InMux I__2121 (
            .O(N__15635),
            .I(N__15629));
    LocalMux I__2120 (
            .O(N__15632),
            .I(N__15626));
    LocalMux I__2119 (
            .O(N__15629),
            .I(N__15621));
    Span4Mux_s2_v I__2118 (
            .O(N__15626),
            .I(N__15618));
    InMux I__2117 (
            .O(N__15625),
            .I(N__15613));
    InMux I__2116 (
            .O(N__15624),
            .I(N__15613));
    Odrv4 I__2115 (
            .O(N__15621),
            .I(data_in_field_71));
    Odrv4 I__2114 (
            .O(N__15618),
            .I(data_in_field_71));
    LocalMux I__2113 (
            .O(N__15613),
            .I(data_in_field_71));
    InMux I__2112 (
            .O(N__15606),
            .I(N__15599));
    InMux I__2111 (
            .O(N__15605),
            .I(N__15599));
    InMux I__2110 (
            .O(N__15604),
            .I(N__15596));
    LocalMux I__2109 (
            .O(N__15599),
            .I(N__15591));
    LocalMux I__2108 (
            .O(N__15596),
            .I(N__15588));
    InMux I__2107 (
            .O(N__15595),
            .I(N__15585));
    InMux I__2106 (
            .O(N__15594),
            .I(N__15582));
    Span4Mux_v I__2105 (
            .O(N__15591),
            .I(N__15575));
    Span4Mux_v I__2104 (
            .O(N__15588),
            .I(N__15575));
    LocalMux I__2103 (
            .O(N__15585),
            .I(N__15575));
    LocalMux I__2102 (
            .O(N__15582),
            .I(data_in_field_147));
    Odrv4 I__2101 (
            .O(N__15575),
            .I(data_in_field_147));
    CascadeMux I__2100 (
            .O(N__15570),
            .I(N__15565));
    CascadeMux I__2099 (
            .O(N__15569),
            .I(N__15562));
    CascadeMux I__2098 (
            .O(N__15568),
            .I(N__15559));
    InMux I__2097 (
            .O(N__15565),
            .I(N__15555));
    InMux I__2096 (
            .O(N__15562),
            .I(N__15550));
    InMux I__2095 (
            .O(N__15559),
            .I(N__15550));
    InMux I__2094 (
            .O(N__15558),
            .I(N__15547));
    LocalMux I__2093 (
            .O(N__15555),
            .I(N__15542));
    LocalMux I__2092 (
            .O(N__15550),
            .I(N__15542));
    LocalMux I__2091 (
            .O(N__15547),
            .I(data_in_field_127));
    Odrv4 I__2090 (
            .O(N__15542),
            .I(data_in_field_127));
    InMux I__2089 (
            .O(N__15537),
            .I(N__15534));
    LocalMux I__2088 (
            .O(N__15534),
            .I(\c0.n9650 ));
    InMux I__2087 (
            .O(N__15531),
            .I(N__15528));
    LocalMux I__2086 (
            .O(N__15528),
            .I(N__15525));
    Span4Mux_s3_h I__2085 (
            .O(N__15525),
            .I(N__15522));
    Odrv4 I__2084 (
            .O(N__15522),
            .I(\c0.n16_adj_1598 ));
    InMux I__2083 (
            .O(N__15519),
            .I(N__15515));
    InMux I__2082 (
            .O(N__15518),
            .I(N__15512));
    LocalMux I__2081 (
            .O(N__15515),
            .I(N__15509));
    LocalMux I__2080 (
            .O(N__15512),
            .I(N__15506));
    Span4Mux_s2_h I__2079 (
            .O(N__15509),
            .I(N__15501));
    Span4Mux_h I__2078 (
            .O(N__15506),
            .I(N__15501));
    Odrv4 I__2077 (
            .O(N__15501),
            .I(\c0.n9016 ));
    CascadeMux I__2076 (
            .O(N__15498),
            .I(\c0.n6_adj_1645_cascade_ ));
    InMux I__2075 (
            .O(N__15495),
            .I(N__15492));
    LocalMux I__2074 (
            .O(N__15492),
            .I(N__15488));
    InMux I__2073 (
            .O(N__15491),
            .I(N__15485));
    Span4Mux_v I__2072 (
            .O(N__15488),
            .I(N__15480));
    LocalMux I__2071 (
            .O(N__15485),
            .I(N__15480));
    Odrv4 I__2070 (
            .O(N__15480),
            .I(\c0.n4154 ));
    CascadeMux I__2069 (
            .O(N__15477),
            .I(\c0.n10_adj_1640_cascade_ ));
    InMux I__2068 (
            .O(N__15474),
            .I(N__15471));
    LocalMux I__2067 (
            .O(N__15471),
            .I(N__15468));
    Span4Mux_v I__2066 (
            .O(N__15468),
            .I(N__15465));
    Odrv4 I__2065 (
            .O(N__15465),
            .I(\c0.n4434 ));
    CascadeMux I__2064 (
            .O(N__15462),
            .I(\c0.n8933_cascade_ ));
    InMux I__2063 (
            .O(N__15459),
            .I(N__15455));
    InMux I__2062 (
            .O(N__15458),
            .I(N__15452));
    LocalMux I__2061 (
            .O(N__15455),
            .I(N__15449));
    LocalMux I__2060 (
            .O(N__15452),
            .I(\c0.n8822 ));
    Odrv4 I__2059 (
            .O(N__15449),
            .I(\c0.n8822 ));
    CascadeMux I__2058 (
            .O(N__15444),
            .I(\c0.n8314_cascade_ ));
    CascadeMux I__2057 (
            .O(N__15441),
            .I(N__15437));
    InMux I__2056 (
            .O(N__15440),
            .I(N__15431));
    InMux I__2055 (
            .O(N__15437),
            .I(N__15431));
    CascadeMux I__2054 (
            .O(N__15436),
            .I(N__15428));
    LocalMux I__2053 (
            .O(N__15431),
            .I(N__15425));
    InMux I__2052 (
            .O(N__15428),
            .I(N__15422));
    Span4Mux_h I__2051 (
            .O(N__15425),
            .I(N__15416));
    LocalMux I__2050 (
            .O(N__15422),
            .I(N__15416));
    InMux I__2049 (
            .O(N__15421),
            .I(N__15411));
    Span4Mux_v I__2048 (
            .O(N__15416),
            .I(N__15408));
    InMux I__2047 (
            .O(N__15415),
            .I(N__15403));
    InMux I__2046 (
            .O(N__15414),
            .I(N__15403));
    LocalMux I__2045 (
            .O(N__15411),
            .I(N__15400));
    Odrv4 I__2044 (
            .O(N__15408),
            .I(data_in_field_145));
    LocalMux I__2043 (
            .O(N__15403),
            .I(data_in_field_145));
    Odrv4 I__2042 (
            .O(N__15400),
            .I(data_in_field_145));
    InMux I__2041 (
            .O(N__15393),
            .I(N__15390));
    LocalMux I__2040 (
            .O(N__15390),
            .I(N__15387));
    Span4Mux_s3_h I__2039 (
            .O(N__15387),
            .I(N__15383));
    InMux I__2038 (
            .O(N__15386),
            .I(N__15380));
    Odrv4 I__2037 (
            .O(N__15383),
            .I(\c0.n4556 ));
    LocalMux I__2036 (
            .O(N__15380),
            .I(\c0.n4556 ));
    InMux I__2035 (
            .O(N__15375),
            .I(N__15372));
    LocalMux I__2034 (
            .O(N__15372),
            .I(N__15368));
    InMux I__2033 (
            .O(N__15371),
            .I(N__15365));
    Odrv4 I__2032 (
            .O(N__15368),
            .I(\c0.n8861 ));
    LocalMux I__2031 (
            .O(N__15365),
            .I(\c0.n8861 ));
    InMux I__2030 (
            .O(N__15360),
            .I(N__15357));
    LocalMux I__2029 (
            .O(N__15357),
            .I(\c0.n6 ));
    CascadeMux I__2028 (
            .O(N__15354),
            .I(\c0.n4452_cascade_ ));
    CascadeMux I__2027 (
            .O(N__15351),
            .I(N__15347));
    InMux I__2026 (
            .O(N__15350),
            .I(N__15344));
    InMux I__2025 (
            .O(N__15347),
            .I(N__15341));
    LocalMux I__2024 (
            .O(N__15344),
            .I(N__15338));
    LocalMux I__2023 (
            .O(N__15341),
            .I(N__15335));
    Span4Mux_v I__2022 (
            .O(N__15338),
            .I(N__15330));
    Span4Mux_v I__2021 (
            .O(N__15335),
            .I(N__15330));
    Odrv4 I__2020 (
            .O(N__15330),
            .I(\c0.n8906 ));
    InMux I__2019 (
            .O(N__15327),
            .I(N__15324));
    LocalMux I__2018 (
            .O(N__15324),
            .I(N__15321));
    Span4Mux_v I__2017 (
            .O(N__15321),
            .I(N__15318));
    Odrv4 I__2016 (
            .O(N__15318),
            .I(n1892));
    InMux I__2015 (
            .O(N__15315),
            .I(N__15312));
    LocalMux I__2014 (
            .O(N__15312),
            .I(N__15309));
    Span4Mux_h I__2013 (
            .O(N__15309),
            .I(N__15306));
    Span4Mux_s0_h I__2012 (
            .O(N__15306),
            .I(N__15303));
    Odrv4 I__2011 (
            .O(N__15303),
            .I(n1891));
    InMux I__2010 (
            .O(N__15300),
            .I(N__15297));
    LocalMux I__2009 (
            .O(N__15297),
            .I(\c0.n8831 ));
    InMux I__2008 (
            .O(N__15294),
            .I(N__15288));
    InMux I__2007 (
            .O(N__15293),
            .I(N__15285));
    InMux I__2006 (
            .O(N__15292),
            .I(N__15282));
    InMux I__2005 (
            .O(N__15291),
            .I(N__15279));
    LocalMux I__2004 (
            .O(N__15288),
            .I(\c0.data_in_field_9 ));
    LocalMux I__2003 (
            .O(N__15285),
            .I(\c0.data_in_field_9 ));
    LocalMux I__2002 (
            .O(N__15282),
            .I(\c0.data_in_field_9 ));
    LocalMux I__2001 (
            .O(N__15279),
            .I(\c0.data_in_field_9 ));
    CascadeMux I__2000 (
            .O(N__15270),
            .I(\c0.n8831_cascade_ ));
    InMux I__1999 (
            .O(N__15267),
            .I(N__15264));
    LocalMux I__1998 (
            .O(N__15264),
            .I(N__15258));
    InMux I__1997 (
            .O(N__15263),
            .I(N__15255));
    InMux I__1996 (
            .O(N__15262),
            .I(N__15252));
    InMux I__1995 (
            .O(N__15261),
            .I(N__15249));
    Span4Mux_h I__1994 (
            .O(N__15258),
            .I(N__15244));
    LocalMux I__1993 (
            .O(N__15255),
            .I(N__15244));
    LocalMux I__1992 (
            .O(N__15252),
            .I(N__15239));
    LocalMux I__1991 (
            .O(N__15249),
            .I(N__15239));
    Span4Mux_v I__1990 (
            .O(N__15244),
            .I(N__15236));
    Odrv4 I__1989 (
            .O(N__15239),
            .I(data_in_1_0));
    Odrv4 I__1988 (
            .O(N__15236),
            .I(data_in_1_0));
    InMux I__1987 (
            .O(N__15231),
            .I(N__15228));
    LocalMux I__1986 (
            .O(N__15228),
            .I(N__15225));
    Span4Mux_h I__1985 (
            .O(N__15225),
            .I(N__15222));
    Span4Mux_s1_h I__1984 (
            .O(N__15222),
            .I(N__15219));
    Odrv4 I__1983 (
            .O(N__15219),
            .I(n1888));
    InMux I__1982 (
            .O(N__15216),
            .I(N__15212));
    InMux I__1981 (
            .O(N__15215),
            .I(N__15208));
    LocalMux I__1980 (
            .O(N__15212),
            .I(N__15205));
    InMux I__1979 (
            .O(N__15211),
            .I(N__15202));
    LocalMux I__1978 (
            .O(N__15208),
            .I(N__15199));
    Odrv12 I__1977 (
            .O(N__15205),
            .I(data_in_5_3));
    LocalMux I__1976 (
            .O(N__15202),
            .I(data_in_5_3));
    Odrv4 I__1975 (
            .O(N__15199),
            .I(data_in_5_3));
    InMux I__1974 (
            .O(N__15192),
            .I(N__15189));
    LocalMux I__1973 (
            .O(N__15189),
            .I(N__15186));
    Span4Mux_v I__1972 (
            .O(N__15186),
            .I(N__15182));
    InMux I__1971 (
            .O(N__15185),
            .I(N__15179));
    Span4Mux_s2_h I__1970 (
            .O(N__15182),
            .I(N__15175));
    LocalMux I__1969 (
            .O(N__15179),
            .I(N__15172));
    InMux I__1968 (
            .O(N__15178),
            .I(N__15169));
    Odrv4 I__1967 (
            .O(N__15175),
            .I(data_in_4_3));
    Odrv4 I__1966 (
            .O(N__15172),
            .I(data_in_4_3));
    LocalMux I__1965 (
            .O(N__15169),
            .I(data_in_4_3));
    InMux I__1964 (
            .O(N__15162),
            .I(N__15157));
    InMux I__1963 (
            .O(N__15161),
            .I(N__15154));
    InMux I__1962 (
            .O(N__15160),
            .I(N__15151));
    LocalMux I__1961 (
            .O(N__15157),
            .I(\c0.n4131 ));
    LocalMux I__1960 (
            .O(N__15154),
            .I(\c0.n4131 ));
    LocalMux I__1959 (
            .O(N__15151),
            .I(\c0.n4131 ));
    CascadeMux I__1958 (
            .O(N__15144),
            .I(N__15141));
    InMux I__1957 (
            .O(N__15141),
            .I(N__15138));
    LocalMux I__1956 (
            .O(N__15138),
            .I(N__15133));
    InMux I__1955 (
            .O(N__15137),
            .I(N__15130));
    InMux I__1954 (
            .O(N__15136),
            .I(N__15127));
    Span4Mux_h I__1953 (
            .O(N__15133),
            .I(N__15124));
    LocalMux I__1952 (
            .O(N__15130),
            .I(\c0.n4224 ));
    LocalMux I__1951 (
            .O(N__15127),
            .I(\c0.n4224 ));
    Odrv4 I__1950 (
            .O(N__15124),
            .I(\c0.n4224 ));
    InMux I__1949 (
            .O(N__15117),
            .I(N__15114));
    LocalMux I__1948 (
            .O(N__15114),
            .I(N__15111));
    Odrv12 I__1947 (
            .O(N__15111),
            .I(\c0.n4127 ));
    CascadeMux I__1946 (
            .O(N__15108),
            .I(N__15105));
    InMux I__1945 (
            .O(N__15105),
            .I(N__15102));
    LocalMux I__1944 (
            .O(N__15102),
            .I(N__15097));
    InMux I__1943 (
            .O(N__15101),
            .I(N__15092));
    InMux I__1942 (
            .O(N__15100),
            .I(N__15092));
    Odrv4 I__1941 (
            .O(N__15097),
            .I(data_in_0_3));
    LocalMux I__1940 (
            .O(N__15092),
            .I(data_in_0_3));
    InMux I__1939 (
            .O(N__15087),
            .I(N__15081));
    InMux I__1938 (
            .O(N__15086),
            .I(N__15078));
    InMux I__1937 (
            .O(N__15085),
            .I(N__15075));
    InMux I__1936 (
            .O(N__15084),
            .I(N__15072));
    LocalMux I__1935 (
            .O(N__15081),
            .I(N__15069));
    LocalMux I__1934 (
            .O(N__15078),
            .I(N__15064));
    LocalMux I__1933 (
            .O(N__15075),
            .I(N__15064));
    LocalMux I__1932 (
            .O(N__15072),
            .I(N__15058));
    Span4Mux_v I__1931 (
            .O(N__15069),
            .I(N__15058));
    Span4Mux_s3_h I__1930 (
            .O(N__15064),
            .I(N__15055));
    InMux I__1929 (
            .O(N__15063),
            .I(N__15052));
    Odrv4 I__1928 (
            .O(N__15058),
            .I(\c0.data_in_field_3 ));
    Odrv4 I__1927 (
            .O(N__15055),
            .I(\c0.data_in_field_3 ));
    LocalMux I__1926 (
            .O(N__15052),
            .I(\c0.data_in_field_3 ));
    InMux I__1925 (
            .O(N__15045),
            .I(N__15042));
    LocalMux I__1924 (
            .O(N__15042),
            .I(N__15039));
    Odrv4 I__1923 (
            .O(N__15039),
            .I(\c0.n20_adj_1597 ));
    InMux I__1922 (
            .O(N__15036),
            .I(N__15033));
    LocalMux I__1921 (
            .O(N__15033),
            .I(N__15030));
    Odrv12 I__1920 (
            .O(N__15030),
            .I(\c0.n22_adj_1595 ));
    InMux I__1919 (
            .O(N__15027),
            .I(N__15023));
    InMux I__1918 (
            .O(N__15026),
            .I(N__15019));
    LocalMux I__1917 (
            .O(N__15023),
            .I(N__15015));
    InMux I__1916 (
            .O(N__15022),
            .I(N__15012));
    LocalMux I__1915 (
            .O(N__15019),
            .I(N__15009));
    InMux I__1914 (
            .O(N__15018),
            .I(N__15006));
    Odrv4 I__1913 (
            .O(N__15015),
            .I(data_in_2_6));
    LocalMux I__1912 (
            .O(N__15012),
            .I(data_in_2_6));
    Odrv12 I__1911 (
            .O(N__15009),
            .I(data_in_2_6));
    LocalMux I__1910 (
            .O(N__15006),
            .I(data_in_2_6));
    CascadeMux I__1909 (
            .O(N__14997),
            .I(n9069_cascade_));
    InMux I__1908 (
            .O(N__14994),
            .I(N__14990));
    InMux I__1907 (
            .O(N__14993),
            .I(N__14986));
    LocalMux I__1906 (
            .O(N__14990),
            .I(N__14982));
    InMux I__1905 (
            .O(N__14989),
            .I(N__14979));
    LocalMux I__1904 (
            .O(N__14986),
            .I(N__14976));
    InMux I__1903 (
            .O(N__14985),
            .I(N__14973));
    Span4Mux_s3_h I__1902 (
            .O(N__14982),
            .I(N__14970));
    LocalMux I__1901 (
            .O(N__14979),
            .I(N__14965));
    Span4Mux_s3_h I__1900 (
            .O(N__14976),
            .I(N__14965));
    LocalMux I__1899 (
            .O(N__14973),
            .I(data_in_3_3));
    Odrv4 I__1898 (
            .O(N__14970),
            .I(data_in_3_3));
    Odrv4 I__1897 (
            .O(N__14965),
            .I(data_in_3_3));
    InMux I__1896 (
            .O(N__14958),
            .I(N__14955));
    LocalMux I__1895 (
            .O(N__14955),
            .I(N__14952));
    Odrv4 I__1894 (
            .O(N__14952),
            .I(\c0.n8849 ));
    CascadeMux I__1893 (
            .O(N__14949),
            .I(n4_adj_1750_cascade_));
    InMux I__1892 (
            .O(N__14946),
            .I(N__14943));
    LocalMux I__1891 (
            .O(N__14943),
            .I(N__14938));
    InMux I__1890 (
            .O(N__14942),
            .I(N__14935));
    InMux I__1889 (
            .O(N__14941),
            .I(N__14931));
    Span4Mux_v I__1888 (
            .O(N__14938),
            .I(N__14928));
    LocalMux I__1887 (
            .O(N__14935),
            .I(N__14925));
    InMux I__1886 (
            .O(N__14934),
            .I(N__14922));
    LocalMux I__1885 (
            .O(N__14931),
            .I(\c0.data_in_field_2 ));
    Odrv4 I__1884 (
            .O(N__14928),
            .I(\c0.data_in_field_2 ));
    Odrv4 I__1883 (
            .O(N__14925),
            .I(\c0.data_in_field_2 ));
    LocalMux I__1882 (
            .O(N__14922),
            .I(\c0.data_in_field_2 ));
    InMux I__1881 (
            .O(N__14913),
            .I(N__14909));
    InMux I__1880 (
            .O(N__14912),
            .I(N__14906));
    LocalMux I__1879 (
            .O(N__14909),
            .I(N__14902));
    LocalMux I__1878 (
            .O(N__14906),
            .I(N__14899));
    InMux I__1877 (
            .O(N__14905),
            .I(N__14894));
    Span4Mux_s3_h I__1876 (
            .O(N__14902),
            .I(N__14889));
    Span4Mux_s3_h I__1875 (
            .O(N__14899),
            .I(N__14889));
    InMux I__1874 (
            .O(N__14898),
            .I(N__14886));
    InMux I__1873 (
            .O(N__14897),
            .I(N__14883));
    LocalMux I__1872 (
            .O(N__14894),
            .I(\c0.data_in_field_33 ));
    Odrv4 I__1871 (
            .O(N__14889),
            .I(\c0.data_in_field_33 ));
    LocalMux I__1870 (
            .O(N__14886),
            .I(\c0.data_in_field_33 ));
    LocalMux I__1869 (
            .O(N__14883),
            .I(\c0.data_in_field_33 ));
    CascadeMux I__1868 (
            .O(N__14874),
            .I(\c0.n6_adj_1632_cascade_ ));
    InMux I__1867 (
            .O(N__14871),
            .I(N__14868));
    LocalMux I__1866 (
            .O(N__14868),
            .I(\c0.n8804 ));
    InMux I__1865 (
            .O(N__14865),
            .I(N__14862));
    LocalMux I__1864 (
            .O(N__14862),
            .I(N__14858));
    InMux I__1863 (
            .O(N__14861),
            .I(N__14853));
    Span4Mux_v I__1862 (
            .O(N__14858),
            .I(N__14850));
    InMux I__1861 (
            .O(N__14857),
            .I(N__14847));
    InMux I__1860 (
            .O(N__14856),
            .I(N__14844));
    LocalMux I__1859 (
            .O(N__14853),
            .I(data_in_1_6));
    Odrv4 I__1858 (
            .O(N__14850),
            .I(data_in_1_6));
    LocalMux I__1857 (
            .O(N__14847),
            .I(data_in_1_6));
    LocalMux I__1856 (
            .O(N__14844),
            .I(data_in_1_6));
    CascadeMux I__1855 (
            .O(N__14835),
            .I(N__14832));
    InMux I__1854 (
            .O(N__14832),
            .I(N__14827));
    InMux I__1853 (
            .O(N__14831),
            .I(N__14824));
    CascadeMux I__1852 (
            .O(N__14830),
            .I(N__14821));
    LocalMux I__1851 (
            .O(N__14827),
            .I(N__14817));
    LocalMux I__1850 (
            .O(N__14824),
            .I(N__14814));
    InMux I__1849 (
            .O(N__14821),
            .I(N__14809));
    InMux I__1848 (
            .O(N__14820),
            .I(N__14809));
    Span4Mux_h I__1847 (
            .O(N__14817),
            .I(N__14806));
    Span4Mux_v I__1846 (
            .O(N__14814),
            .I(N__14803));
    LocalMux I__1845 (
            .O(N__14809),
            .I(data_in_3_7));
    Odrv4 I__1844 (
            .O(N__14806),
            .I(data_in_3_7));
    Odrv4 I__1843 (
            .O(N__14803),
            .I(data_in_3_7));
    InMux I__1842 (
            .O(N__14796),
            .I(N__14793));
    LocalMux I__1841 (
            .O(N__14793),
            .I(N__14789));
    InMux I__1840 (
            .O(N__14792),
            .I(N__14786));
    Odrv4 I__1839 (
            .O(N__14789),
            .I(data_in_13_0));
    LocalMux I__1838 (
            .O(N__14786),
            .I(data_in_13_0));
    InMux I__1837 (
            .O(N__14781),
            .I(N__14778));
    LocalMux I__1836 (
            .O(N__14778),
            .I(N__14773));
    InMux I__1835 (
            .O(N__14777),
            .I(N__14770));
    InMux I__1834 (
            .O(N__14776),
            .I(N__14767));
    Odrv4 I__1833 (
            .O(N__14773),
            .I(data_in_4_0));
    LocalMux I__1832 (
            .O(N__14770),
            .I(data_in_4_0));
    LocalMux I__1831 (
            .O(N__14767),
            .I(data_in_4_0));
    InMux I__1830 (
            .O(N__14760),
            .I(N__14757));
    LocalMux I__1829 (
            .O(N__14757),
            .I(\c0.n13_adj_1671 ));
    InMux I__1828 (
            .O(N__14754),
            .I(N__14751));
    LocalMux I__1827 (
            .O(N__14751),
            .I(\c0.n13_adj_1672 ));
    InMux I__1826 (
            .O(N__14748),
            .I(N__14744));
    InMux I__1825 (
            .O(N__14747),
            .I(N__14741));
    LocalMux I__1824 (
            .O(N__14744),
            .I(N__14737));
    LocalMux I__1823 (
            .O(N__14741),
            .I(N__14734));
    CascadeMux I__1822 (
            .O(N__14740),
            .I(N__14730));
    Span4Mux_v I__1821 (
            .O(N__14737),
            .I(N__14727));
    Span4Mux_s3_h I__1820 (
            .O(N__14734),
            .I(N__14724));
    InMux I__1819 (
            .O(N__14733),
            .I(N__14721));
    InMux I__1818 (
            .O(N__14730),
            .I(N__14718));
    Odrv4 I__1817 (
            .O(N__14727),
            .I(data_in_1_2));
    Odrv4 I__1816 (
            .O(N__14724),
            .I(data_in_1_2));
    LocalMux I__1815 (
            .O(N__14721),
            .I(data_in_1_2));
    LocalMux I__1814 (
            .O(N__14718),
            .I(data_in_1_2));
    InMux I__1813 (
            .O(N__14709),
            .I(N__14706));
    LocalMux I__1812 (
            .O(N__14706),
            .I(N__14701));
    InMux I__1811 (
            .O(N__14705),
            .I(N__14696));
    InMux I__1810 (
            .O(N__14704),
            .I(N__14696));
    Odrv4 I__1809 (
            .O(N__14701),
            .I(data_in_6_3));
    LocalMux I__1808 (
            .O(N__14696),
            .I(data_in_6_3));
    CascadeMux I__1807 (
            .O(N__14691),
            .I(N__14688));
    InMux I__1806 (
            .O(N__14688),
            .I(N__14685));
    LocalMux I__1805 (
            .O(N__14685),
            .I(N__14682));
    Span4Mux_v I__1804 (
            .O(N__14682),
            .I(N__14676));
    InMux I__1803 (
            .O(N__14681),
            .I(N__14669));
    InMux I__1802 (
            .O(N__14680),
            .I(N__14669));
    InMux I__1801 (
            .O(N__14679),
            .I(N__14669));
    Odrv4 I__1800 (
            .O(N__14676),
            .I(data_in_1_3));
    LocalMux I__1799 (
            .O(N__14669),
            .I(data_in_1_3));
    InMux I__1798 (
            .O(N__14664),
            .I(N__14661));
    LocalMux I__1797 (
            .O(N__14661),
            .I(N__14657));
    CascadeMux I__1796 (
            .O(N__14660),
            .I(N__14654));
    Span4Mux_s3_h I__1795 (
            .O(N__14657),
            .I(N__14649));
    InMux I__1794 (
            .O(N__14654),
            .I(N__14642));
    InMux I__1793 (
            .O(N__14653),
            .I(N__14642));
    InMux I__1792 (
            .O(N__14652),
            .I(N__14642));
    Odrv4 I__1791 (
            .O(N__14649),
            .I(data_in_2_3));
    LocalMux I__1790 (
            .O(N__14642),
            .I(data_in_2_3));
    CascadeMux I__1789 (
            .O(N__14637),
            .I(N__14634));
    InMux I__1788 (
            .O(N__14634),
            .I(N__14631));
    LocalMux I__1787 (
            .O(N__14631),
            .I(N__14628));
    Odrv4 I__1786 (
            .O(N__14628),
            .I(\c0.n4495 ));
    InMux I__1785 (
            .O(N__14625),
            .I(N__14621));
    InMux I__1784 (
            .O(N__14624),
            .I(N__14618));
    LocalMux I__1783 (
            .O(N__14621),
            .I(data_in_15_6));
    LocalMux I__1782 (
            .O(N__14618),
            .I(data_in_15_6));
    InMux I__1781 (
            .O(N__14613),
            .I(N__14609));
    InMux I__1780 (
            .O(N__14612),
            .I(N__14606));
    LocalMux I__1779 (
            .O(N__14609),
            .I(data_in_14_6));
    LocalMux I__1778 (
            .O(N__14606),
            .I(data_in_14_6));
    InMux I__1777 (
            .O(N__14601),
            .I(N__14597));
    InMux I__1776 (
            .O(N__14600),
            .I(N__14594));
    LocalMux I__1775 (
            .O(N__14597),
            .I(data_in_20_4));
    LocalMux I__1774 (
            .O(N__14594),
            .I(data_in_20_4));
    InMux I__1773 (
            .O(N__14589),
            .I(N__14585));
    InMux I__1772 (
            .O(N__14588),
            .I(N__14580));
    LocalMux I__1771 (
            .O(N__14585),
            .I(N__14577));
    CascadeMux I__1770 (
            .O(N__14584),
            .I(N__14574));
    InMux I__1769 (
            .O(N__14583),
            .I(N__14571));
    LocalMux I__1768 (
            .O(N__14580),
            .I(N__14566));
    Span4Mux_v I__1767 (
            .O(N__14577),
            .I(N__14566));
    InMux I__1766 (
            .O(N__14574),
            .I(N__14563));
    LocalMux I__1765 (
            .O(N__14571),
            .I(data_in_3_0));
    Odrv4 I__1764 (
            .O(N__14566),
            .I(data_in_3_0));
    LocalMux I__1763 (
            .O(N__14563),
            .I(data_in_3_0));
    InMux I__1762 (
            .O(N__14556),
            .I(N__14552));
    InMux I__1761 (
            .O(N__14555),
            .I(N__14548));
    LocalMux I__1760 (
            .O(N__14552),
            .I(N__14545));
    InMux I__1759 (
            .O(N__14551),
            .I(N__14542));
    LocalMux I__1758 (
            .O(N__14548),
            .I(data_in_0_5));
    Odrv4 I__1757 (
            .O(N__14545),
            .I(data_in_0_5));
    LocalMux I__1756 (
            .O(N__14542),
            .I(data_in_0_5));
    CascadeMux I__1755 (
            .O(N__14535),
            .I(\c0.n28_adj_1668_cascade_ ));
    InMux I__1754 (
            .O(N__14532),
            .I(N__14529));
    LocalMux I__1753 (
            .O(N__14529),
            .I(\c0.n30_adj_1674 ));
    InMux I__1752 (
            .O(N__14526),
            .I(N__14523));
    LocalMux I__1751 (
            .O(N__14523),
            .I(\c0.n22_adj_1667 ));
    InMux I__1750 (
            .O(N__14520),
            .I(N__14517));
    LocalMux I__1749 (
            .O(N__14517),
            .I(N__14514));
    Span4Mux_s3_h I__1748 (
            .O(N__14514),
            .I(N__14509));
    InMux I__1747 (
            .O(N__14513),
            .I(N__14504));
    InMux I__1746 (
            .O(N__14512),
            .I(N__14504));
    Odrv4 I__1745 (
            .O(N__14509),
            .I(data_in_0_0));
    LocalMux I__1744 (
            .O(N__14504),
            .I(data_in_0_0));
    InMux I__1743 (
            .O(N__14499),
            .I(N__14496));
    LocalMux I__1742 (
            .O(N__14496),
            .I(N__14493));
    Span4Mux_s3_h I__1741 (
            .O(N__14493),
            .I(N__14489));
    InMux I__1740 (
            .O(N__14492),
            .I(N__14486));
    Odrv4 I__1739 (
            .O(N__14489),
            .I(data_in_13_7));
    LocalMux I__1738 (
            .O(N__14486),
            .I(data_in_13_7));
    InMux I__1737 (
            .O(N__14481),
            .I(N__14475));
    InMux I__1736 (
            .O(N__14480),
            .I(N__14475));
    LocalMux I__1735 (
            .O(N__14475),
            .I(data_in_16_6));
    InMux I__1734 (
            .O(N__14472),
            .I(N__14468));
    InMux I__1733 (
            .O(N__14471),
            .I(N__14465));
    LocalMux I__1732 (
            .O(N__14468),
            .I(data_in_9_6));
    LocalMux I__1731 (
            .O(N__14465),
            .I(data_in_9_6));
    InMux I__1730 (
            .O(N__14460),
            .I(N__14454));
    InMux I__1729 (
            .O(N__14459),
            .I(N__14454));
    LocalMux I__1728 (
            .O(N__14454),
            .I(data_in_10_6));
    InMux I__1727 (
            .O(N__14451),
            .I(N__14445));
    InMux I__1726 (
            .O(N__14450),
            .I(N__14445));
    LocalMux I__1725 (
            .O(N__14445),
            .I(data_in_11_6));
    InMux I__1724 (
            .O(N__14442),
            .I(N__14438));
    InMux I__1723 (
            .O(N__14441),
            .I(N__14435));
    LocalMux I__1722 (
            .O(N__14438),
            .I(data_in_13_6));
    LocalMux I__1721 (
            .O(N__14435),
            .I(data_in_13_6));
    InMux I__1720 (
            .O(N__14430),
            .I(N__14424));
    InMux I__1719 (
            .O(N__14429),
            .I(N__14424));
    LocalMux I__1718 (
            .O(N__14424),
            .I(data_in_12_6));
    CascadeMux I__1717 (
            .O(N__14421),
            .I(\c0.n9752_cascade_ ));
    InMux I__1716 (
            .O(N__14418),
            .I(N__14414));
    InMux I__1715 (
            .O(N__14417),
            .I(N__14410));
    LocalMux I__1714 (
            .O(N__14414),
            .I(N__14406));
    InMux I__1713 (
            .O(N__14413),
            .I(N__14403));
    LocalMux I__1712 (
            .O(N__14410),
            .I(N__14400));
    InMux I__1711 (
            .O(N__14409),
            .I(N__14396));
    Span12Mux_s3_v I__1710 (
            .O(N__14406),
            .I(N__14393));
    LocalMux I__1709 (
            .O(N__14403),
            .I(N__14388));
    Span4Mux_v I__1708 (
            .O(N__14400),
            .I(N__14388));
    InMux I__1707 (
            .O(N__14399),
            .I(N__14385));
    LocalMux I__1706 (
            .O(N__14396),
            .I(\c0.data_in_field_39 ));
    Odrv12 I__1705 (
            .O(N__14393),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__1704 (
            .O(N__14388),
            .I(\c0.data_in_field_39 ));
    LocalMux I__1703 (
            .O(N__14385),
            .I(\c0.data_in_field_39 ));
    InMux I__1702 (
            .O(N__14376),
            .I(N__14373));
    LocalMux I__1701 (
            .O(N__14373),
            .I(\c0.n9120 ));
    InMux I__1700 (
            .O(N__14370),
            .I(N__14367));
    LocalMux I__1699 (
            .O(N__14367),
            .I(N__14364));
    Span4Mux_s2_v I__1698 (
            .O(N__14364),
            .I(N__14361));
    Odrv4 I__1697 (
            .O(N__14361),
            .I(\c0.tx2.r_Tx_Data_3 ));
    InMux I__1696 (
            .O(N__14358),
            .I(N__14355));
    LocalMux I__1695 (
            .O(N__14355),
            .I(N__14352));
    Span4Mux_h I__1694 (
            .O(N__14352),
            .I(N__14349));
    Odrv4 I__1693 (
            .O(N__14349),
            .I(\c0.tx2.r_Tx_Data_1 ));
    CascadeMux I__1692 (
            .O(N__14346),
            .I(\c0.tx2.n9692_cascade_ ));
    CascadeMux I__1691 (
            .O(N__14343),
            .I(\c0.tx2.n9695_cascade_ ));
    CascadeMux I__1690 (
            .O(N__14340),
            .I(\c0.tx2.o_Tx_Serial_N_1511_cascade_ ));
    CascadeMux I__1689 (
            .O(N__14337),
            .I(n2207_cascade_));
    InMux I__1688 (
            .O(N__14334),
            .I(N__14327));
    InMux I__1687 (
            .O(N__14333),
            .I(N__14327));
    InMux I__1686 (
            .O(N__14332),
            .I(N__14324));
    LocalMux I__1685 (
            .O(N__14327),
            .I(r_Bit_Index_2_adj_1741));
    LocalMux I__1684 (
            .O(N__14324),
            .I(r_Bit_Index_2_adj_1741));
    CascadeMux I__1683 (
            .O(N__14319),
            .I(N__14311));
    InMux I__1682 (
            .O(N__14318),
            .I(N__14308));
    CascadeMux I__1681 (
            .O(N__14317),
            .I(N__14305));
    CascadeMux I__1680 (
            .O(N__14316),
            .I(N__14301));
    InMux I__1679 (
            .O(N__14315),
            .I(N__14292));
    InMux I__1678 (
            .O(N__14314),
            .I(N__14292));
    InMux I__1677 (
            .O(N__14311),
            .I(N__14292));
    LocalMux I__1676 (
            .O(N__14308),
            .I(N__14289));
    InMux I__1675 (
            .O(N__14305),
            .I(N__14284));
    InMux I__1674 (
            .O(N__14304),
            .I(N__14284));
    InMux I__1673 (
            .O(N__14301),
            .I(N__14277));
    InMux I__1672 (
            .O(N__14300),
            .I(N__14277));
    InMux I__1671 (
            .O(N__14299),
            .I(N__14277));
    LocalMux I__1670 (
            .O(N__14292),
            .I(r_SM_Main_0_adj_1740));
    Odrv4 I__1669 (
            .O(N__14289),
            .I(r_SM_Main_0_adj_1740));
    LocalMux I__1668 (
            .O(N__14284),
            .I(r_SM_Main_0_adj_1740));
    LocalMux I__1667 (
            .O(N__14277),
            .I(r_SM_Main_0_adj_1740));
    InMux I__1666 (
            .O(N__14268),
            .I(N__14261));
    InMux I__1665 (
            .O(N__14267),
            .I(N__14252));
    InMux I__1664 (
            .O(N__14266),
            .I(N__14252));
    InMux I__1663 (
            .O(N__14265),
            .I(N__14252));
    InMux I__1662 (
            .O(N__14264),
            .I(N__14252));
    LocalMux I__1661 (
            .O(N__14261),
            .I(r_SM_Main_2_N_1480_1_adj_1744));
    LocalMux I__1660 (
            .O(N__14252),
            .I(r_SM_Main_2_N_1480_1_adj_1744));
    InMux I__1659 (
            .O(N__14247),
            .I(N__14241));
    InMux I__1658 (
            .O(N__14246),
            .I(N__14238));
    InMux I__1657 (
            .O(N__14245),
            .I(N__14233));
    InMux I__1656 (
            .O(N__14244),
            .I(N__14233));
    LocalMux I__1655 (
            .O(N__14241),
            .I(N__14230));
    LocalMux I__1654 (
            .O(N__14238),
            .I(data_in_field_83));
    LocalMux I__1653 (
            .O(N__14233),
            .I(data_in_field_83));
    Odrv4 I__1652 (
            .O(N__14230),
            .I(data_in_field_83));
    InMux I__1651 (
            .O(N__14223),
            .I(N__14220));
    LocalMux I__1650 (
            .O(N__14220),
            .I(N__14217));
    Odrv4 I__1649 (
            .O(N__14217),
            .I(\c0.n9126 ));
    CascadeMux I__1648 (
            .O(N__14214),
            .I(\c0.n9123_cascade_ ));
    InMux I__1647 (
            .O(N__14211),
            .I(N__14208));
    LocalMux I__1646 (
            .O(N__14208),
            .I(N__14205));
    Span4Mux_s2_v I__1645 (
            .O(N__14205),
            .I(N__14202));
    Odrv4 I__1644 (
            .O(N__14202),
            .I(\c0.n9240 ));
    CascadeMux I__1643 (
            .O(N__14199),
            .I(\c0.n9644_cascade_ ));
    CascadeMux I__1642 (
            .O(N__14196),
            .I(\c0.n9647_cascade_ ));
    InMux I__1641 (
            .O(N__14193),
            .I(N__14190));
    LocalMux I__1640 (
            .O(N__14190),
            .I(\c0.n9656 ));
    InMux I__1639 (
            .O(N__14187),
            .I(N__14184));
    LocalMux I__1638 (
            .O(N__14184),
            .I(n6164));
    InMux I__1637 (
            .O(N__14181),
            .I(N__14178));
    LocalMux I__1636 (
            .O(N__14178),
            .I(N__14173));
    InMux I__1635 (
            .O(N__14177),
            .I(N__14168));
    InMux I__1634 (
            .O(N__14176),
            .I(N__14168));
    Odrv12 I__1633 (
            .O(N__14173),
            .I(data_in_field_105));
    LocalMux I__1632 (
            .O(N__14168),
            .I(data_in_field_105));
    CascadeMux I__1631 (
            .O(N__14163),
            .I(\c0.n8890_cascade_ ));
    InMux I__1630 (
            .O(N__14160),
            .I(N__14157));
    LocalMux I__1629 (
            .O(N__14157),
            .I(N__14154));
    Span4Mux_h I__1628 (
            .O(N__14154),
            .I(N__14151));
    Span4Mux_v I__1627 (
            .O(N__14151),
            .I(N__14148));
    Odrv4 I__1626 (
            .O(N__14148),
            .I(\c0.n14_adj_1638 ));
    InMux I__1625 (
            .O(N__14145),
            .I(N__14142));
    LocalMux I__1624 (
            .O(N__14142),
            .I(N__14139));
    Odrv4 I__1623 (
            .O(N__14139),
            .I(\c0.n4285 ));
    InMux I__1622 (
            .O(N__14136),
            .I(N__14132));
    InMux I__1621 (
            .O(N__14135),
            .I(N__14129));
    LocalMux I__1620 (
            .O(N__14132),
            .I(N__14126));
    LocalMux I__1619 (
            .O(N__14129),
            .I(N__14123));
    Odrv12 I__1618 (
            .O(N__14126),
            .I(\c0.n9007 ));
    Odrv4 I__1617 (
            .O(N__14123),
            .I(\c0.n9007 ));
    CascadeMux I__1616 (
            .O(N__14118),
            .I(\c0.n18_adj_1589_cascade_ ));
    CascadeMux I__1615 (
            .O(N__14115),
            .I(\c0.n20_adj_1590_cascade_ ));
    InMux I__1614 (
            .O(N__14112),
            .I(N__14109));
    LocalMux I__1613 (
            .O(N__14109),
            .I(N__14105));
    InMux I__1612 (
            .O(N__14108),
            .I(N__14102));
    Sp12to4 I__1611 (
            .O(N__14105),
            .I(N__14097));
    LocalMux I__1610 (
            .O(N__14102),
            .I(N__14097));
    Odrv12 I__1609 (
            .O(N__14097),
            .I(\c0.n29 ));
    InMux I__1608 (
            .O(N__14094),
            .I(N__14091));
    LocalMux I__1607 (
            .O(N__14091),
            .I(N__14088));
    Odrv4 I__1606 (
            .O(N__14088),
            .I(\c0.n4114 ));
    InMux I__1605 (
            .O(N__14085),
            .I(N__14082));
    LocalMux I__1604 (
            .O(N__14082),
            .I(\c0.n4448 ));
    InMux I__1603 (
            .O(N__14079),
            .I(N__14076));
    LocalMux I__1602 (
            .O(N__14076),
            .I(\c0.n4445 ));
    CascadeMux I__1601 (
            .O(N__14073),
            .I(N__14070));
    InMux I__1600 (
            .O(N__14070),
            .I(N__14067));
    LocalMux I__1599 (
            .O(N__14067),
            .I(N__14063));
    InMux I__1598 (
            .O(N__14066),
            .I(N__14060));
    Odrv12 I__1597 (
            .O(N__14063),
            .I(\c0.n8896 ));
    LocalMux I__1596 (
            .O(N__14060),
            .I(\c0.n8896 ));
    CascadeMux I__1595 (
            .O(N__14055),
            .I(\c0.n10_adj_1647_cascade_ ));
    CascadeMux I__1594 (
            .O(N__14052),
            .I(N__14049));
    InMux I__1593 (
            .O(N__14049),
            .I(N__14046));
    LocalMux I__1592 (
            .O(N__14046),
            .I(N__14043));
    Odrv4 I__1591 (
            .O(N__14043),
            .I(\c0.data_in_frame_19_1 ));
    CascadeMux I__1590 (
            .O(N__14040),
            .I(\c0.n9704_cascade_ ));
    InMux I__1589 (
            .O(N__14037),
            .I(N__14034));
    LocalMux I__1588 (
            .O(N__14034),
            .I(N__14031));
    Span4Mux_v I__1587 (
            .O(N__14031),
            .I(N__14028));
    Span4Mux_h I__1586 (
            .O(N__14028),
            .I(N__14025));
    Odrv4 I__1585 (
            .O(N__14025),
            .I(\c0.data_in_frame_20_1 ));
    CascadeMux I__1584 (
            .O(N__14022),
            .I(\c0.n9707_cascade_ ));
    InMux I__1583 (
            .O(N__14019),
            .I(N__14016));
    LocalMux I__1582 (
            .O(N__14016),
            .I(N__14013));
    Span4Mux_s3_h I__1581 (
            .O(N__14013),
            .I(N__14010));
    Odrv4 I__1580 (
            .O(N__14010),
            .I(\c0.n22_adj_1682 ));
    CascadeMux I__1579 (
            .O(N__14007),
            .I(\c0.n9722_cascade_ ));
    InMux I__1578 (
            .O(N__14004),
            .I(N__14000));
    InMux I__1577 (
            .O(N__14003),
            .I(N__13995));
    LocalMux I__1576 (
            .O(N__14000),
            .I(N__13992));
    InMux I__1575 (
            .O(N__13999),
            .I(N__13987));
    InMux I__1574 (
            .O(N__13998),
            .I(N__13987));
    LocalMux I__1573 (
            .O(N__13995),
            .I(\c0.data_in_field_7 ));
    Odrv4 I__1572 (
            .O(N__13992),
            .I(\c0.data_in_field_7 ));
    LocalMux I__1571 (
            .O(N__13987),
            .I(\c0.data_in_field_7 ));
    CascadeMux I__1570 (
            .O(N__13980),
            .I(N__13976));
    InMux I__1569 (
            .O(N__13979),
            .I(N__13973));
    InMux I__1568 (
            .O(N__13976),
            .I(N__13968));
    LocalMux I__1567 (
            .O(N__13973),
            .I(N__13965));
    InMux I__1566 (
            .O(N__13972),
            .I(N__13960));
    InMux I__1565 (
            .O(N__13971),
            .I(N__13960));
    LocalMux I__1564 (
            .O(N__13968),
            .I(\c0.data_in_field_23 ));
    Odrv4 I__1563 (
            .O(N__13965),
            .I(\c0.data_in_field_23 ));
    LocalMux I__1562 (
            .O(N__13960),
            .I(\c0.data_in_field_23 ));
    InMux I__1561 (
            .O(N__13953),
            .I(N__13949));
    InMux I__1560 (
            .O(N__13952),
            .I(N__13946));
    LocalMux I__1559 (
            .O(N__13949),
            .I(N__13943));
    LocalMux I__1558 (
            .O(N__13946),
            .I(\c0.n4514 ));
    Odrv12 I__1557 (
            .O(N__13943),
            .I(\c0.n4514 ));
    CascadeMux I__1556 (
            .O(N__13938),
            .I(N__13935));
    InMux I__1555 (
            .O(N__13935),
            .I(N__13928));
    InMux I__1554 (
            .O(N__13934),
            .I(N__13921));
    InMux I__1553 (
            .O(N__13933),
            .I(N__13921));
    InMux I__1552 (
            .O(N__13932),
            .I(N__13921));
    InMux I__1551 (
            .O(N__13931),
            .I(N__13918));
    LocalMux I__1550 (
            .O(N__13928),
            .I(N__13913));
    LocalMux I__1549 (
            .O(N__13921),
            .I(N__13913));
    LocalMux I__1548 (
            .O(N__13918),
            .I(\c0.data_in_field_4 ));
    Odrv4 I__1547 (
            .O(N__13913),
            .I(\c0.data_in_field_4 ));
    InMux I__1546 (
            .O(N__13908),
            .I(N__13905));
    LocalMux I__1545 (
            .O(N__13905),
            .I(N__13900));
    CascadeMux I__1544 (
            .O(N__13904),
            .I(N__13897));
    InMux I__1543 (
            .O(N__13903),
            .I(N__13894));
    Span4Mux_v I__1542 (
            .O(N__13900),
            .I(N__13891));
    InMux I__1541 (
            .O(N__13897),
            .I(N__13888));
    LocalMux I__1540 (
            .O(N__13894),
            .I(data_in_0_7));
    Odrv4 I__1539 (
            .O(N__13891),
            .I(data_in_0_7));
    LocalMux I__1538 (
            .O(N__13888),
            .I(data_in_0_7));
    InMux I__1537 (
            .O(N__13881),
            .I(N__13878));
    LocalMux I__1536 (
            .O(N__13878),
            .I(N__13873));
    InMux I__1535 (
            .O(N__13877),
            .I(N__13868));
    InMux I__1534 (
            .O(N__13876),
            .I(N__13868));
    Odrv4 I__1533 (
            .O(N__13873),
            .I(\c0.n8776 ));
    LocalMux I__1532 (
            .O(N__13868),
            .I(\c0.n8776 ));
    CascadeMux I__1531 (
            .O(N__13863),
            .I(\c0.n4131_cascade_ ));
    CascadeMux I__1530 (
            .O(N__13860),
            .I(\c0.n8927_cascade_ ));
    InMux I__1529 (
            .O(N__13857),
            .I(N__13854));
    LocalMux I__1528 (
            .O(N__13854),
            .I(N__13851));
    Span4Mux_v I__1527 (
            .O(N__13851),
            .I(N__13848));
    Odrv4 I__1526 (
            .O(N__13848),
            .I(n1896));
    InMux I__1525 (
            .O(N__13845),
            .I(N__13842));
    LocalMux I__1524 (
            .O(N__13842),
            .I(N__13839));
    Span4Mux_h I__1523 (
            .O(N__13839),
            .I(N__13833));
    InMux I__1522 (
            .O(N__13838),
            .I(N__13828));
    InMux I__1521 (
            .O(N__13837),
            .I(N__13828));
    InMux I__1520 (
            .O(N__13836),
            .I(N__13825));
    Odrv4 I__1519 (
            .O(N__13833),
            .I(data_in_2_7));
    LocalMux I__1518 (
            .O(N__13828),
            .I(data_in_2_7));
    LocalMux I__1517 (
            .O(N__13825),
            .I(data_in_2_7));
    InMux I__1516 (
            .O(N__13818),
            .I(N__13814));
    InMux I__1515 (
            .O(N__13817),
            .I(N__13810));
    LocalMux I__1514 (
            .O(N__13814),
            .I(N__13807));
    InMux I__1513 (
            .O(N__13813),
            .I(N__13804));
    LocalMux I__1512 (
            .O(N__13810),
            .I(data_in_0_6));
    Odrv4 I__1511 (
            .O(N__13807),
            .I(data_in_0_6));
    LocalMux I__1510 (
            .O(N__13804),
            .I(data_in_0_6));
    InMux I__1509 (
            .O(N__13797),
            .I(N__13793));
    InMux I__1508 (
            .O(N__13796),
            .I(N__13787));
    LocalMux I__1507 (
            .O(N__13793),
            .I(N__13784));
    InMux I__1506 (
            .O(N__13792),
            .I(N__13777));
    InMux I__1505 (
            .O(N__13791),
            .I(N__13777));
    InMux I__1504 (
            .O(N__13790),
            .I(N__13777));
    LocalMux I__1503 (
            .O(N__13787),
            .I(\c0.data_in_field_19 ));
    Odrv4 I__1502 (
            .O(N__13784),
            .I(\c0.data_in_field_19 ));
    LocalMux I__1501 (
            .O(N__13777),
            .I(\c0.data_in_field_19 ));
    InMux I__1500 (
            .O(N__13770),
            .I(N__13767));
    LocalMux I__1499 (
            .O(N__13767),
            .I(\c0.n14 ));
    CascadeMux I__1498 (
            .O(N__13764),
            .I(\c0.n10_adj_1631_cascade_ ));
    InMux I__1497 (
            .O(N__13761),
            .I(N__13757));
    CascadeMux I__1496 (
            .O(N__13760),
            .I(N__13754));
    LocalMux I__1495 (
            .O(N__13757),
            .I(N__13749));
    InMux I__1494 (
            .O(N__13754),
            .I(N__13742));
    InMux I__1493 (
            .O(N__13753),
            .I(N__13742));
    InMux I__1492 (
            .O(N__13752),
            .I(N__13742));
    Odrv4 I__1491 (
            .O(N__13749),
            .I(data_in_1_1));
    LocalMux I__1490 (
            .O(N__13742),
            .I(data_in_1_1));
    InMux I__1489 (
            .O(N__13737),
            .I(N__13734));
    LocalMux I__1488 (
            .O(N__13734),
            .I(N__13730));
    InMux I__1487 (
            .O(N__13733),
            .I(N__13727));
    Span4Mux_v I__1486 (
            .O(N__13730),
            .I(N__13724));
    LocalMux I__1485 (
            .O(N__13727),
            .I(N__13721));
    Span4Mux_v I__1484 (
            .O(N__13724),
            .I(N__13717));
    Sp12to4 I__1483 (
            .O(N__13721),
            .I(N__13714));
    InMux I__1482 (
            .O(N__13720),
            .I(N__13711));
    Odrv4 I__1481 (
            .O(N__13717),
            .I(data_in_4_7));
    Odrv12 I__1480 (
            .O(N__13714),
            .I(data_in_4_7));
    LocalMux I__1479 (
            .O(N__13711),
            .I(data_in_4_7));
    CascadeMux I__1478 (
            .O(N__13704),
            .I(N__13701));
    InMux I__1477 (
            .O(N__13701),
            .I(N__13698));
    LocalMux I__1476 (
            .O(N__13698),
            .I(N__13695));
    Span4Mux_s2_h I__1475 (
            .O(N__13695),
            .I(N__13692));
    Odrv4 I__1474 (
            .O(N__13692),
            .I(\c0.n47 ));
    InMux I__1473 (
            .O(N__13689),
            .I(N__13686));
    LocalMux I__1472 (
            .O(N__13686),
            .I(N__13681));
    InMux I__1471 (
            .O(N__13685),
            .I(N__13678));
    InMux I__1470 (
            .O(N__13684),
            .I(N__13675));
    Odrv4 I__1469 (
            .O(N__13681),
            .I(data_in_0_2));
    LocalMux I__1468 (
            .O(N__13678),
            .I(data_in_0_2));
    LocalMux I__1467 (
            .O(N__13675),
            .I(data_in_0_2));
    InMux I__1466 (
            .O(N__13668),
            .I(N__13665));
    LocalMux I__1465 (
            .O(N__13665),
            .I(\c0.n4381 ));
    CascadeMux I__1464 (
            .O(N__13662),
            .I(\c0.n4381_cascade_ ));
    InMux I__1463 (
            .O(N__13659),
            .I(N__13648));
    InMux I__1462 (
            .O(N__13658),
            .I(N__13648));
    InMux I__1461 (
            .O(N__13657),
            .I(N__13648));
    InMux I__1460 (
            .O(N__13656),
            .I(N__13643));
    InMux I__1459 (
            .O(N__13655),
            .I(N__13643));
    LocalMux I__1458 (
            .O(N__13648),
            .I(\c0.data_in_field_20 ));
    LocalMux I__1457 (
            .O(N__13643),
            .I(\c0.data_in_field_20 ));
    CascadeMux I__1456 (
            .O(N__13638),
            .I(N__13635));
    InMux I__1455 (
            .O(N__13635),
            .I(N__13632));
    LocalMux I__1454 (
            .O(N__13632),
            .I(N__13629));
    Span4Mux_v I__1453 (
            .O(N__13629),
            .I(N__13624));
    InMux I__1452 (
            .O(N__13628),
            .I(N__13619));
    InMux I__1451 (
            .O(N__13627),
            .I(N__13619));
    IoSpan4Mux I__1450 (
            .O(N__13624),
            .I(N__13616));
    LocalMux I__1449 (
            .O(N__13619),
            .I(data_in_4_1));
    Odrv4 I__1448 (
            .O(N__13616),
            .I(data_in_4_1));
    InMux I__1447 (
            .O(N__13611),
            .I(N__13607));
    InMux I__1446 (
            .O(N__13610),
            .I(N__13601));
    LocalMux I__1445 (
            .O(N__13607),
            .I(N__13598));
    InMux I__1444 (
            .O(N__13606),
            .I(N__13591));
    InMux I__1443 (
            .O(N__13605),
            .I(N__13591));
    InMux I__1442 (
            .O(N__13604),
            .I(N__13591));
    LocalMux I__1441 (
            .O(N__13601),
            .I(\c0.data_in_field_35 ));
    Odrv4 I__1440 (
            .O(N__13598),
            .I(\c0.data_in_field_35 ));
    LocalMux I__1439 (
            .O(N__13591),
            .I(\c0.data_in_field_35 ));
    CascadeMux I__1438 (
            .O(N__13584),
            .I(\c0.n4154_cascade_ ));
    CascadeMux I__1437 (
            .O(N__13581),
            .I(N__13578));
    InMux I__1436 (
            .O(N__13578),
            .I(N__13575));
    LocalMux I__1435 (
            .O(N__13575),
            .I(\c0.n9578 ));
    InMux I__1434 (
            .O(N__13572),
            .I(N__13569));
    LocalMux I__1433 (
            .O(N__13569),
            .I(\c0.n8794 ));
    InMux I__1432 (
            .O(N__13566),
            .I(N__13562));
    CascadeMux I__1431 (
            .O(N__13565),
            .I(N__13558));
    LocalMux I__1430 (
            .O(N__13562),
            .I(N__13554));
    InMux I__1429 (
            .O(N__13561),
            .I(N__13549));
    InMux I__1428 (
            .O(N__13558),
            .I(N__13549));
    InMux I__1427 (
            .O(N__13557),
            .I(N__13546));
    Span4Mux_h I__1426 (
            .O(N__13554),
            .I(N__13543));
    LocalMux I__1425 (
            .O(N__13549),
            .I(N__13540));
    LocalMux I__1424 (
            .O(N__13546),
            .I(data_in_3_1));
    Odrv4 I__1423 (
            .O(N__13543),
            .I(data_in_3_1));
    Odrv4 I__1422 (
            .O(N__13540),
            .I(data_in_3_1));
    InMux I__1421 (
            .O(N__13533),
            .I(N__13529));
    InMux I__1420 (
            .O(N__13532),
            .I(N__13526));
    LocalMux I__1419 (
            .O(N__13529),
            .I(data_in_9_0));
    LocalMux I__1418 (
            .O(N__13526),
            .I(data_in_9_0));
    InMux I__1417 (
            .O(N__13521),
            .I(N__13517));
    InMux I__1416 (
            .O(N__13520),
            .I(N__13514));
    LocalMux I__1415 (
            .O(N__13517),
            .I(data_in_8_0));
    LocalMux I__1414 (
            .O(N__13514),
            .I(data_in_8_0));
    InMux I__1413 (
            .O(N__13509),
            .I(N__13503));
    InMux I__1412 (
            .O(N__13508),
            .I(N__13503));
    LocalMux I__1411 (
            .O(N__13503),
            .I(data_in_7_0));
    CascadeMux I__1410 (
            .O(N__13500),
            .I(N__13497));
    InMux I__1409 (
            .O(N__13497),
            .I(N__13493));
    CascadeMux I__1408 (
            .O(N__13496),
            .I(N__13488));
    LocalMux I__1407 (
            .O(N__13493),
            .I(N__13485));
    InMux I__1406 (
            .O(N__13492),
            .I(N__13482));
    InMux I__1405 (
            .O(N__13491),
            .I(N__13477));
    InMux I__1404 (
            .O(N__13488),
            .I(N__13477));
    Odrv4 I__1403 (
            .O(N__13485),
            .I(data_in_1_5));
    LocalMux I__1402 (
            .O(N__13482),
            .I(data_in_1_5));
    LocalMux I__1401 (
            .O(N__13477),
            .I(data_in_1_5));
    InMux I__1400 (
            .O(N__13470),
            .I(N__13467));
    LocalMux I__1399 (
            .O(N__13467),
            .I(N__13463));
    InMux I__1398 (
            .O(N__13466),
            .I(N__13460));
    Odrv4 I__1397 (
            .O(N__13463),
            .I(data_in_12_0));
    LocalMux I__1396 (
            .O(N__13460),
            .I(data_in_12_0));
    InMux I__1395 (
            .O(N__13455),
            .I(N__13452));
    LocalMux I__1394 (
            .O(N__13452),
            .I(N__13449));
    Span4Mux_v I__1393 (
            .O(N__13449),
            .I(N__13446));
    Odrv4 I__1392 (
            .O(N__13446),
            .I(\c0.n14_adj_1670 ));
    CascadeMux I__1391 (
            .O(N__13443),
            .I(N__13440));
    InMux I__1390 (
            .O(N__13440),
            .I(N__13437));
    LocalMux I__1389 (
            .O(N__13437),
            .I(\c0.n14_adj_1669 ));
    InMux I__1388 (
            .O(N__13434),
            .I(N__13431));
    LocalMux I__1387 (
            .O(N__13431),
            .I(N__13428));
    Span4Mux_v I__1386 (
            .O(N__13428),
            .I(N__13425));
    Odrv4 I__1385 (
            .O(N__13425),
            .I(\c0.n26_adj_1673 ));
    InMux I__1384 (
            .O(N__13422),
            .I(N__13419));
    LocalMux I__1383 (
            .O(N__13419),
            .I(\c0.n25_adj_1675 ));
    CascadeMux I__1382 (
            .O(N__13416),
            .I(\c0.n9033_cascade_ ));
    CascadeMux I__1381 (
            .O(N__13413),
            .I(n3220_cascade_));
    InMux I__1380 (
            .O(N__13410),
            .I(N__13406));
    InMux I__1379 (
            .O(N__13409),
            .I(N__13403));
    LocalMux I__1378 (
            .O(N__13406),
            .I(data_in_9_7));
    LocalMux I__1377 (
            .O(N__13403),
            .I(data_in_9_7));
    InMux I__1376 (
            .O(N__13398),
            .I(N__13394));
    InMux I__1375 (
            .O(N__13397),
            .I(N__13391));
    LocalMux I__1374 (
            .O(N__13394),
            .I(data_in_8_7));
    LocalMux I__1373 (
            .O(N__13391),
            .I(data_in_8_7));
    InMux I__1372 (
            .O(N__13386),
            .I(N__13383));
    LocalMux I__1371 (
            .O(N__13383),
            .I(N__13380));
    Span4Mux_v I__1370 (
            .O(N__13380),
            .I(N__13377));
    Odrv4 I__1369 (
            .O(N__13377),
            .I(n1900));
    InMux I__1368 (
            .O(N__13374),
            .I(N__13368));
    InMux I__1367 (
            .O(N__13373),
            .I(N__13368));
    LocalMux I__1366 (
            .O(N__13368),
            .I(data_in_7_3));
    InMux I__1365 (
            .O(N__13365),
            .I(N__13359));
    InMux I__1364 (
            .O(N__13364),
            .I(N__13359));
    LocalMux I__1363 (
            .O(N__13359),
            .I(data_in_8_3));
    InMux I__1362 (
            .O(N__13356),
            .I(N__13352));
    InMux I__1361 (
            .O(N__13355),
            .I(N__13349));
    LocalMux I__1360 (
            .O(N__13352),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1359 (
            .O(N__13349),
            .I(\c0.tx2.r_Clock_Count_5 ));
    CascadeMux I__1358 (
            .O(N__13344),
            .I(\c0.tx2.n5_cascade_ ));
    InMux I__1357 (
            .O(N__13341),
            .I(N__13337));
    InMux I__1356 (
            .O(N__13340),
            .I(N__13334));
    LocalMux I__1355 (
            .O(N__13337),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1354 (
            .O(N__13334),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__1353 (
            .O(N__13329),
            .I(N__13326));
    LocalMux I__1352 (
            .O(N__13326),
            .I(\c0.tx2.n4081 ));
    CascadeMux I__1351 (
            .O(N__13323),
            .I(\c0.tx2.n4081_cascade_ ));
    InMux I__1350 (
            .O(N__13320),
            .I(N__13317));
    LocalMux I__1349 (
            .O(N__13317),
            .I(\c0.tx2.n7 ));
    CascadeMux I__1348 (
            .O(N__13314),
            .I(\c0.tx2.n8196_cascade_ ));
    SRMux I__1347 (
            .O(N__13311),
            .I(N__13308));
    LocalMux I__1346 (
            .O(N__13308),
            .I(N__13304));
    SRMux I__1345 (
            .O(N__13307),
            .I(N__13301));
    Span4Mux_s1_h I__1344 (
            .O(N__13304),
            .I(N__13298));
    LocalMux I__1343 (
            .O(N__13301),
            .I(N__13295));
    Odrv4 I__1342 (
            .O(N__13298),
            .I(\c0.tx2.n5146 ));
    Odrv12 I__1341 (
            .O(N__13295),
            .I(\c0.tx2.n5146 ));
    CascadeMux I__1340 (
            .O(N__13290),
            .I(n9075_cascade_));
    InMux I__1339 (
            .O(N__13287),
            .I(N__13280));
    InMux I__1338 (
            .O(N__13286),
            .I(N__13277));
    InMux I__1337 (
            .O(N__13285),
            .I(N__13270));
    InMux I__1336 (
            .O(N__13284),
            .I(N__13270));
    InMux I__1335 (
            .O(N__13283),
            .I(N__13270));
    LocalMux I__1334 (
            .O(N__13280),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1333 (
            .O(N__13277),
            .I(\c0.tx2.r_Clock_Count_8 ));
    LocalMux I__1332 (
            .O(N__13270),
            .I(\c0.tx2.r_Clock_Count_8 ));
    InMux I__1331 (
            .O(N__13263),
            .I(N__13253));
    InMux I__1330 (
            .O(N__13262),
            .I(N__13253));
    InMux I__1329 (
            .O(N__13261),
            .I(N__13253));
    InMux I__1328 (
            .O(N__13260),
            .I(N__13250));
    LocalMux I__1327 (
            .O(N__13253),
            .I(\c0.tx2.n7399 ));
    LocalMux I__1326 (
            .O(N__13250),
            .I(\c0.tx2.n7399 ));
    InMux I__1325 (
            .O(N__13245),
            .I(N__13242));
    LocalMux I__1324 (
            .O(N__13242),
            .I(\c0.tx2.n7236 ));
    CascadeMux I__1323 (
            .O(N__13239),
            .I(\c0.tx2.n7236_cascade_ ));
    InMux I__1322 (
            .O(N__13236),
            .I(N__13233));
    LocalMux I__1321 (
            .O(N__13233),
            .I(N__13230));
    Span4Mux_v I__1320 (
            .O(N__13230),
            .I(N__13227));
    Odrv4 I__1319 (
            .O(N__13227),
            .I(\c0.n4577 ));
    InMux I__1318 (
            .O(N__13224),
            .I(N__13221));
    LocalMux I__1317 (
            .O(N__13221),
            .I(\c0.n4282 ));
    CascadeMux I__1316 (
            .O(N__13218),
            .I(\c0.n4476_cascade_ ));
    InMux I__1315 (
            .O(N__13215),
            .I(N__13212));
    LocalMux I__1314 (
            .O(N__13212),
            .I(N__13209));
    Span4Mux_v I__1313 (
            .O(N__13209),
            .I(N__13206));
    Odrv4 I__1312 (
            .O(N__13206),
            .I(\c0.n19_adj_1623 ));
    InMux I__1311 (
            .O(N__13203),
            .I(N__13199));
    InMux I__1310 (
            .O(N__13202),
            .I(N__13196));
    LocalMux I__1309 (
            .O(N__13199),
            .I(N__13190));
    LocalMux I__1308 (
            .O(N__13196),
            .I(N__13190));
    InMux I__1307 (
            .O(N__13195),
            .I(N__13187));
    Span4Mux_v I__1306 (
            .O(N__13190),
            .I(N__13184));
    LocalMux I__1305 (
            .O(N__13187),
            .I(data_in_5_7));
    Odrv4 I__1304 (
            .O(N__13184),
            .I(data_in_5_7));
    IoInMux I__1303 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__1302 (
            .O(N__13176),
            .I(N__13173));
    Span4Mux_s1_h I__1301 (
            .O(N__13173),
            .I(N__13170));
    Odrv4 I__1300 (
            .O(N__13170),
            .I(tx2_enable));
    InMux I__1299 (
            .O(N__13167),
            .I(N__13163));
    InMux I__1298 (
            .O(N__13166),
            .I(N__13160));
    LocalMux I__1297 (
            .O(N__13163),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1296 (
            .O(N__13160),
            .I(\c0.tx2.r_Clock_Count_2 ));
    InMux I__1295 (
            .O(N__13155),
            .I(N__13151));
    InMux I__1294 (
            .O(N__13154),
            .I(N__13148));
    LocalMux I__1293 (
            .O(N__13151),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1292 (
            .O(N__13148),
            .I(\c0.tx2.r_Clock_Count_6 ));
    CascadeMux I__1291 (
            .O(N__13143),
            .I(N__13139));
    InMux I__1290 (
            .O(N__13142),
            .I(N__13136));
    InMux I__1289 (
            .O(N__13139),
            .I(N__13133));
    LocalMux I__1288 (
            .O(N__13136),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1287 (
            .O(N__13133),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__1286 (
            .O(N__13128),
            .I(N__13124));
    InMux I__1285 (
            .O(N__13127),
            .I(N__13121));
    LocalMux I__1284 (
            .O(N__13124),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1283 (
            .O(N__13121),
            .I(\c0.tx2.r_Clock_Count_3 ));
    InMux I__1282 (
            .O(N__13116),
            .I(N__13112));
    InMux I__1281 (
            .O(N__13115),
            .I(N__13109));
    LocalMux I__1280 (
            .O(N__13112),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1279 (
            .O(N__13109),
            .I(\c0.tx2.r_Clock_Count_4 ));
    CascadeMux I__1278 (
            .O(N__13104),
            .I(\c0.n4568_cascade_ ));
    InMux I__1277 (
            .O(N__13101),
            .I(N__13098));
    LocalMux I__1276 (
            .O(N__13098),
            .I(\c0.n46 ));
    InMux I__1275 (
            .O(N__13095),
            .I(N__13091));
    InMux I__1274 (
            .O(N__13094),
            .I(N__13088));
    LocalMux I__1273 (
            .O(N__13091),
            .I(N__13084));
    LocalMux I__1272 (
            .O(N__13088),
            .I(N__13081));
    InMux I__1271 (
            .O(N__13087),
            .I(N__13078));
    Span12Mux_s1_h I__1270 (
            .O(N__13084),
            .I(N__13073));
    Span12Mux_s5_v I__1269 (
            .O(N__13081),
            .I(N__13073));
    LocalMux I__1268 (
            .O(N__13078),
            .I(data_in_6_7));
    Odrv12 I__1267 (
            .O(N__13073),
            .I(data_in_6_7));
    InMux I__1266 (
            .O(N__13068),
            .I(N__13065));
    LocalMux I__1265 (
            .O(N__13065),
            .I(\c0.n8816 ));
    CascadeMux I__1264 (
            .O(N__13062),
            .I(\c0.n4282_cascade_ ));
    InMux I__1263 (
            .O(N__13059),
            .I(N__13056));
    LocalMux I__1262 (
            .O(N__13056),
            .I(N__13053));
    Span4Mux_s2_h I__1261 (
            .O(N__13053),
            .I(N__13050));
    Span4Mux_h I__1260 (
            .O(N__13050),
            .I(N__13047));
    Odrv4 I__1259 (
            .O(N__13047),
            .I(\c0.data_in_frame_20_5 ));
    CascadeMux I__1258 (
            .O(N__13044),
            .I(\c0.n4215_cascade_ ));
    CascadeMux I__1257 (
            .O(N__13041),
            .I(\c0.n18_adj_1593_cascade_ ));
    InMux I__1256 (
            .O(N__13038),
            .I(N__13035));
    LocalMux I__1255 (
            .O(N__13035),
            .I(\c0.n20_adj_1596 ));
    CascadeMux I__1254 (
            .O(N__13032),
            .I(\c0.n17_cascade_ ));
    CascadeMux I__1253 (
            .O(N__13029),
            .I(\c0.n4324_cascade_ ));
    InMux I__1252 (
            .O(N__13026),
            .I(N__13023));
    LocalMux I__1251 (
            .O(N__13023),
            .I(\c0.n8951 ));
    CascadeMux I__1250 (
            .O(N__13020),
            .I(\c0.n8951_cascade_ ));
    InMux I__1249 (
            .O(N__13017),
            .I(N__13014));
    LocalMux I__1248 (
            .O(N__13014),
            .I(N__13011));
    Odrv4 I__1247 (
            .O(N__13011),
            .I(\c0.n48 ));
    InMux I__1246 (
            .O(N__13008),
            .I(N__13005));
    LocalMux I__1245 (
            .O(N__13005),
            .I(\c0.n4406 ));
    CascadeMux I__1244 (
            .O(N__13002),
            .I(\c0.n4406_cascade_ ));
    InMux I__1243 (
            .O(N__12999),
            .I(N__12996));
    LocalMux I__1242 (
            .O(N__12996),
            .I(N__12993));
    Odrv4 I__1241 (
            .O(N__12993),
            .I(\c0.n43_adj_1610 ));
    InMux I__1240 (
            .O(N__12990),
            .I(N__12987));
    LocalMux I__1239 (
            .O(N__12987),
            .I(N__12984));
    Span4Mux_h I__1238 (
            .O(N__12984),
            .I(N__12981));
    Odrv4 I__1237 (
            .O(N__12981),
            .I(n1894));
    CascadeMux I__1236 (
            .O(N__12978),
            .I(\c0.n9542_cascade_ ));
    InMux I__1235 (
            .O(N__12975),
            .I(N__12972));
    LocalMux I__1234 (
            .O(N__12972),
            .I(N__12969));
    Span4Mux_v I__1233 (
            .O(N__12969),
            .I(N__12966));
    Odrv4 I__1232 (
            .O(N__12966),
            .I(\c0.n9180 ));
    CascadeMux I__1231 (
            .O(N__12963),
            .I(\c0.n4114_cascade_ ));
    CascadeMux I__1230 (
            .O(N__12960),
            .I(\c0.n8801_cascade_ ));
    InMux I__1229 (
            .O(N__12957),
            .I(N__12954));
    LocalMux I__1228 (
            .O(N__12954),
            .I(N__12948));
    InMux I__1227 (
            .O(N__12953),
            .I(N__12941));
    InMux I__1226 (
            .O(N__12952),
            .I(N__12941));
    InMux I__1225 (
            .O(N__12951),
            .I(N__12941));
    Odrv4 I__1224 (
            .O(N__12948),
            .I(\c0.data_in_field_11 ));
    LocalMux I__1223 (
            .O(N__12941),
            .I(\c0.data_in_field_11 ));
    CascadeMux I__1222 (
            .O(N__12936),
            .I(N__12933));
    InMux I__1221 (
            .O(N__12933),
            .I(N__12930));
    LocalMux I__1220 (
            .O(N__12930),
            .I(\c0.n4276 ));
    CascadeMux I__1219 (
            .O(N__12927),
            .I(\c0.n4276_cascade_ ));
    CascadeMux I__1218 (
            .O(N__12924),
            .I(\c0.n12_adj_1633_cascade_ ));
    InMux I__1217 (
            .O(N__12921),
            .I(N__12917));
    InMux I__1216 (
            .O(N__12920),
            .I(N__12914));
    LocalMux I__1215 (
            .O(N__12917),
            .I(\c0.n4327 ));
    LocalMux I__1214 (
            .O(N__12914),
            .I(\c0.n4327 ));
    CascadeMux I__1213 (
            .O(N__12909),
            .I(\c0.n4434_cascade_ ));
    InMux I__1212 (
            .O(N__12906),
            .I(N__12903));
    LocalMux I__1211 (
            .O(N__12903),
            .I(\c0.n8766 ));
    CascadeMux I__1210 (
            .O(N__12900),
            .I(\c0.n9482_cascade_ ));
    InMux I__1209 (
            .O(N__12897),
            .I(N__12894));
    LocalMux I__1208 (
            .O(N__12894),
            .I(N__12891));
    Span4Mux_v I__1207 (
            .O(N__12891),
            .I(N__12888));
    Odrv4 I__1206 (
            .O(N__12888),
            .I(\c0.n9207 ));
    CascadeMux I__1205 (
            .O(N__12885),
            .I(\c0.n9548_cascade_ ));
    InMux I__1204 (
            .O(N__12882),
            .I(N__12879));
    LocalMux I__1203 (
            .O(N__12879),
            .I(N__12876));
    Span4Mux_s3_v I__1202 (
            .O(N__12876),
            .I(N__12873));
    Span4Mux_v I__1201 (
            .O(N__12873),
            .I(N__12870));
    Odrv4 I__1200 (
            .O(N__12870),
            .I(\c0.n9177 ));
    InMux I__1199 (
            .O(N__12867),
            .I(N__12863));
    InMux I__1198 (
            .O(N__12866),
            .I(N__12858));
    LocalMux I__1197 (
            .O(N__12863),
            .I(N__12855));
    InMux I__1196 (
            .O(N__12862),
            .I(N__12850));
    InMux I__1195 (
            .O(N__12861),
            .I(N__12850));
    LocalMux I__1194 (
            .O(N__12858),
            .I(N__12847));
    Odrv4 I__1193 (
            .O(N__12855),
            .I(\c0.data_in_field_10 ));
    LocalMux I__1192 (
            .O(N__12850),
            .I(\c0.data_in_field_10 ));
    Odrv4 I__1191 (
            .O(N__12847),
            .I(\c0.data_in_field_10 ));
    InMux I__1190 (
            .O(N__12840),
            .I(N__12834));
    InMux I__1189 (
            .O(N__12839),
            .I(N__12834));
    LocalMux I__1188 (
            .O(N__12834),
            .I(data_in_12_7));
    InMux I__1187 (
            .O(N__12831),
            .I(N__12827));
    InMux I__1186 (
            .O(N__12830),
            .I(N__12824));
    LocalMux I__1185 (
            .O(N__12827),
            .I(data_in_13_4));
    LocalMux I__1184 (
            .O(N__12824),
            .I(data_in_13_4));
    InMux I__1183 (
            .O(N__12819),
            .I(N__12813));
    InMux I__1182 (
            .O(N__12818),
            .I(N__12813));
    LocalMux I__1181 (
            .O(N__12813),
            .I(data_in_14_4));
    InMux I__1180 (
            .O(N__12810),
            .I(N__12804));
    InMux I__1179 (
            .O(N__12809),
            .I(N__12804));
    LocalMux I__1178 (
            .O(N__12804),
            .I(data_in_10_0));
    InMux I__1177 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__1176 (
            .O(N__12798),
            .I(N__12794));
    InMux I__1175 (
            .O(N__12797),
            .I(N__12791));
    Odrv4 I__1174 (
            .O(N__12794),
            .I(data_in_11_0));
    LocalMux I__1173 (
            .O(N__12791),
            .I(data_in_11_0));
    InMux I__1172 (
            .O(N__12786),
            .I(\c0.tx2.n8109 ));
    InMux I__1171 (
            .O(N__12783),
            .I(\c0.tx2.n8110 ));
    InMux I__1170 (
            .O(N__12780),
            .I(\c0.tx2.n8111 ));
    InMux I__1169 (
            .O(N__12777),
            .I(bfn_1_32_0_));
    InMux I__1168 (
            .O(N__12774),
            .I(N__12768));
    InMux I__1167 (
            .O(N__12773),
            .I(N__12768));
    LocalMux I__1166 (
            .O(N__12768),
            .I(data_in_7_7));
    InMux I__1165 (
            .O(N__12765),
            .I(N__12759));
    InMux I__1164 (
            .O(N__12764),
            .I(N__12759));
    LocalMux I__1163 (
            .O(N__12759),
            .I(data_in_10_7));
    InMux I__1162 (
            .O(N__12756),
            .I(N__12750));
    InMux I__1161 (
            .O(N__12755),
            .I(N__12750));
    LocalMux I__1160 (
            .O(N__12750),
            .I(data_in_11_7));
    CascadeMux I__1159 (
            .O(N__12747),
            .I(\c0.n9524_cascade_ ));
    InMux I__1158 (
            .O(N__12744),
            .I(N__12741));
    LocalMux I__1157 (
            .O(N__12741),
            .I(\c0.n9183 ));
    CascadeMux I__1156 (
            .O(N__12738),
            .I(\c0.n9186_cascade_ ));
    CascadeMux I__1155 (
            .O(N__12735),
            .I(\c0.n9518_cascade_ ));
    InMux I__1154 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__1153 (
            .O(N__12729),
            .I(N__12726));
    Odrv12 I__1152 (
            .O(N__12726),
            .I(\c0.n22_adj_1680 ));
    CascadeMux I__1151 (
            .O(N__12723),
            .I(\c0.n9521_cascade_ ));
    InMux I__1150 (
            .O(N__12720),
            .I(N__12717));
    LocalMux I__1149 (
            .O(N__12717),
            .I(\c0.tx2.r_Clock_Count_0 ));
    InMux I__1148 (
            .O(N__12714),
            .I(bfn_1_31_0_));
    InMux I__1147 (
            .O(N__12711),
            .I(\c0.tx2.n8105 ));
    InMux I__1146 (
            .O(N__12708),
            .I(\c0.tx2.n8106 ));
    InMux I__1145 (
            .O(N__12705),
            .I(\c0.tx2.n8107 ));
    InMux I__1144 (
            .O(N__12702),
            .I(\c0.tx2.n8108 ));
    CascadeMux I__1143 (
            .O(N__12699),
            .I(\c0.n9464_cascade_ ));
    CascadeMux I__1142 (
            .O(N__12696),
            .I(\c0.n9470_cascade_ ));
    InMux I__1141 (
            .O(N__12693),
            .I(N__12690));
    LocalMux I__1140 (
            .O(N__12690),
            .I(\c0.n9216 ));
    CascadeMux I__1139 (
            .O(N__12687),
            .I(\c0.n9213_cascade_ ));
    InMux I__1138 (
            .O(N__12684),
            .I(N__12681));
    LocalMux I__1137 (
            .O(N__12681),
            .I(N__12678));
    Odrv4 I__1136 (
            .O(N__12678),
            .I(\c0.n9210 ));
    CascadeMux I__1135 (
            .O(N__12675),
            .I(\c0.n9458_cascade_ ));
    CascadeMux I__1134 (
            .O(N__12672),
            .I(\c0.n9461_cascade_ ));
    CascadeMux I__1133 (
            .O(N__12669),
            .I(\c0.n9530_cascade_ ));
    CascadeMux I__1132 (
            .O(N__12666),
            .I(\c0.n54_cascade_ ));
    InMux I__1131 (
            .O(N__12663),
            .I(N__12660));
    LocalMux I__1130 (
            .O(N__12660),
            .I(\c0.n49 ));
    InMux I__1129 (
            .O(N__12657),
            .I(N__12654));
    LocalMux I__1128 (
            .O(N__12654),
            .I(\c0.n9001 ));
    CascadeMux I__1127 (
            .O(N__12651),
            .I(\c0.n9001_cascade_ ));
    CascadeMux I__1126 (
            .O(N__12648),
            .I(\c0.n10_adj_1637_cascade_ ));
    CascadeMux I__1125 (
            .O(N__12645),
            .I(N__12642));
    InMux I__1124 (
            .O(N__12642),
            .I(N__12639));
    LocalMux I__1123 (
            .O(N__12639),
            .I(\c0.data_in_frame_19_3 ));
    CascadeMux I__1122 (
            .O(N__12636),
            .I(\c0.n9686_cascade_ ));
    CascadeMux I__1121 (
            .O(N__12633),
            .I(\c0.n9689_cascade_ ));
    InMux I__1120 (
            .O(N__12630),
            .I(N__12627));
    LocalMux I__1119 (
            .O(N__12627),
            .I(N__12624));
    Odrv4 I__1118 (
            .O(N__12624),
            .I(\c0.n10_adj_1646 ));
    InMux I__1117 (
            .O(N__12621),
            .I(N__12617));
    InMux I__1116 (
            .O(N__12620),
            .I(N__12614));
    LocalMux I__1115 (
            .O(N__12617),
            .I(N__12611));
    LocalMux I__1114 (
            .O(N__12614),
            .I(\c0.n8779 ));
    Odrv4 I__1113 (
            .O(N__12611),
            .I(\c0.n8779 ));
    CascadeMux I__1112 (
            .O(N__12606),
            .I(\c0.n9674_cascade_ ));
    CascadeMux I__1111 (
            .O(N__12603),
            .I(\c0.n9677_cascade_ ));
    InMux I__1110 (
            .O(N__12600),
            .I(N__12597));
    LocalMux I__1109 (
            .O(N__12597),
            .I(N__12594));
    Odrv12 I__1108 (
            .O(N__12594),
            .I(\c0.n4431 ));
    CascadeMux I__1107 (
            .O(N__12591),
            .I(\c0.n8849_cascade_ ));
    CascadeMux I__1106 (
            .O(N__12588),
            .I(\c0.n20_adj_1622_cascade_ ));
    CascadeMux I__1105 (
            .O(N__12585),
            .I(N__12582));
    InMux I__1104 (
            .O(N__12582),
            .I(N__12579));
    LocalMux I__1103 (
            .O(N__12579),
            .I(\c0.data_in_frame_19_5 ));
    CascadeMux I__1102 (
            .O(N__12576),
            .I(\c0.n4431_cascade_ ));
    InMux I__1101 (
            .O(N__12573),
            .I(N__12570));
    LocalMux I__1100 (
            .O(N__12570),
            .I(n1902));
    InMux I__1099 (
            .O(N__12567),
            .I(N__12564));
    LocalMux I__1098 (
            .O(N__12564),
            .I(N__12559));
    InMux I__1097 (
            .O(N__12563),
            .I(N__12556));
    InMux I__1096 (
            .O(N__12562),
            .I(N__12553));
    Span4Mux_v I__1095 (
            .O(N__12559),
            .I(N__12550));
    LocalMux I__1094 (
            .O(N__12556),
            .I(data_in_6_4));
    LocalMux I__1093 (
            .O(N__12553),
            .I(data_in_6_4));
    Odrv4 I__1092 (
            .O(N__12550),
            .I(data_in_6_4));
    CascadeMux I__1091 (
            .O(N__12543),
            .I(\c0.n24_cascade_ ));
    CascadeMux I__1090 (
            .O(N__12540),
            .I(\c0.n4_adj_1594_cascade_ ));
    InMux I__1089 (
            .O(N__12537),
            .I(N__12528));
    InMux I__1088 (
            .O(N__12536),
            .I(N__12528));
    InMux I__1087 (
            .O(N__12535),
            .I(N__12528));
    LocalMux I__1086 (
            .O(N__12528),
            .I(data_in_5_1));
    InMux I__1085 (
            .O(N__12525),
            .I(N__12520));
    InMux I__1084 (
            .O(N__12524),
            .I(N__12515));
    InMux I__1083 (
            .O(N__12523),
            .I(N__12515));
    LocalMux I__1082 (
            .O(N__12520),
            .I(data_in_6_1));
    LocalMux I__1081 (
            .O(N__12515),
            .I(data_in_6_1));
    InMux I__1080 (
            .O(N__12510),
            .I(N__12504));
    InMux I__1079 (
            .O(N__12509),
            .I(N__12504));
    LocalMux I__1078 (
            .O(N__12504),
            .I(data_in_7_1));
    InMux I__1077 (
            .O(N__12501),
            .I(N__12498));
    LocalMux I__1076 (
            .O(N__12498),
            .I(N__12494));
    InMux I__1075 (
            .O(N__12497),
            .I(N__12491));
    Odrv12 I__1074 (
            .O(N__12494),
            .I(data_in_9_1));
    LocalMux I__1073 (
            .O(N__12491),
            .I(data_in_9_1));
    InMux I__1072 (
            .O(N__12486),
            .I(N__12480));
    InMux I__1071 (
            .O(N__12485),
            .I(N__12480));
    LocalMux I__1070 (
            .O(N__12480),
            .I(data_in_8_1));
    InMux I__1069 (
            .O(N__12477),
            .I(N__12471));
    InMux I__1068 (
            .O(N__12476),
            .I(N__12471));
    LocalMux I__1067 (
            .O(N__12471),
            .I(data_in_13_1));
    InMux I__1066 (
            .O(N__12468),
            .I(N__12462));
    InMux I__1065 (
            .O(N__12467),
            .I(N__12462));
    LocalMux I__1064 (
            .O(N__12462),
            .I(data_in_12_1));
    InMux I__1063 (
            .O(N__12459),
            .I(N__12453));
    InMux I__1062 (
            .O(N__12458),
            .I(N__12453));
    LocalMux I__1061 (
            .O(N__12453),
            .I(data_in_7_4));
    InMux I__1060 (
            .O(N__12450),
            .I(N__12444));
    InMux I__1059 (
            .O(N__12449),
            .I(N__12444));
    LocalMux I__1058 (
            .O(N__12444),
            .I(data_in_8_4));
    InMux I__1057 (
            .O(N__12441),
            .I(N__12435));
    InMux I__1056 (
            .O(N__12440),
            .I(N__12435));
    LocalMux I__1055 (
            .O(N__12435),
            .I(data_in_9_4));
    InMux I__1054 (
            .O(N__12432),
            .I(N__12426));
    InMux I__1053 (
            .O(N__12431),
            .I(N__12426));
    LocalMux I__1052 (
            .O(N__12426),
            .I(data_in_10_4));
    InMux I__1051 (
            .O(N__12423),
            .I(N__12417));
    InMux I__1050 (
            .O(N__12422),
            .I(N__12417));
    LocalMux I__1049 (
            .O(N__12417),
            .I(data_in_11_4));
    InMux I__1048 (
            .O(N__12414),
            .I(N__12408));
    InMux I__1047 (
            .O(N__12413),
            .I(N__12408));
    LocalMux I__1046 (
            .O(N__12408),
            .I(data_in_12_4));
    InMux I__1045 (
            .O(N__12405),
            .I(N__12399));
    InMux I__1044 (
            .O(N__12404),
            .I(N__12399));
    LocalMux I__1043 (
            .O(N__12399),
            .I(data_in_10_1));
    InMux I__1042 (
            .O(N__12396),
            .I(N__12390));
    InMux I__1041 (
            .O(N__12395),
            .I(N__12390));
    LocalMux I__1040 (
            .O(N__12390),
            .I(data_in_11_1));
    InMux I__1039 (
            .O(N__12387),
            .I(N__12381));
    InMux I__1038 (
            .O(N__12386),
            .I(N__12381));
    LocalMux I__1037 (
            .O(N__12381),
            .I(data_in_14_1));
    IoInMux I__1036 (
            .O(N__12378),
            .I(N__12375));
    LocalMux I__1035 (
            .O(N__12375),
            .I(N__12372));
    IoSpan4Mux I__1034 (
            .O(N__12372),
            .I(N__12369));
    IoSpan4Mux I__1033 (
            .O(N__12369),
            .I(N__12366));
    IoSpan4Mux I__1032 (
            .O(N__12366),
            .I(N__12363));
    Odrv4 I__1031 (
            .O(N__12363),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_6_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_27_0_));
    defparam IN_MUX_bfv_6_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_28_0_ (
            .carryinitin(n8162),
            .carryinitout(bfn_6_28_0_));
    defparam IN_MUX_bfv_6_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_29_0_ (
            .carryinitin(n8170),
            .carryinitout(bfn_6_29_0_));
    defparam IN_MUX_bfv_6_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_30_0_ (
            .carryinitin(n8178),
            .carryinitout(bfn_6_30_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(\c0.tx2.n8112 ),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_15_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_30_0_));
    defparam IN_MUX_bfv_15_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_31_0_ (
            .carryinitin(\c0.tx.n8097 ),
            .carryinitout(bfn_15_31_0_));
    defparam IN_MUX_bfv_11_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_31_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_16_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_26_0_ (
            .carryinitin(\c0.n8127 ),
            .carryinitout(bfn_16_26_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_11_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_27_0_));
    defparam IN_MUX_bfv_11_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_28_0_ (
            .carryinitin(n8137),
            .carryinitout(bfn_11_28_0_));
    defparam IN_MUX_bfv_11_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_29_0_ (
            .carryinitin(n8145),
            .carryinitout(bfn_11_29_0_));
    defparam IN_MUX_bfv_11_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_30_0_ (
            .carryinitin(n8153),
            .carryinitout(bfn_11_30_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__12378),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.data_in_0___i74_LC_1_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i74_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i74_LC_1_19_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i74_LC_1_19_0  (
            .in0(N__12405),
            .in1(N__29627),
            .in2(_gnd_net_),
            .in3(N__12497),
            .lcout(data_in_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i82_LC_1_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i82_LC_1_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i82_LC_1_19_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i82_LC_1_19_1  (
            .in0(N__12396),
            .in1(_gnd_net_),
            .in2(N__29843),
            .in3(N__12404),
            .lcout(data_in_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i90_LC_1_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i90_LC_1_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i90_LC_1_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i90_LC_1_19_2  (
            .in0(N__29631),
            .in1(N__12468),
            .in2(_gnd_net_),
            .in3(N__12395),
            .lcout(data_in_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i106_LC_1_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i106_LC_1_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i106_LC_1_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i106_LC_1_19_4  (
            .in0(N__12387),
            .in1(N__29626),
            .in2(_gnd_net_),
            .in3(N__12476),
            .lcout(data_in_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i114_LC_1_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i114_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i114_LC_1_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i114_LC_1_19_5  (
            .in0(N__29625),
            .in1(N__16068),
            .in2(_gnd_net_),
            .in3(N__12386),
            .lcout(data_in_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i98_LC_1_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i98_LC_1_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i98_LC_1_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i98_LC_1_19_6  (
            .in0(N__29632),
            .in1(N__12477),
            .in2(_gnd_net_),
            .in3(N__12467),
            .lcout(data_in_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i53_LC_1_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i53_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i53_LC_1_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i53_LC_1_20_0  (
            .in0(N__12459),
            .in1(N__29779),
            .in2(_gnd_net_),
            .in3(N__12562),
            .lcout(data_in_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i61_LC_1_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i61_LC_1_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i61_LC_1_20_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i61_LC_1_20_1  (
            .in0(N__12450),
            .in1(N__29776),
            .in2(_gnd_net_),
            .in3(N__12458),
            .lcout(data_in_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i69_LC_1_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i69_LC_1_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i69_LC_1_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i69_LC_1_20_2  (
            .in0(N__12441),
            .in1(N__29780),
            .in2(_gnd_net_),
            .in3(N__12449),
            .lcout(data_in_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i77_LC_1_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i77_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i77_LC_1_20_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i77_LC_1_20_3  (
            .in0(N__12432),
            .in1(N__29777),
            .in2(_gnd_net_),
            .in3(N__12440),
            .lcout(data_in_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i85_LC_1_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i85_LC_1_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i85_LC_1_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i85_LC_1_20_4  (
            .in0(N__12423),
            .in1(N__29781),
            .in2(_gnd_net_),
            .in3(N__12431),
            .lcout(data_in_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i93_LC_1_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i93_LC_1_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i93_LC_1_20_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i93_LC_1_20_5  (
            .in0(N__12414),
            .in1(N__29778),
            .in2(_gnd_net_),
            .in3(N__12422),
            .lcout(data_in_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i101_LC_1_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i101_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i101_LC_1_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i101_LC_1_20_6  (
            .in0(N__29775),
            .in1(N__12831),
            .in2(_gnd_net_),
            .in3(N__12413),
            .lcout(data_in_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i45_LC_1_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i45_LC_1_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i45_LC_1_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i45_LC_1_21_1  (
            .in0(N__29929),
            .in1(N__12563),
            .in2(_gnd_net_),
            .in3(N__16036),
            .lcout(data_in_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35295),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_41_i1_3_lut_LC_1_22_0 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_41_i1_3_lut_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_41_i1_3_lut_LC_1_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_41_i1_3_lut_LC_1_22_0  (
            .in0(N__12535),
            .in1(N__19601),
            .in2(_gnd_net_),
            .in3(N__23419),
            .lcout(n1902),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i42_LC_1_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i42_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i42_LC_1_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i42_LC_1_22_1  (
            .in0(N__12525),
            .in1(N__12536),
            .in2(_gnd_net_),
            .in3(N__29931),
            .lcout(data_in_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i34_LC_1_22_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i34_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i34_LC_1_22_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i34_LC_1_22_2  (
            .in0(N__12537),
            .in1(_gnd_net_),
            .in2(N__30018),
            .in3(N__13628),
            .lcout(data_in_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_1_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_1_22_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i26_LC_1_22_3  (
            .in0(N__13627),
            .in1(N__29930),
            .in2(_gnd_net_),
            .in3(N__13557),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i50_LC_1_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i50_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i50_LC_1_22_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i50_LC_1_22_4  (
            .in0(N__12524),
            .in1(_gnd_net_),
            .in2(N__30019),
            .in3(N__12510),
            .lcout(data_in_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_49_i1_3_lut_LC_1_22_5 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_49_i1_3_lut_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_49_i1_3_lut_LC_1_22_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.mux_358_Mux_49_i1_3_lut_LC_1_22_5  (
            .in0(N__23418),
            .in1(N__12523),
            .in2(_gnd_net_),
            .in3(N__19856),
            .lcout(n1894),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i58_LC_1_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i58_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i58_LC_1_22_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_0___i58_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(N__12485),
            .in2(N__30020),
            .in3(N__12509),
            .lcout(data_in_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i66_LC_1_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i66_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i66_LC_1_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i66_LC_1_22_7  (
            .in0(N__12486),
            .in1(N__12501),
            .in2(_gnd_net_),
            .in3(N__29932),
            .lcout(data_in_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_677_LC_1_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_677_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_677_LC_1_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_677_LC_1_23_0  (
            .in0(N__24754),
            .in1(N__18601),
            .in2(N__28300),
            .in3(N__28240),
            .lcout(\c0.n4431 ),
            .ltout(\c0.n4431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_511_LC_1_23_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_511_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_511_LC_1_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_511_LC_1_23_1  (
            .in0(N__22358),
            .in1(N__16712),
            .in2(N__12576),
            .in3(N__22476),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_667_LC_1_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_667_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_667_LC_1_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_667_LC_1_23_2  (
            .in0(N__24755),
            .in1(N__16847),
            .in2(_gnd_net_),
            .in3(N__18602),
            .lcout(\c0.n8878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i42_LC_1_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i42_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i42_LC_1_23_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_in_frame_0___i42_LC_1_23_3  (
            .in0(N__24776),
            .in1(N__12573),
            .in2(N__19152),
            .in3(_gnd_net_),
            .lcout(data_in_field_41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35304),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_52_i1_3_lut_LC_1_23_4 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_52_i1_3_lut_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_52_i1_3_lut_LC_1_23_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_52_i1_3_lut_LC_1_23_4  (
            .in0(N__12567),
            .in1(N__24336),
            .in2(_gnd_net_),
            .in3(N__23420),
            .lcout(n1891),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_1_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_658_LC_1_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_658_LC_1_23_6  (
            .in0(N__17305),
            .in1(N__16496),
            .in2(_gnd_net_),
            .in3(N__18716),
            .lcout(\c0.n24 ),
            .ltout(\c0.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_706_LC_1_23_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_706_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_706_LC_1_23_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_706_LC_1_23_7  (
            .in0(N__12921),
            .in1(N__14912),
            .in2(N__12543),
            .in3(N__15085),
            .lcout(\c0.n8858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_1_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_1_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_1_24_0  (
            .in0(N__22674),
            .in1(N__18759),
            .in2(N__22984),
            .in3(N__22200),
            .lcout(),
            .ltout(\c0.n4_adj_1594_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_519_LC_1_24_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_519_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_519_LC_1_24_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i7_4_lut_adj_519_LC_1_24_1  (
            .in0(N__23027),
            .in1(N__22976),
            .in2(N__12540),
            .in3(N__12621),
            .lcout(\c0.n22_adj_1595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i44_LC_1_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i44_LC_1_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i44_LC_1_24_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0___i44_LC_1_24_2  (
            .in0(N__22977),
            .in1(N__19154),
            .in2(_gnd_net_),
            .in3(N__13386),
            .lcout(data_in_field_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35310),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_741_LC_1_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_741_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_741_LC_1_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_741_LC_1_24_3  (
            .in0(N__22199),
            .in1(N__22673),
            .in2(_gnd_net_),
            .in3(N__22972),
            .lcout(\c0.n8766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9512_bdd_4_lut_LC_1_24_4 .C_ON=1'b0;
    defparam \c0.n9512_bdd_4_lut_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.n9512_bdd_4_lut_LC_1_24_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9512_bdd_4_lut_LC_1_24_4  (
            .in0(N__33151),
            .in1(N__12862),
            .in2(N__16779),
            .in3(N__14946),
            .lcout(\c0.n9192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i14_LC_1_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i14_LC_1_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i14_LC_1_24_5 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \c0.data_in_frame_0___i14_LC_1_24_5  (
            .in0(N__23516),
            .in1(N__22207),
            .in2(N__13500),
            .in3(N__19147),
            .lcout(\c0.data_in_field_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35310),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_636_LC_1_24_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_636_LC_1_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_636_LC_1_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_636_LC_1_24_6  (
            .in0(N__15117),
            .in1(N__12861),
            .in2(N__12936),
            .in3(N__22614),
            .lcout(\c0.n10_adj_1646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i11_LC_1_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i11_LC_1_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i11_LC_1_24_7 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \c0.data_in_frame_0___i11_LC_1_24_7  (
            .in0(N__19153),
            .in1(N__14748),
            .in2(N__23558),
            .in3(N__12867),
            .lcout(\c0.data_in_field_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35310),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7970_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7970_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7970_LC_1_25_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7970_LC_1_25_0  (
            .in0(N__19770),
            .in1(N__32985),
            .in2(N__12585),
            .in3(N__32014),
            .lcout(),
            .ltout(\c0.n9674_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9674_bdd_4_lut_LC_1_25_1 .C_ON=1'b0;
    defparam \c0.n9674_bdd_4_lut_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9674_bdd_4_lut_LC_1_25_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9674_bdd_4_lut_LC_1_25_1  (
            .in0(N__32986),
            .in1(N__32606),
            .in2(N__12606),
            .in3(N__19932),
            .lcout(),
            .ltout(\c0.n9677_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2  (
            .in0(N__13059),
            .in1(N__31377),
            .in2(N__12603),
            .in3(N__31204),
            .lcout(\c0.n22_adj_1678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_666_LC_1_25_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_666_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_666_LC_1_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_666_LC_1_25_3  (
            .in0(N__12957),
            .in1(N__14413),
            .in2(_gnd_net_),
            .in3(N__12600),
            .lcout(\c0.n8849 ),
            .ltout(\c0.n8849_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_575_LC_1_25_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_575_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_575_LC_1_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_575_LC_1_25_4  (
            .in0(N__27371),
            .in1(N__22068),
            .in2(N__12591),
            .in3(N__19686),
            .lcout(),
            .ltout(\c0.n20_adj_1622_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i158_LC_1_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i158_LC_1_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i158_LC_1_25_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.data_in_frame_0___i158_LC_1_25_5  (
            .in0(_gnd_net_),
            .in1(N__13215),
            .in2(N__12588),
            .in3(N__21105),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35316),
            .ce(N__29066),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_1_26_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_LC_1_26_0  (
            .in0(_gnd_net_),
            .in1(N__17472),
            .in2(_gnd_net_),
            .in3(N__12620),
            .lcout(),
            .ltout(\c0.n10_adj_1637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i156_LC_1_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i156_LC_1_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i156_LC_1_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i156_LC_1_26_1  (
            .in0(N__26757),
            .in1(N__14160),
            .in2(N__12648),
            .in3(N__20630),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35323),
            .ce(N__29004),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7984_LC_1_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7984_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7984_LC_1_26_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7984_LC_1_26_2  (
            .in0(N__33208),
            .in1(N__15604),
            .in2(N__12645),
            .in3(N__32040),
            .lcout(),
            .ltout(\c0.n9686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9686_bdd_4_lut_LC_1_26_3 .C_ON=1'b0;
    defparam \c0.n9686_bdd_4_lut_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9686_bdd_4_lut_LC_1_26_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9686_bdd_4_lut_LC_1_26_3  (
            .in0(N__17398),
            .in1(N__33209),
            .in2(N__12636),
            .in3(N__23782),
            .lcout(),
            .ltout(\c0.n9689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_1_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_1_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_1_26_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_1_26_4  (
            .in0(N__17847),
            .in1(N__31376),
            .in2(N__12633),
            .in3(N__31231),
            .lcout(\c0.n22_adj_1680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_1_26_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_1_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_1_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_LC_1_26_5  (
            .in0(N__12630),
            .in1(N__14417),
            .in2(_gnd_net_),
            .in3(N__13979),
            .lcout(\c0.n8779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_1_27_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_1_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_1_27_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i8_LC_1_27_0  (
            .in0(N__16973),
            .in1(_gnd_net_),
            .in2(N__30036),
            .in3(N__13903),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_1_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_1_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_1_27_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i16_LC_1_27_1  (
            .in0(N__13838),
            .in1(N__30021),
            .in2(_gnd_net_),
            .in3(N__16972),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_697_LC_1_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_697_LC_1_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_697_LC_1_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_697_LC_1_27_2  (
            .in0(N__22532),
            .in1(N__13008),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(\c0.n6_adj_1654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9476_bdd_4_lut_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.n9476_bdd_4_lut_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.n9476_bdd_4_lut_LC_1_27_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9476_bdd_4_lut_LC_1_27_4  (
            .in0(N__33173),
            .in1(N__24780),
            .in2(N__20310),
            .in3(N__14913),
            .lcout(\c0.n9210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_1_27_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_1_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_1_27_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_0___i32_LC_1_27_5  (
            .in0(N__13733),
            .in1(_gnd_net_),
            .in2(N__14830),
            .in3(N__30022),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_1_27_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_1_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_1_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i24_LC_1_27_6  (
            .in0(N__30024),
            .in1(N__14820),
            .in2(_gnd_net_),
            .in3(N__13837),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i48_LC_1_27_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i48_LC_1_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i48_LC_1_27_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i48_LC_1_27_7  (
            .in0(N__13095),
            .in1(N__30023),
            .in2(_gnd_net_),
            .in3(N__13195),
            .lcout(data_in_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_LC_1_28_0 .C_ON=1'b0;
    defparam \c0.i26_4_lut_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_LC_1_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_LC_1_28_0  (
            .in0(N__13101),
            .in1(N__17274),
            .in2(N__13704),
            .in3(N__13017),
            .lcout(),
            .ltout(\c0.n54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i162_LC_1_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i162_LC_1_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i162_LC_1_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i162_LC_1_28_1  (
            .in0(N__12999),
            .in1(N__22179),
            .in2(N__12666),
            .in3(N__12663),
            .lcout(\c0.data_in_frame_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35337),
            .ce(N__29067),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_1_28_2 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_1_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_1_28_2  (
            .in0(N__27186),
            .in1(N__12657),
            .in2(N__17637),
            .in3(N__18780),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_714_LC_1_28_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_714_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_714_LC_1_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_714_LC_1_28_3  (
            .in0(N__24561),
            .in1(N__18470),
            .in2(N__24503),
            .in3(N__17468),
            .lcout(\c0.n9001 ),
            .ltout(\c0.n9001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_546_LC_1_28_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_546_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_546_LC_1_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_546_LC_1_28_4  (
            .in0(N__25083),
            .in1(N__17832),
            .in2(N__12651),
            .in3(N__15519),
            .lcout(\c0.n28_adj_1612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7795_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7795_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7795_LC_1_29_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7795_LC_1_29_0  (
            .in0(N__33190),
            .in1(N__32041),
            .in2(N__19818),
            .in3(N__21622),
            .lcout(),
            .ltout(\c0.n9464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9464_bdd_4_lut_LC_1_29_1 .C_ON=1'b0;
    defparam \c0.n9464_bdd_4_lut_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9464_bdd_4_lut_LC_1_29_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n9464_bdd_4_lut_LC_1_29_1  (
            .in0(N__27791),
            .in1(N__14181),
            .in2(N__12699),
            .in3(N__33191),
            .lcout(\c0.n9216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7800_LC_1_29_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7800_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7800_LC_1_29_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7800_LC_1_29_2  (
            .in0(N__33192),
            .in1(N__15869),
            .in2(N__17955),
            .in3(N__32042),
            .lcout(),
            .ltout(\c0.n9470_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9470_bdd_4_lut_LC_1_29_3 .C_ON=1'b0;
    defparam \c0.n9470_bdd_4_lut_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9470_bdd_4_lut_LC_1_29_3 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n9470_bdd_4_lut_LC_1_29_3  (
            .in0(N__24490),
            .in1(N__20751),
            .in2(N__12696),
            .in3(N__33193),
            .lcout(),
            .ltout(\c0.n9213_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7810_LC_1_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7810_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7810_LC_1_29_4 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7810_LC_1_29_4  (
            .in0(N__31617),
            .in1(N__12693),
            .in2(N__12687),
            .in3(N__31229),
            .lcout(),
            .ltout(\c0.n9458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9458_bdd_4_lut_LC_1_29_5 .C_ON=1'b0;
    defparam \c0.n9458_bdd_4_lut_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9458_bdd_4_lut_LC_1_29_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n9458_bdd_4_lut_LC_1_29_5  (
            .in0(N__12897),
            .in1(N__12684),
            .in2(N__12675),
            .in3(N__31618),
            .lcout(),
            .ltout(\c0.n9461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_29_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_29_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_1_29_6  (
            .in0(N__31619),
            .in1(N__14019),
            .in2(N__12672),
            .in3(N__32377),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35344),
            .ce(N__32273),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7850_LC_1_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7850_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7850_LC_1_30_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7850_LC_1_30_0  (
            .in0(N__33199),
            .in1(N__14247),
            .in2(N__21894),
            .in3(N__32057),
            .lcout(),
            .ltout(\c0.n9530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9530_bdd_4_lut_LC_1_30_1 .C_ON=1'b0;
    defparam \c0.n9530_bdd_4_lut_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9530_bdd_4_lut_LC_1_30_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n9530_bdd_4_lut_LC_1_30_1  (
            .in0(N__17130),
            .in1(N__17103),
            .in2(N__12669),
            .in3(N__33200),
            .lcout(\c0.n9183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7845_LC_1_30_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7845_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7845_LC_1_30_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7845_LC_1_30_2  (
            .in0(N__33201),
            .in1(N__15669),
            .in2(N__26691),
            .in3(N__32058),
            .lcout(),
            .ltout(\c0.n9524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9524_bdd_4_lut_LC_1_30_3 .C_ON=1'b0;
    defparam \c0.n9524_bdd_4_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9524_bdd_4_lut_LC_1_30_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n9524_bdd_4_lut_LC_1_30_3  (
            .in0(N__23852),
            .in1(N__33202),
            .in2(N__12747),
            .in3(N__17732),
            .lcout(),
            .ltout(\c0.n9186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7865_LC_1_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7865_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7865_LC_1_30_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7865_LC_1_30_4  (
            .in0(N__12744),
            .in1(N__31630),
            .in2(N__12738),
            .in3(N__31230),
            .lcout(),
            .ltout(\c0.n9518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9518_bdd_4_lut_LC_1_30_5 .C_ON=1'b0;
    defparam \c0.n9518_bdd_4_lut_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9518_bdd_4_lut_LC_1_30_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9518_bdd_4_lut_LC_1_30_5  (
            .in0(N__31631),
            .in1(N__12882),
            .in2(N__12735),
            .in3(N__12975),
            .lcout(),
            .ltout(\c0.n9521_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_1_30_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_1_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_1_30_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_1_30_6  (
            .in0(N__12732),
            .in1(N__31632),
            .in2(N__12723),
            .in3(N__32388),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35352),
            .ce(N__32264),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_31_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__12720),
            .in2(_gnd_net_),
            .in3(N__12714),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(\c0.tx2.n8105 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i1_LC_1_31_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i1_LC_1_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_1_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_1_31_1  (
            .in0(_gnd_net_),
            .in1(N__13142),
            .in2(_gnd_net_),
            .in3(N__12711),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx2.n8105 ),
            .carryout(\c0.tx2.n8106 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i2_LC_1_31_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i2_LC_1_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_1_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_1_31_2  (
            .in0(_gnd_net_),
            .in1(N__13167),
            .in2(_gnd_net_),
            .in3(N__12708),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx2.n8106 ),
            .carryout(\c0.tx2.n8107 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_31_3 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__13128),
            .in2(_gnd_net_),
            .in3(N__12705),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx2.n8107 ),
            .carryout(\c0.tx2.n8108 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_31_4 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_1_31_4  (
            .in0(_gnd_net_),
            .in1(N__13116),
            .in2(_gnd_net_),
            .in3(N__12702),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx2.n8108 ),
            .carryout(\c0.tx2.n8109 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_31_5 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_1_31_5  (
            .in0(_gnd_net_),
            .in1(N__13356),
            .in2(_gnd_net_),
            .in3(N__12786),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx2.n8109 ),
            .carryout(\c0.tx2.n8110 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_31_6 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_1_31_6  (
            .in0(_gnd_net_),
            .in1(N__13155),
            .in2(_gnd_net_),
            .in3(N__12783),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx2.n8110 ),
            .carryout(\c0.tx2.n8111 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_31_7 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_1_31_7  (
            .in0(_gnd_net_),
            .in1(N__13341),
            .in2(_gnd_net_),
            .in3(N__12780),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx2.n8111 ),
            .carryout(\c0.tx2.n8112 ),
            .clk(N__35359),
            .ce(N__26876),
            .sr(N__13307));
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_1_32_0  (
            .in0(_gnd_net_),
            .in1(N__13287),
            .in2(_gnd_net_),
            .in3(N__12777),
            .lcout(\c0.tx2.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(N__26880),
            .sr(N__13311));
    defparam \c0.data_in_0___i56_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i56_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i56_LC_2_19_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i56_LC_2_19_0  (
            .in0(N__12774),
            .in1(_gnd_net_),
            .in2(N__29844),
            .in3(N__13087),
            .lcout(data_in_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i64_LC_2_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i64_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i64_LC_2_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i64_LC_2_19_1  (
            .in0(N__29642),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__12773),
            .lcout(data_in_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i80_LC_2_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i80_LC_2_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i80_LC_2_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i80_LC_2_19_3  (
            .in0(N__12765),
            .in1(N__29634),
            .in2(_gnd_net_),
            .in3(N__13409),
            .lcout(data_in_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i88_LC_2_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i88_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i88_LC_2_19_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i88_LC_2_19_4  (
            .in0(N__12756),
            .in1(_gnd_net_),
            .in2(N__29845),
            .in3(N__12764),
            .lcout(data_in_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i96_LC_2_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i96_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i96_LC_2_19_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i96_LC_2_19_5  (
            .in0(N__12840),
            .in1(N__29635),
            .in2(_gnd_net_),
            .in3(N__12755),
            .lcout(data_in_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i104_LC_2_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i104_LC_2_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i104_LC_2_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i104_LC_2_19_6  (
            .in0(N__29633),
            .in1(N__12839),
            .in2(_gnd_net_),
            .in3(N__14499),
            .lcout(data_in_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i109_LC_2_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i109_LC_2_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i109_LC_2_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i109_LC_2_20_0  (
            .in0(N__29570),
            .in1(N__12830),
            .in2(_gnd_net_),
            .in3(N__12819),
            .lcout(data_in_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i73_LC_2_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i73_LC_2_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i73_LC_2_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i73_LC_2_20_4  (
            .in0(N__12810),
            .in1(N__29713),
            .in2(_gnd_net_),
            .in3(N__13532),
            .lcout(data_in_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i117_LC_2_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i117_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i117_LC_2_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i117_LC_2_20_6  (
            .in0(N__29571),
            .in1(N__16335),
            .in2(_gnd_net_),
            .in3(N__12818),
            .lcout(data_in_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i81_LC_2_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i81_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i81_LC_2_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i81_LC_2_20_7  (
            .in0(N__29712),
            .in1(N__12801),
            .in2(_gnd_net_),
            .in3(N__12809),
            .lcout(data_in_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_2_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_2_21_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i3_LC_2_21_4  (
            .in0(N__29492),
            .in1(N__13685),
            .in2(_gnd_net_),
            .in3(N__14747),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_679_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_679_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_679_LC_2_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_679_LC_2_22_0  (
            .in0(N__18449),
            .in1(N__13752),
            .in2(N__13496),
            .in3(N__16642),
            .lcout(\c0.n14_adj_1669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_2_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_2_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_2_22_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_0___i2_LC_2_22_1  (
            .in0(N__29485),
            .in1(_gnd_net_),
            .in2(N__13760),
            .in3(N__16646),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_2_22_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_2_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_2_22_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i10_LC_2_22_2  (
            .in0(N__16750),
            .in1(N__29486),
            .in2(_gnd_net_),
            .in3(N__13753),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i89_LC_2_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i89_LC_2_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i89_LC_2_22_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i89_LC_2_22_3  (
            .in0(N__13470),
            .in1(_gnd_net_),
            .in2(N__29700),
            .in3(N__12797),
            .lcout(data_in_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_2_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_2_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_2_22_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i14_LC_2_22_4  (
            .in0(N__13491),
            .in1(N__29487),
            .in2(_gnd_net_),
            .in3(N__16262),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_2_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_2_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i18_LC_2_22_5  (
            .in0(N__29488),
            .in1(N__13561),
            .in2(_gnd_net_),
            .in3(N__16749),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_683_LC_2_22_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_683_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_683_LC_2_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_683_LC_2_22_6  (
            .in0(N__14831),
            .in1(N__14856),
            .in2(N__13565),
            .in3(N__13684),
            .lcout(\c0.n26_adj_1673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_46_i1_3_lut_LC_2_22_7 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_46_i1_3_lut_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_46_i1_3_lut_LC_2_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_358_Mux_46_i1_3_lut_LC_2_22_7  (
            .in0(N__22305),
            .in1(N__16224),
            .in2(_gnd_net_),
            .in3(N__23325),
            .lcout(n1897),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7870_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7870_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7870_LC_2_23_0 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7870_LC_2_23_0  (
            .in0(N__32038),
            .in1(N__33034),
            .in2(N__28305),
            .in3(N__13792),
            .lcout(),
            .ltout(\c0.n9548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9548_bdd_4_lut_LC_2_23_1 .C_ON=1'b0;
    defparam \c0.n9548_bdd_4_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9548_bdd_4_lut_LC_2_23_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9548_bdd_4_lut_LC_2_23_1  (
            .in0(N__12952),
            .in1(N__33064),
            .in2(N__12885),
            .in3(N__15086),
            .lcout(\c0.n9177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9578_bdd_4_lut_LC_2_23_2 .C_ON=1'b0;
    defparam \c0.n9578_bdd_4_lut_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.n9578_bdd_4_lut_LC_2_23_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n9578_bdd_4_lut_LC_2_23_2  (
            .in0(N__13934),
            .in1(N__33033),
            .in2(N__13581),
            .in3(N__18813),
            .lcout(\c0.n9162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_712_LC_2_23_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_712_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_712_LC_2_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_712_LC_2_23_3  (
            .in0(N__13790),
            .in1(N__13932),
            .in2(N__18857),
            .in3(N__17068),
            .lcout(\c0.n4327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_736_LC_2_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_736_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_736_LC_2_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_736_LC_2_23_4  (
            .in0(N__12866),
            .in1(N__12951),
            .in2(_gnd_net_),
            .in3(N__16839),
            .lcout(\c0.n4224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_731_LC_2_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_731_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_731_LC_2_23_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_731_LC_2_23_5  (
            .in0(N__13791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13933),
            .lcout(),
            .ltout(\c0.n8801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_2_23_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_2_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_2_23_6  (
            .in0(N__13572),
            .in1(N__15137),
            .in2(N__12960),
            .in3(N__16816),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i12_LC_2_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i12_LC_2_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i12_LC_2_23_7 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \c0.data_in_frame_0___i12_LC_2_23_7  (
            .in0(N__12953),
            .in1(N__23429),
            .in2(N__14691),
            .in3(N__19146),
            .lcout(\c0.data_in_field_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35311),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_631_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_631_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_631_LC_2_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_631_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__28229),
            .in2(_gnd_net_),
            .in3(N__15291),
            .lcout(\c0.n4276 ),
            .ltout(\c0.n4276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_598_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_598_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_598_LC_2_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_598_LC_2_24_1  (
            .in0(N__27975),
            .in1(N__17312),
            .in2(N__12927),
            .in3(N__13668),
            .lcout(),
            .ltout(\c0.n12_adj_1633_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_603_LC_2_24_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_603_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_603_LC_2_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_603_LC_2_24_2  (
            .in0(N__21315),
            .in1(N__16728),
            .in2(N__12924),
            .in3(N__12920),
            .lcout(\c0.n4434 ),
            .ltout(\c0.n4434_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_593_LC_2_24_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_593_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_593_LC_2_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_593_LC_2_24_3  (
            .in0(N__18773),
            .in1(N__15845),
            .in2(N__12909),
            .in3(N__12906),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7815_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7815_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7815_LC_2_24_5 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7815_LC_2_24_5  (
            .in0(N__28230),
            .in1(N__32039),
            .in2(N__33174),
            .in3(N__17313),
            .lcout(),
            .ltout(\c0.n9482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9482_bdd_4_lut_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.n9482_bdd_4_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.n9482_bdd_4_lut_LC_2_24_6 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n9482_bdd_4_lut_LC_2_24_6  (
            .in0(N__15293),
            .in1(N__16626),
            .in2(N__12900),
            .in3(N__33115),
            .lcout(\c0.n9207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i50_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i50_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i50_LC_2_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i50_LC_2_24_7  (
            .in0(N__22368),
            .in1(N__12990),
            .in2(_gnd_net_),
            .in3(N__19108),
            .lcout(data_in_field_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7860_LC_2_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7860_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7860_LC_2_25_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7860_LC_2_25_0  (
            .in0(N__17503),
            .in1(N__32891),
            .in2(N__17549),
            .in3(N__31992),
            .lcout(),
            .ltout(\c0.n9542_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9542_bdd_4_lut_LC_2_25_1 .C_ON=1'b0;
    defparam \c0.n9542_bdd_4_lut_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9542_bdd_4_lut_LC_2_25_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n9542_bdd_4_lut_LC_2_25_1  (
            .in0(N__13605),
            .in1(N__32892),
            .in2(N__12978),
            .in3(N__22983),
            .lcout(\c0.n9180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i36_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i36_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i36_LC_2_25_2 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \c0.data_in_frame_0___i36_LC_2_25_2  (
            .in0(N__23484),
            .in1(N__15192),
            .in2(N__19158),
            .in3(N__13606),
            .lcout(\c0.data_in_field_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_2_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_711_LC_2_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_711_LC_2_25_3  (
            .in0(N__21409),
            .in1(N__17502),
            .in2(_gnd_net_),
            .in3(N__15827),
            .lcout(\c0.n8855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_579_LC_2_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_579_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_579_LC_2_25_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_579_LC_2_25_4  (
            .in0(_gnd_net_),
            .in1(N__23781),
            .in2(_gnd_net_),
            .in3(N__26685),
            .lcout(\c0.n4577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_2_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_2_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i9_LC_2_25_5  (
            .in0(N__29614),
            .in1(N__16883),
            .in2(_gnd_net_),
            .in3(N__15261),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_687_LC_2_25_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_687_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_687_LC_2_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_687_LC_2_25_6  (
            .in0(N__17057),
            .in1(N__13604),
            .in2(N__21322),
            .in3(N__14898),
            .lcout(\c0.n4114 ),
            .ltout(\c0.n4114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_664_LC_2_25_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_664_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_664_LC_2_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_664_LC_2_25_7  (
            .in0(_gnd_net_),
            .in1(N__15826),
            .in2(N__12963),
            .in3(N__21367),
            .lcout(\c0.n8864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_2_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_2_26_0  (
            .in0(N__25677),
            .in1(N__13026),
            .in2(N__15351),
            .in3(N__17511),
            .lcout(),
            .ltout(\c0.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i168_LC_2_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i168_LC_2_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i168_LC_2_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i168_LC_2_26_1  (
            .in0(N__32457),
            .in1(N__15681),
            .in2(N__13032),
            .in3(N__14136),
            .lcout(\c0.data_in_frame_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35331),
            .ce(N__29003),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_628_LC_2_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_628_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_628_LC_2_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_628_LC_2_26_2  (
            .in0(N__17228),
            .in1(N__13797),
            .in2(_gnd_net_),
            .in3(N__16379),
            .lcout(\c0.n4324 ),
            .ltout(\c0.n4324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_2_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_2_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_2_26_3  (
            .in0(N__31733),
            .in1(N__27666),
            .in2(N__13029),
            .in3(N__17762),
            .lcout(\c0.n8951 ),
            .ltout(\c0.n8951_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_2_26_4 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_2_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_2_26_4  (
            .in0(N__26787),
            .in1(N__28206),
            .in2(N__13020),
            .in3(N__17204),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_2_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_2_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_2_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_735_LC_2_26_5  (
            .in0(N__31734),
            .in1(N__27667),
            .in2(_gnd_net_),
            .in3(N__17763),
            .lcout(\c0.n4479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_662_LC_2_26_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_662_LC_2_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_662_LC_2_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_662_LC_2_26_6  (
            .in0(N__14942),
            .in1(N__13952),
            .in2(N__17265),
            .in3(N__15087),
            .lcout(\c0.n8930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_680_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_680_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_680_LC_2_27_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_680_LC_2_27_0  (
            .in0(N__16971),
            .in1(N__13813),
            .in2(N__13904),
            .in3(N__13836),
            .lcout(\c0.n14_adj_1670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_703_LC_2_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_703_LC_2_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_703_LC_2_27_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_703_LC_2_27_1  (
            .in0(N__17099),
            .in1(_gnd_net_),
            .in2(N__17603),
            .in3(N__15595),
            .lcout(\c0.n4406 ),
            .ltout(\c0.n4406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_2_27_2 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_2_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_2_27_2  (
            .in0(N__17406),
            .in1(N__27792),
            .in2(N__13002),
            .in3(N__14112),
            .lcout(\c0.n43_adj_1610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i108_LC_2_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i108_LC_2_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i108_LC_2_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i108_LC_2_27_3  (
            .in0(N__19565),
            .in1(N__17728),
            .in2(_gnd_net_),
            .in3(N__29032),
            .lcout(data_in_field_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i90_LC_2_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i90_LC_2_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i90_LC_2_27_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i90_LC_2_27_4  (
            .in0(N__21669),
            .in1(_gnd_net_),
            .in2(N__29069),
            .in3(N__17944),
            .lcout(data_in_field_89),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_580_LC_2_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_580_LC_2_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_580_LC_2_27_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_580_LC_2_27_5  (
            .in0(N__17098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15624),
            .lcout(\c0.n8921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i72_LC_2_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i72_LC_2_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i72_LC_2_27_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0___i72_LC_2_27_6  (
            .in0(N__15625),
            .in1(_gnd_net_),
            .in2(N__29068),
            .in3(N__21085),
            .lcout(data_in_field_71),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i102_LC_2_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i102_LC_2_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i102_LC_2_27_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i102_LC_2_27_7  (
            .in0(N__24158),
            .in1(N__19303),
            .in2(_gnd_net_),
            .in3(N__29031),
            .lcout(data_in_field_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i166_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i166_LC_2_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i166_LC_2_28_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_in_frame_0___i166_LC_2_28_0  (
            .in0(N__15531),
            .in1(N__15350),
            .in2(N__22101),
            .in3(N__13038),
            .lcout(\c0.data_in_frame_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(N__29026),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_2_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_2_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_715_LC_2_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_715_LC_2_28_1  (
            .in0(N__20631),
            .in1(N__26081),
            .in2(_gnd_net_),
            .in3(N__14066),
            .lcout(\c0.n4215 ),
            .ltout(\c0.n4215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_518_LC_2_28_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_518_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_518_LC_2_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_518_LC_2_28_2  (
            .in0(N__13068),
            .in1(N__17358),
            .in2(N__13044),
            .in3(N__16680),
            .lcout(),
            .ltout(\c0.n18_adj_1593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_520_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_520_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_520_LC_2_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_520_LC_2_28_3  (
            .in0(N__14145),
            .in1(N__17966),
            .in2(N__13041),
            .in3(N__22375),
            .lcout(\c0.n20_adj_1596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_611_LC_2_28_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_611_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_611_LC_2_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_611_LC_2_28_4  (
            .in0(N__26409),
            .in1(N__32172),
            .in2(_gnd_net_),
            .in3(N__26329),
            .lcout(),
            .ltout(\c0.n4568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_2_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_2_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_2_28_5  (
            .in0(N__24605),
            .in1(N__15393),
            .in2(N__13104),
            .in3(N__24861),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_47_i1_3_lut_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_47_i1_3_lut_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_47_i1_3_lut_LC_2_29_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_358_Mux_47_i1_3_lut_LC_2_29_0  (
            .in0(N__19506),
            .in1(N__13202),
            .in2(_gnd_net_),
            .in3(N__23266),
            .lcout(n1896),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state__i0_LC_2_29_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state__i0_LC_2_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state__i0_LC_2_29_1 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \c0.FRAME_MATCHER_state__i0_LC_2_29_1  (
            .in0(_gnd_net_),
            .in1(N__23676),
            .in2(N__23326),
            .in3(N__23616),
            .lcout(FRAME_MATCHER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35353),
            .ce(N__20808),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_55_i1_3_lut_LC_2_29_3 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_55_i1_3_lut_LC_2_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_55_i1_3_lut_LC_2_29_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.mux_358_Mux_55_i1_3_lut_LC_2_29_3  (
            .in0(N__23262),
            .in1(N__13094),
            .in2(_gnd_net_),
            .in3(N__19714),
            .lcout(n1888),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4613_3_lut_LC_2_29_4.C_ON=1'b0;
    defparam i4613_3_lut_LC_2_29_4.SEQ_MODE=4'b0000;
    defparam i4613_3_lut_LC_2_29_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 i4613_3_lut_LC_2_29_4 (
            .in0(N__21507),
            .in1(N__16050),
            .in2(_gnd_net_),
            .in3(N__23267),
            .lcout(n6164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_527_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_527_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_527_LC_2_29_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_527_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__24488),
            .in2(_gnd_net_),
            .in3(N__28397),
            .lcout(\c0.n9004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_540_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_540_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_540_LC_2_29_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_540_LC_2_29_6  (
            .in0(_gnd_net_),
            .in1(N__21950),
            .in2(_gnd_net_),
            .in3(N__21893),
            .lcout(\c0.n8816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_642_LC_2_30_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_642_LC_2_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_642_LC_2_30_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_642_LC_2_30_0  (
            .in0(_gnd_net_),
            .in1(N__17589),
            .in2(_gnd_net_),
            .in3(N__15606),
            .lcout(\c0.n8807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_574_LC_2_30_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_574_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_574_LC_2_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_574_LC_2_30_1  (
            .in0(N__15605),
            .in1(N__19635),
            .in2(N__15436),
            .in3(N__27729),
            .lcout(\c0.n4282 ),
            .ltout(\c0.n4282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_2_30_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_LC_2_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13062),
            .in3(N__24560),
            .lcout(\c0.n9007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_629_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_629_LC_2_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_629_LC_2_30_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_629_LC_2_30_3  (
            .in0(_gnd_net_),
            .in1(N__15871),
            .in2(_gnd_net_),
            .in3(N__14246),
            .lcout(),
            .ltout(\c0.n4476_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_576_LC_2_30_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_576_LC_2_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_576_LC_2_30_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_576_LC_2_30_4  (
            .in0(N__13236),
            .in1(N__13224),
            .in2(N__13218),
            .in3(N__21951),
            .lcout(\c0.n19_adj_1623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i40_LC_2_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i40_LC_2_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i40_LC_2_30_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i40_LC_2_30_5  (
            .in0(N__13720),
            .in1(N__29396),
            .in2(_gnd_net_),
            .in3(N__13203),
            .lcout(data_in_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35360),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i82_LC_2_30_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i82_LC_2_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i82_LC_2_30_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i82_LC_2_30_7  (
            .in0(N__19857),
            .in1(N__15872),
            .in2(_gnd_net_),
            .in3(N__29070),
            .lcout(data_in_field_81),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35360),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_31_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_31_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_31_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15782),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_LC_2_31_1 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_LC_2_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_LC_2_31_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx2.i2_2_lut_LC_2_31_1  (
            .in0(_gnd_net_),
            .in1(N__14304),
            .in2(_gnd_net_),
            .in3(N__13283),
            .lcout(\c0.tx2.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_2_31_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_31_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_2_31_2  (
            .in0(N__13285),
            .in1(N__13329),
            .in2(N__14317),
            .in3(N__13263),
            .lcout(r_SM_Main_2_adj_1738),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_2_31_3 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_2_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_2_31_3 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx2.i1_4_lut_LC_2_31_3  (
            .in0(N__13166),
            .in1(N__13154),
            .in2(N__13143),
            .in3(N__13127),
            .lcout(),
            .ltout(\c0.tx2.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5854_4_lut_LC_2_31_4 .C_ON=1'b0;
    defparam \c0.tx2.i5854_4_lut_LC_2_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5854_4_lut_LC_2_31_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx2.i5854_4_lut_LC_2_31_4  (
            .in0(N__13115),
            .in1(N__13355),
            .in2(N__13344),
            .in3(N__13340),
            .lcout(\c0.tx2.n7399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_2_lut_LC_2_31_5 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_2_lut_LC_2_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_2_lut_LC_2_31_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx2.i1_2_lut_2_lut_LC_2_31_5  (
            .in0(_gnd_net_),
            .in1(N__26917),
            .in2(_gnd_net_),
            .in3(N__15940),
            .lcout(\c0.tx2.n4081 ),
            .ltout(\c0.tx2.n4081_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_4_lut_LC_2_31_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_4_lut_LC_2_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_4_lut_LC_2_31_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i2_4_lut_LC_2_31_6  (
            .in0(N__13284),
            .in1(N__14318),
            .in2(N__13323),
            .in3(N__13261),
            .lcout(),
            .ltout(\c0.tx2.n8196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7758_4_lut_4_lut_LC_2_31_7 .C_ON=1'b0;
    defparam \c0.tx2.i7758_4_lut_4_lut_LC_2_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7758_4_lut_4_lut_LC_2_31_7 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \c0.tx2.i7758_4_lut_4_lut_LC_2_31_7  (
            .in0(N__13262),
            .in1(N__13320),
            .in2(N__13314),
            .in3(N__26918),
            .lcout(\c0.tx2.n5146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7404_4_lut_LC_2_32_0 .C_ON=1'b0;
    defparam \c0.tx2.i7404_4_lut_LC_2_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7404_4_lut_LC_2_32_0 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \c0.tx2.i7404_4_lut_LC_2_32_0  (
            .in0(N__26919),
            .in1(N__15941),
            .in2(N__14319),
            .in3(N__14264),
            .lcout(n9075),
            .ltout(n9075_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7412_3_lut_LC_2_32_1 .C_ON=1'b0;
    defparam \c0.tx2.i7412_3_lut_LC_2_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7412_3_lut_LC_2_32_1 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \c0.tx2.i7412_3_lut_LC_2_32_1  (
            .in0(N__15942),
            .in1(_gnd_net_),
            .in2(N__13290),
            .in3(N__13245),
            .lcout(n5346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5868_2_lut_LC_2_32_2 .C_ON=1'b0;
    defparam \c0.tx2.i5868_2_lut_LC_2_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5868_2_lut_LC_2_32_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.i5868_2_lut_LC_2_32_2  (
            .in0(_gnd_net_),
            .in1(N__13286),
            .in2(_gnd_net_),
            .in3(N__13260),
            .lcout(r_SM_Main_2_N_1480_1_adj_1744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_LC_2_32_3 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_2_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_2_32_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_LC_2_32_3  (
            .in0(N__16110),
            .in1(N__14332),
            .in2(_gnd_net_),
            .in3(N__16179),
            .lcout(\c0.tx2.n7236 ),
            .ltout(\c0.tx2.n7236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1673_4_lut_LC_2_32_4 .C_ON=1'b0;
    defparam \c0.tx2.i1673_4_lut_LC_2_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1673_4_lut_LC_2_32_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \c0.tx2.i1673_4_lut_LC_2_32_4  (
            .in0(N__20473),
            .in1(N__15943),
            .in2(N__13239),
            .in3(N__14265),
            .lcout(),
            .ltout(n3220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_2_32_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_2_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_2_32_5 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_2_32_5  (
            .in0(N__14267),
            .in1(N__14315),
            .in2(N__13413),
            .in3(N__26920),
            .lcout(r_SM_Main_0_adj_1740),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_7 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_2_32_7  (
            .in0(N__14266),
            .in1(N__14314),
            .in2(N__15950),
            .in3(N__26921),
            .lcout(r_SM_Main_1_adj_1739),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i72_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i72_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i72_LC_3_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i72_LC_3_19_2  (
            .in0(N__29650),
            .in1(N__13410),
            .in2(_gnd_net_),
            .in3(N__13397),
            .lcout(data_in_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35297),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_43_i1_3_lut_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_43_i1_3_lut_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_43_i1_3_lut_LC_3_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_358_Mux_43_i1_3_lut_LC_3_20_0  (
            .in0(N__19566),
            .in1(N__15215),
            .in2(_gnd_net_),
            .in3(N__23541),
            .lcout(n1900),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i71_LC_3_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i71_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i71_LC_3_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i71_LC_3_20_1  (
            .in0(N__29861),
            .in1(N__14472),
            .in2(_gnd_net_),
            .in3(N__16580),
            .lcout(data_in_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i111_LC_3_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i111_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i111_LC_3_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i111_LC_3_20_2  (
            .in0(N__14613),
            .in1(N__29862),
            .in2(_gnd_net_),
            .in3(N__14441),
            .lcout(data_in_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i52_LC_3_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i52_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i52_LC_3_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i52_LC_3_20_3  (
            .in0(N__29859),
            .in1(N__13374),
            .in2(_gnd_net_),
            .in3(N__14705),
            .lcout(data_in_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_51_i1_3_lut_LC_3_20_4 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_51_i1_3_lut_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_51_i1_3_lut_LC_3_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_51_i1_3_lut_LC_3_20_4  (
            .in0(N__14704),
            .in1(N__19438),
            .in2(_gnd_net_),
            .in3(N__23540),
            .lcout(n1892),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i60_LC_3_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i60_LC_3_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i60_LC_3_20_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i60_LC_3_20_5  (
            .in0(N__13365),
            .in1(_gnd_net_),
            .in2(N__29986),
            .in3(N__13373),
            .lcout(data_in_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i68_LC_3_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i68_LC_3_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i68_LC_3_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i68_LC_3_20_6  (
            .in0(N__29759),
            .in1(N__18129),
            .in2(_gnd_net_),
            .in3(N__13364),
            .lcout(data_in_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i65_LC_3_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i65_LC_3_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i65_LC_3_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i65_LC_3_20_7  (
            .in0(N__29860),
            .in1(N__13533),
            .in2(_gnd_net_),
            .in3(N__13520),
            .lcout(data_in_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i49_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i49_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i49_LC_3_21_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i49_LC_3_21_0  (
            .in0(N__13509),
            .in1(N__29493),
            .in2(_gnd_net_),
            .in3(N__20545),
            .lcout(data_in_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i57_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i57_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i57_LC_3_21_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i57_LC_3_21_1  (
            .in0(N__13521),
            .in1(_gnd_net_),
            .in2(N__29701),
            .in3(N__13508),
            .lcout(data_in_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_3_21_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i6_LC_3_21_2  (
            .in0(N__14555),
            .in1(N__13492),
            .in2(_gnd_net_),
            .in3(N__29497),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i97_LC_3_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i97_LC_3_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i97_LC_3_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i97_LC_3_21_4  (
            .in0(N__29358),
            .in1(N__14796),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(data_in_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_704_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_704_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_704_LC_3_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_704_LC_3_21_5  (
            .in0(N__14993),
            .in1(N__18515),
            .in2(N__14740),
            .in3(N__18552),
            .lcout(\c0.n25_adj_1675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7366_4_lut_LC_3_21_6 .C_ON=1'b0;
    defparam \c0.i7366_4_lut_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7366_4_lut_LC_3_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i7366_4_lut_LC_3_21_6  (
            .in0(N__13455),
            .in1(N__14760),
            .in2(N__13443),
            .in3(N__14754),
            .lcout(),
            .ltout(\c0.n9033_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_723_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_723_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_723_LC_3_21_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_4_lut_adj_723_LC_3_21_7  (
            .in0(N__13434),
            .in1(N__13422),
            .in2(N__13416),
            .in3(N__14532),
            .lcout(\c0.n8449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_3_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_3_22_0  (
            .in0(N__33313),
            .in1(N__26461),
            .in2(N__17636),
            .in3(N__27936),
            .lcout(\c0.n20_adj_1659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i152_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i152_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i152_LC_3_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i152_LC_3_22_1  (
            .in0(N__21089),
            .in1(N__25170),
            .in2(_gnd_net_),
            .in3(N__29064),
            .lcout(data_in_field_151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i21_LC_3_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i21_LC_3_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i21_LC_3_22_2 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \c0.data_in_frame_0___i21_LC_3_22_2  (
            .in0(N__13659),
            .in1(N__23564),
            .in2(N__18519),
            .in3(N__19149),
            .lcout(\c0.data_in_field_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_3_22_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i17_LC_3_22_3  (
            .in0(N__14588),
            .in1(N__29616),
            .in2(_gnd_net_),
            .in3(N__16878),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7895_LC_3_22_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7895_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7895_LC_3_22_4 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7895_LC_3_22_4  (
            .in0(N__13658),
            .in1(N__32000),
            .in2(N__33031),
            .in3(N__18758),
            .lcout(\c0.n9578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_732_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_732_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_732_LC_3_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_732_LC_3_22_5  (
            .in0(_gnd_net_),
            .in1(N__16371),
            .in2(_gnd_net_),
            .in3(N__13657),
            .lcout(\c0.n8794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_3_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_3_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_3_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i15_LC_3_22_7  (
            .in0(N__15027),
            .in1(N__14857),
            .in2(_gnd_net_),
            .in3(N__29615),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i27_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i27_LC_3_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i27_LC_3_23_0 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \c0.data_in_frame_0___i27_LC_3_23_0  (
            .in0(N__23479),
            .in1(N__18551),
            .in2(N__19132),
            .in3(N__16846),
            .lcout(\c0.data_in_field_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i26_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i26_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i26_LC_3_23_1 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_in_frame_0___i26_LC_3_23_1  (
            .in0(N__13566),
            .in1(N__23482),
            .in2(N__28244),
            .in3(N__19084),
            .lcout(\c0.data_in_field_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i33_LC_3_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i33_LC_3_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i33_LC_3_23_2 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \c0.data_in_frame_0___i33_LC_3_23_2  (
            .in0(N__23480),
            .in1(N__18715),
            .in2(N__19133),
            .in3(N__14781),
            .lcout(\c0.data_in_field_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i28_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i28_LC_3_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i28_LC_3_23_3 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_in_frame_0___i28_LC_3_23_3  (
            .in0(N__14994),
            .in1(N__23483),
            .in2(N__28299),
            .in3(N__19085),
            .lcout(\c0.data_in_field_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i3_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i3_LC_3_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i3_LC_3_23_4 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \c0.data_in_frame_0___i3_LC_3_23_4  (
            .in0(N__23481),
            .in1(N__13689),
            .in2(N__19134),
            .in3(N__14941),
            .lcout(\c0.data_in_field_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_3_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_694_LC_3_23_5  (
            .in0(N__13655),
            .in1(N__16358),
            .in2(_gnd_net_),
            .in3(N__16435),
            .lcout(\c0.n4381 ),
            .ltout(\c0.n4381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_685_LC_3_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_685_LC_3_23_6  (
            .in0(N__17069),
            .in1(N__13611),
            .in2(N__13662),
            .in3(N__14004),
            .lcout(\c0.n8899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_583_LC_3_23_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_583_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_583_LC_3_23_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_583_LC_3_23_7  (
            .in0(N__13656),
            .in1(N__16806),
            .in2(N__13938),
            .in3(N__18711),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i1_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i1_LC_3_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i1_LC_3_24_0 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \c0.data_in_frame_0___i1_LC_3_24_0  (
            .in0(N__14520),
            .in1(N__27982),
            .in2(N__23546),
            .in3(N__19045),
            .lcout(\c0.data_in_field_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i7_LC_3_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i7_LC_3_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i7_LC_3_24_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.data_in_frame_0___i7_LC_3_24_1  (
            .in0(N__19040),
            .in1(N__13818),
            .in2(N__16378),
            .in3(N__23478),
            .lcout(\c0.data_in_field_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i34_LC_3_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i34_LC_3_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i34_LC_3_24_2 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \c0.data_in_frame_0___i34_LC_3_24_2  (
            .in0(N__23472),
            .in1(N__19041),
            .in2(N__13638),
            .in3(N__14905),
            .lcout(\c0.data_in_field_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_607_LC_3_24_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_607_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_607_LC_3_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_607_LC_3_24_3  (
            .in0(N__13610),
            .in1(N__15300),
            .in2(N__21375),
            .in3(N__13953),
            .lcout(\c0.n4154 ),
            .ltout(\c0.n4154_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_591_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_591_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_591_LC_3_24_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_591_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13584),
            .in3(N__24785),
            .lcout(\c0.n4200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i6_LC_3_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i6_LC_3_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i6_LC_3_24_5 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.data_in_frame_0___i6_LC_3_24_5  (
            .in0(N__19039),
            .in1(N__14556),
            .in2(N__21326),
            .in3(N__23477),
            .lcout(\c0.data_in_field_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_641_LC_3_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_641_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_641_LC_3_24_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_641_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__15136),
            .in2(_gnd_net_),
            .in3(N__18642),
            .lcout(\c0.n8776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i20_LC_3_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i20_LC_3_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i20_LC_3_24_7 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \c0.data_in_frame_0___i20_LC_3_24_7  (
            .in0(N__14664),
            .in1(N__23473),
            .in2(N__19127),
            .in3(N__13796),
            .lcout(\c0.data_in_field_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_3_25_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_3_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_3_25_0  (
            .in0(N__13876),
            .in1(N__15162),
            .in2(_gnd_net_),
            .in3(N__17006),
            .lcout(),
            .ltout(\c0.n10_adj_1631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_594_LC_3_25_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_594_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_594_LC_3_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_594_LC_3_25_1  (
            .in0(N__28292),
            .in1(N__13770),
            .in2(N__13764),
            .in3(N__15720),
            .lcout(\c0.n8427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i25_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i25_LC_3_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i25_LC_3_25_2 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.data_in_frame_0___i25_LC_3_25_2  (
            .in0(N__19046),
            .in1(N__14589),
            .in2(N__28079),
            .in3(N__23493),
            .lcout(\c0.data_in_field_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i10_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i10_LC_3_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i10_LC_3_25_3 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \c0.data_in_frame_0___i10_LC_3_25_3  (
            .in0(N__13761),
            .in1(N__15294),
            .in2(N__23547),
            .in3(N__19053),
            .lcout(\c0.data_in_field_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i40_LC_3_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i40_LC_3_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i40_LC_3_25_4 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \c0.data_in_frame_0___i40_LC_3_25_4  (
            .in0(N__13737),
            .in1(N__23486),
            .in2(N__19129),
            .in3(N__14409),
            .lcout(\c0.data_in_field_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_3_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_LC_3_25_5  (
            .in0(N__15375),
            .in1(N__23733),
            .in2(N__14637),
            .in3(N__13877),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i35_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i35_LC_3_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i35_LC_3_25_6 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \c0.data_in_frame_0___i35_LC_3_25_6  (
            .in0(N__26982),
            .in1(N__23485),
            .in2(N__19128),
            .in3(N__17067),
            .lcout(\c0.data_in_field_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i5_LC_3_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i5_LC_3_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i5_LC_3_25_7 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \c0.data_in_frame_0___i5_LC_3_25_7  (
            .in0(N__18450),
            .in1(N__13931),
            .in2(N__23548),
            .in3(N__19054),
            .lcout(\c0.data_in_field_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i30_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i30_LC_3_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i30_LC_3_26_0 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_in_frame_0___i30_LC_3_26_0  (
            .in0(N__16554),
            .in1(N__23527),
            .in2(N__21429),
            .in3(N__19125),
            .lcout(\c0.data_in_field_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i8_LC_3_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i8_LC_3_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i8_LC_3_26_1 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \c0.data_in_frame_0___i8_LC_3_26_1  (
            .in0(N__23525),
            .in1(N__13908),
            .in2(N__19151),
            .in3(N__14003),
            .lcout(\c0.data_in_field_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_655_LC_3_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_655_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_655_LC_3_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_655_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__28069),
            .in2(_gnd_net_),
            .in3(N__14399),
            .lcout(\c0.n4131 ),
            .ltout(\c0.n4131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_3_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_700_LC_3_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_700_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__13881),
            .in2(N__13863),
            .in3(N__22615),
            .lcout(\c0.n8927 ),
            .ltout(\c0.n8927_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_3_26_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i5_4_lut_LC_3_26_4  (
            .in0(N__15371),
            .in1(N__18681),
            .in2(N__13860),
            .in3(N__17254),
            .lcout(\c0.n20_adj_1597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i48_LC_3_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i48_LC_3_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i48_LC_3_26_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0___i48_LC_3_26_5  (
            .in0(N__19120),
            .in1(N__13857),
            .in2(_gnd_net_),
            .in3(N__15837),
            .lcout(data_in_field_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i24_LC_3_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i24_LC_3_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i24_LC_3_26_6 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_in_frame_0___i24_LC_3_26_6  (
            .in0(N__13845),
            .in1(N__23526),
            .in2(N__13980),
            .in3(N__19124),
            .lcout(\c0.data_in_field_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_3_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_3_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_3_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i7_LC_3_26_7  (
            .in0(N__29380),
            .in1(N__14865),
            .in2(_gnd_net_),
            .in3(N__13817),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_637_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_637_LC_3_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_637_LC_3_27_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_637_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__19817),
            .in2(_gnd_net_),
            .in3(N__27854),
            .lcout(),
            .ltout(\c0.n10_adj_1647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i154_LC_3_27_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i154_LC_3_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i154_LC_3_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i154_LC_3_27_1  (
            .in0(N__25346),
            .in1(N__15753),
            .in2(N__14055),
            .in3(N__31469),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(N__28996),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8004_LC_3_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8004_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8004_LC_3_27_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_8004_LC_3_27_2  (
            .in0(N__15421),
            .in1(N__33116),
            .in2(N__14052),
            .in3(N__32033),
            .lcout(),
            .ltout(\c0.n9704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9704_bdd_4_lut_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.n9704_bdd_4_lut_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9704_bdd_4_lut_LC_3_27_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9704_bdd_4_lut_LC_3_27_3  (
            .in0(N__33120),
            .in1(N__20629),
            .in2(N__14040),
            .in3(N__17709),
            .lcout(),
            .ltout(\c0.n9707_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_27_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_27_4  (
            .in0(N__31378),
            .in1(N__14037),
            .in2(N__14022),
            .in3(N__31245),
            .lcout(\c0.n22_adj_1682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8014_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8014_LC_3_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8014_LC_3_27_5 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_8014_LC_3_27_5  (
            .in0(N__32032),
            .in1(N__13972),
            .in2(N__33175),
            .in3(N__16500),
            .lcout(),
            .ltout(\c0.n9722_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9722_bdd_4_lut_LC_3_27_6 .C_ON=1'b0;
    defparam \c0.n9722_bdd_4_lut_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.n9722_bdd_4_lut_LC_3_27_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9722_bdd_4_lut_LC_3_27_6  (
            .in0(N__33121),
            .in1(N__13999),
            .in2(N__14007),
            .in3(N__16953),
            .lcout(\c0.n9240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_661_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_661_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_661_LC_3_27_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_661_LC_3_27_7  (
            .in0(N__13998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13971),
            .lcout(\c0.n4514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_513_LC_3_28_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_513_LC_3_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_513_LC_3_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_513_LC_3_28_0  (
            .in0(N__14079),
            .in1(N__14085),
            .in2(N__14073),
            .in3(N__15458),
            .lcout(),
            .ltout(\c0.n18_adj_1589_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_514_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_514_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_514_LC_3_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_514_LC_3_28_1  (
            .in0(N__24606),
            .in1(N__14135),
            .in2(N__14118),
            .in3(N__26082),
            .lcout(),
            .ltout(\c0.n20_adj_1590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i167_LC_3_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i167_LC_3_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i167_LC_3_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i167_LC_3_28_2  (
            .in0(N__22097),
            .in1(N__24351),
            .in2(N__14115),
            .in3(N__18471),
            .lcout(\c0.data_in_frame_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35354),
            .ce(N__29025),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_592_LC_3_28_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_592_LC_3_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_592_LC_3_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_592_LC_3_28_3  (
            .in0(N__14108),
            .in1(N__14094),
            .in2(_gnd_net_),
            .in3(N__22685),
            .lcout(\c0.n8822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_651_LC_3_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_651_LC_3_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_651_LC_3_28_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_651_LC_3_28_4  (
            .in0(_gnd_net_),
            .in1(N__26397),
            .in2(_gnd_net_),
            .in3(N__25481),
            .lcout(\c0.n4448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_742_LC_3_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_742_LC_3_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_742_LC_3_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_742_LC_3_28_5  (
            .in0(N__32118),
            .in1(N__26619),
            .in2(_gnd_net_),
            .in3(N__17942),
            .lcout(\c0.n4445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_739_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_739_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_739_LC_3_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_739_LC_3_28_6  (
            .in0(N__17943),
            .in1(N__17450),
            .in2(N__26627),
            .in3(N__32119),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9650_bdd_4_lut_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.n9650_bdd_4_lut_LC_3_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.n9650_bdd_4_lut_LC_3_29_0 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n9650_bdd_4_lut_LC_3_29_0  (
            .in0(N__15537),
            .in1(N__17756),
            .in2(N__32555),
            .in3(N__33176),
            .lcout(\c0.n9126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i64_LC_3_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i64_LC_3_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i64_LC_3_29_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i64_LC_3_29_1  (
            .in0(N__17595),
            .in1(N__21591),
            .in2(_gnd_net_),
            .in3(N__28990),
            .lcout(data_in_field_63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_717_LC_3_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_717_LC_3_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_717_LC_3_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_717_LC_3_29_2  (
            .in0(N__22016),
            .in1(N__22524),
            .in2(N__24960),
            .in3(N__27853),
            .lcout(\c0.n8896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i45_LC_3_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i45_LC_3_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i45_LC_3_29_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i45_LC_3_29_3  (
            .in0(N__22463),
            .in1(N__14187),
            .in2(_gnd_net_),
            .in3(N__19150),
            .lcout(data_in_field_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_627_LC_3_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_627_LC_3_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_627_LC_3_29_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_627_LC_3_29_4  (
            .in0(_gnd_net_),
            .in1(N__14176),
            .in2(_gnd_net_),
            .in3(N__18057),
            .lcout(\c0.n9016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i106_LC_3_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i106_LC_3_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i106_LC_3_29_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_frame_0___i106_LC_3_29_5  (
            .in0(N__14177),
            .in1(_gnd_net_),
            .in2(N__19611),
            .in3(N__28986),
            .lcout(data_in_field_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i128_LC_3_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i128_LC_3_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i128_LC_3_29_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i128_LC_3_29_6  (
            .in0(N__21590),
            .in1(_gnd_net_),
            .in2(N__29062),
            .in3(N__15558),
            .lcout(data_in_field_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i74_LC_3_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i74_LC_3_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i74_LC_3_29_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i74_LC_3_29_7  (
            .in0(N__19610),
            .in1(N__24489),
            .in2(_gnd_net_),
            .in3(N__28991),
            .lcout(data_in_field_73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_601_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_601_LC_3_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_601_LC_3_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_601_LC_3_30_0  (
            .in0(N__18061),
            .in1(N__19684),
            .in2(N__19737),
            .in3(N__21627),
            .lcout(\c0.n8890 ),
            .ltout(\c0.n8890_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_606_LC_3_30_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_606_LC_3_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_606_LC_3_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_606_LC_3_30_1  (
            .in0(N__24713),
            .in1(N__15740),
            .in2(N__14163),
            .in3(N__22261),
            .lcout(\c0.n14_adj_1638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_720_LC_3_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_720_LC_3_30_2  (
            .in0(N__15666),
            .in1(N__22017),
            .in2(N__15441),
            .in3(N__21549),
            .lcout(\c0.n8936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_600_LC_3_30_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_600_LC_3_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_600_LC_3_30_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_600_LC_3_30_3  (
            .in0(N__21550),
            .in1(N__15440),
            .in2(_gnd_net_),
            .in3(N__15667),
            .lcout(\c0.n4285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i136_LC_3_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i136_LC_3_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i136_LC_3_30_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i136_LC_3_30_4  (
            .in0(N__18062),
            .in1(N__21090),
            .in2(_gnd_net_),
            .in3(N__28992),
            .lcout(data_in_field_135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i84_LC_3_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i84_LC_3_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i84_LC_3_30_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0___i84_LC_3_30_5  (
            .in0(N__14245),
            .in1(_gnd_net_),
            .in2(N__29063),
            .in3(N__19440),
            .lcout(data_in_field_83),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_710_LC_3_30_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_710_LC_3_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_710_LC_3_30_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_710_LC_3_30_6  (
            .in0(N__17446),
            .in1(N__15870),
            .in2(_gnd_net_),
            .in3(N__14244),
            .lcout(\c0.n8785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7885_LC_3_30_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7885_LC_3_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7885_LC_3_30_7 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7885_LC_3_30_7  (
            .in0(N__33137),
            .in1(N__25275),
            .in2(N__21793),
            .in3(N__32031),
            .lcout(\c0.n9572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9656_bdd_4_lut_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.n9656_bdd_4_lut_LC_3_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.n9656_bdd_4_lut_LC_3_31_0 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n9656_bdd_4_lut_LC_3_31_0  (
            .in0(N__33182),
            .in1(N__15636),
            .in2(N__17451),
            .in3(N__14193),
            .lcout(),
            .ltout(\c0.n9123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_8009_LC_3_31_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_8009_LC_3_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_8009_LC_3_31_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_8009_LC_3_31_1  (
            .in0(N__14223),
            .in1(N__31627),
            .in2(N__14214),
            .in3(N__31244),
            .lcout(),
            .ltout(\c0.n9644_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9644_bdd_4_lut_LC_3_31_2 .C_ON=1'b0;
    defparam \c0.n9644_bdd_4_lut_LC_3_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.n9644_bdd_4_lut_LC_3_31_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9644_bdd_4_lut_LC_3_31_2  (
            .in0(N__31628),
            .in1(N__14211),
            .in2(N__14199),
            .in3(N__14376),
            .lcout(),
            .ltout(\c0.n9647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_31_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_31_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_3_31_3  (
            .in0(N__18111),
            .in1(N__31629),
            .in2(N__14196),
            .in3(N__32384),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35376),
            .ce(N__32228),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7955_LC_3_31_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7955_LC_3_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7955_LC_3_31_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7955_LC_3_31_4  (
            .in0(N__27728),
            .in1(N__33177),
            .in2(N__21949),
            .in3(N__32056),
            .lcout(\c0.n9656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_3_31_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_3_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_3_31_5 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_3_31_5  (
            .in0(N__17679),
            .in1(N__17604),
            .in2(N__33203),
            .in3(N__32034),
            .lcout(),
            .ltout(\c0.n9752_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9752_bdd_4_lut_LC_3_31_6 .C_ON=1'b0;
    defparam \c0.n9752_bdd_4_lut_LC_3_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.n9752_bdd_4_lut_LC_3_31_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9752_bdd_4_lut_LC_3_31_6  (
            .in0(N__33181),
            .in1(N__15841),
            .in2(N__14421),
            .in3(N__14418),
            .lcout(\c0.n9120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_7999_LC_3_32_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_7999_LC_3_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_7999_LC_3_32_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_7999_LC_3_32_0  (
            .in0(N__14370),
            .in1(N__32292),
            .in2(N__16109),
            .in3(N__16172),
            .lcout(),
            .ltout(\c0.tx2.n9692_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n9692_bdd_4_lut_LC_3_32_1 .C_ON=1'b0;
    defparam \c0.tx2.n9692_bdd_4_lut_LC_3_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n9692_bdd_4_lut_LC_3_32_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.tx2.n9692_bdd_4_lut_LC_3_32_1  (
            .in0(N__30054),
            .in1(N__14358),
            .in2(N__14346),
            .in3(N__16102),
            .lcout(),
            .ltout(\c0.tx2.n9695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i590722_i1_3_lut_LC_3_32_2 .C_ON=1'b0;
    defparam \c0.tx2.i590722_i1_3_lut_LC_3_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i590722_i1_3_lut_LC_3_32_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.tx2.i590722_i1_3_lut_LC_3_32_2  (
            .in0(_gnd_net_),
            .in1(N__14333),
            .in2(N__14343),
            .in3(N__15891),
            .lcout(),
            .ltout(\c0.tx2.o_Tx_Serial_N_1511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_3_32_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_3_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_3_32_3 .LUT_INIT=16'b1111101001010101;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_3_32_3  (
            .in0(N__14300),
            .in1(_gnd_net_),
            .in2(N__14340),
            .in3(N__15939),
            .lcout(n3_adj_1749),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i657_2_lut_LC_3_32_4 .C_ON=1'b0;
    defparam \c0.tx2.i657_2_lut_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i657_2_lut_LC_3_32_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i657_2_lut_LC_3_32_4  (
            .in0(N__16103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16173),
            .lcout(),
            .ltout(n2207_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_32_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_3_32_5 .LUT_INIT=16'b1001101000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_3_32_5  (
            .in0(N__14334),
            .in1(N__16144),
            .in2(N__14337),
            .in3(N__16121),
            .lcout(r_Bit_Index_2_adj_1741),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35383),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_adj_507_LC_3_32_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_adj_507_LC_3_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_4_lut_adj_507_LC_3_32_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_4_lut_adj_507_LC_3_32_6  (
            .in0(N__15937),
            .in1(N__14299),
            .in2(N__26934),
            .in3(N__20475),
            .lcout(\c0.tx2.n3760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7729_3_lut_4_lut_4_lut_LC_3_32_7 .C_ON=1'b0;
    defparam \c0.tx2.i7729_3_lut_4_lut_4_lut_LC_3_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7729_3_lut_4_lut_4_lut_LC_3_32_7 .LUT_INIT=16'b1100001000000010;
    LogicCell40 \c0.tx2.i7729_3_lut_4_lut_4_lut_LC_3_32_7  (
            .in0(N__20474),
            .in1(N__15938),
            .in2(N__14316),
            .in3(N__14268),
            .lcout(n8747),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i138_LC_4_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i138_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i138_LC_4_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i138_LC_4_17_1  (
            .in0(N__29395),
            .in1(N__20133),
            .in2(_gnd_net_),
            .in3(N__16016),
            .lcout(data_in_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i112_LC_4_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i112_LC_4_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i112_LC_4_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i112_LC_4_18_2  (
            .in0(N__29954),
            .in1(N__15993),
            .in2(_gnd_net_),
            .in3(N__14492),
            .lcout(data_in_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35298),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i127_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i127_LC_4_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i127_LC_4_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i127_LC_4_19_1  (
            .in0(N__29697),
            .in1(N__14481),
            .in2(_gnd_net_),
            .in3(N__14624),
            .lcout(data_in_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35302),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i157_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i157_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i157_LC_4_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i157_LC_4_19_4  (
            .in0(N__29699),
            .in1(N__14601),
            .in2(_gnd_net_),
            .in3(N__16286),
            .lcout(data_in_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35302),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i135_LC_4_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i135_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i135_LC_4_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i135_LC_4_19_7  (
            .in0(N__29698),
            .in1(N__18159),
            .in2(_gnd_net_),
            .in3(N__14480),
            .lcout(data_in_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35302),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i79_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i79_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i79_LC_4_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i79_LC_4_20_0  (
            .in0(N__14460),
            .in1(N__29769),
            .in2(_gnd_net_),
            .in3(N__14471),
            .lcout(data_in_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i87_LC_4_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i87_LC_4_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i87_LC_4_20_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i87_LC_4_20_1  (
            .in0(N__14451),
            .in1(_gnd_net_),
            .in2(N__29955),
            .in3(N__14459),
            .lcout(data_in_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i95_LC_4_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i95_LC_4_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i95_LC_4_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i95_LC_4_20_2  (
            .in0(N__14430),
            .in1(N__29770),
            .in2(_gnd_net_),
            .in3(N__14450),
            .lcout(data_in_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i103_LC_4_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i103_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i103_LC_4_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i103_LC_4_20_3  (
            .in0(N__29766),
            .in1(N__14442),
            .in2(_gnd_net_),
            .in3(N__14429),
            .lcout(data_in_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i119_LC_4_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i119_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i119_LC_4_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i119_LC_4_20_5  (
            .in0(N__29767),
            .in1(N__14625),
            .in2(_gnd_net_),
            .in3(N__14612),
            .lcout(data_in_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_4_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_4_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i25_LC_4_20_6  (
            .in0(N__14583),
            .in1(N__14777),
            .in2(_gnd_net_),
            .in3(N__29774),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i165_LC_4_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i165_LC_4_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i165_LC_4_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i165_LC_4_20_7  (
            .in0(N__29768),
            .in1(N__20418),
            .in2(_gnd_net_),
            .in3(N__14600),
            .lcout(data_in_20_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_678_LC_4_21_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_678_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_678_LC_4_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_adj_678_LC_4_21_0  (
            .in0(N__15018),
            .in1(N__16542),
            .in2(N__14584),
            .in3(N__14551),
            .lcout(),
            .ltout(\c0.n28_adj_1668_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_684_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_684_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_684_LC_4_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_684_LC_4_21_1  (
            .in0(N__16760),
            .in1(N__16518),
            .in2(N__14535),
            .in3(N__14526),
            .lcout(\c0.n30_adj_1674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_4_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i6_2_lut_LC_4_21_2  (
            .in0(_gnd_net_),
            .in1(N__18573),
            .in2(_gnd_net_),
            .in3(N__14512),
            .lcout(\c0.n22_adj_1667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_4_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_4_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_4_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i23_LC_4_21_3  (
            .in0(N__15022),
            .in1(N__16520),
            .in2(_gnd_net_),
            .in3(N__29393),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_4_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_4_21_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i31_LC_4_21_4  (
            .in0(N__16519),
            .in1(_gnd_net_),
            .in2(N__29623),
            .in3(N__16196),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_4_21_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_4_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_4_21_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i1_LC_4_21_5  (
            .in0(N__14513),
            .in1(N__29389),
            .in2(_gnd_net_),
            .in3(N__15267),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i105_LC_4_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i105_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i105_LC_4_21_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i105_LC_4_21_6  (
            .in0(N__29388),
            .in1(N__14792),
            .in2(_gnd_net_),
            .in3(N__18411),
            .lcout(data_in_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i33_LC_4_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i33_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i33_LC_4_21_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i33_LC_4_21_7  (
            .in0(N__29840),
            .in1(N__14776),
            .in2(_gnd_net_),
            .in3(N__20526),
            .lcout(data_in_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_681_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_681_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_681_LC_4_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i5_4_lut_adj_681_LC_4_22_0  (
            .in0(N__18379),
            .in1(N__19185),
            .in2(N__16879),
            .in3(N__15263),
            .lcout(\c0.n13_adj_1671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_682_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_682_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_682_LC_4_22_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i5_4_lut_adj_682_LC_4_22_1  (
            .in0(N__15100),
            .in1(N__14652),
            .in2(N__16255),
            .in3(N__14679),
            .lcout(\c0.n13_adj_1672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_4_22_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i11_LC_4_22_2  (
            .in0(N__18380),
            .in1(N__29956),
            .in2(_gnd_net_),
            .in3(N__14733),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i44_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i44_LC_4_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i44_LC_4_22_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i44_LC_4_22_3  (
            .in0(N__14709),
            .in1(_gnd_net_),
            .in2(N__30028),
            .in3(N__15211),
            .lcout(data_in_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_4_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_4_22_4 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \c0.data_in_0___i12_LC_4_22_4  (
            .in0(N__14680),
            .in1(N__29964),
            .in2(N__14660),
            .in3(_gnd_net_),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_4_22_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i4_LC_4_22_5  (
            .in0(N__15101),
            .in1(_gnd_net_),
            .in2(N__30029),
            .in3(N__14681),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_4_22_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i20_LC_4_22_6  (
            .in0(N__14653),
            .in1(N__29957),
            .in2(_gnd_net_),
            .in3(N__14989),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_572_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_572_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_572_LC_4_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_572_LC_4_22_7  (
            .in0(_gnd_net_),
            .in1(N__21234),
            .in2(_gnd_net_),
            .in3(N__25166),
            .lcout(\c0.n4495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i22_LC_4_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i22_LC_4_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i22_LC_4_23_0 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \c0.data_in_frame_0___i22_LC_4_23_0  (
            .in0(N__23560),
            .in1(N__19066),
            .in2(N__16263),
            .in3(N__21357),
            .lcout(\c0.data_in_field_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_614_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_614_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_614_LC_4_23_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_614_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(N__16458),
            .in2(_gnd_net_),
            .in3(N__14934),
            .lcout(\c0.n8902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_4_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_708_LC_4_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_708_LC_4_23_2  (
            .in0(N__14897),
            .in1(N__15063),
            .in2(_gnd_net_),
            .in3(N__28041),
            .lcout(),
            .ltout(\c0.n6_adj_1632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_596_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_596_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_596_LC_4_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_596_LC_4_23_3  (
            .in0(N__16697),
            .in1(N__16805),
            .in2(N__14874),
            .in3(N__14871),
            .lcout(\c0.n4107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_695_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_695_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_695_LC_4_23_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_695_LC_4_23_4  (
            .in0(N__18707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16487),
            .lcout(\c0.n8804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i15_LC_4_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i15_LC_4_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i15_LC_4_23_5 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_in_frame_0___i15_LC_4_23_5  (
            .in0(N__14861),
            .in1(N__23562),
            .in2(N__16413),
            .in3(N__19088),
            .lcout(\c0.data_in_field_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i32_LC_4_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i32_LC_4_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i32_LC_4_23_6 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \c0.data_in_frame_0___i32_LC_4_23_6  (
            .in0(N__23561),
            .in1(N__19067),
            .in2(N__14835),
            .in3(N__16488),
            .lcout(\c0.data_in_field_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i19_LC_4_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i19_LC_4_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i19_LC_4_23_7 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_in_frame_0___i19_LC_4_23_7  (
            .in0(N__18384),
            .in1(N__23563),
            .in2(N__16818),
            .in3(N__19089),
            .lcout(\c0.data_in_field_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i39_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i39_LC_4_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i39_LC_4_24_0 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_in_frame_0___i39_LC_4_24_0  (
            .in0(N__16203),
            .in1(N__23470),
            .in2(N__22619),
            .in3(N__19087),
            .lcout(\c0.data_in_field_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_728_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_728_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_728_LC_4_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_728_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__18636),
            .in2(_gnd_net_),
            .in3(N__25603),
            .lcout(\c0.n4127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i4_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i4_LC_4_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i4_LC_4_24_2 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \c0.data_in_frame_0___i4_LC_4_24_2  (
            .in0(N__19065),
            .in1(N__23471),
            .in2(N__15108),
            .in3(N__15084),
            .lcout(\c0.data_in_field_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_534_LC_4_24_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_534_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_534_LC_4_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i13_4_lut_adj_534_LC_4_24_3  (
            .in0(N__15045),
            .in1(N__15036),
            .in2(N__16659),
            .in3(N__17019),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i38_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i38_LC_4_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i38_LC_4_24_4 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \c0.data_in_frame_0___i38_LC_4_24_4  (
            .in0(N__25604),
            .in1(N__23469),
            .in2(N__18300),
            .in3(N__19086),
            .lcout(data_in_field_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7399_4_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.i7399_4_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7399_4_lut_LC_4_24_5 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \c0.i7399_4_lut_LC_4_24_5  (
            .in0(N__23668),
            .in1(N__20822),
            .in2(N__23545),
            .in3(N__20776),
            .lcout(n9069),
            .ltout(n9069_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i23_LC_4_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i23_LC_4_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i23_LC_4_24_6 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \c0.data_in_frame_0___i23_LC_4_24_6  (
            .in0(N__15026),
            .in1(N__23468),
            .in2(N__14997),
            .in3(N__16439),
            .lcout(\c0.data_in_field_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_4_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_4_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_4_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i28_LC_4_24_7  (
            .in0(N__29394),
            .in1(N__15185),
            .in2(_gnd_net_),
            .in3(N__14985),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_4_25_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_4_25_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_4_25_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 i1_2_lut_3_lut_LC_4_25_0 (
            .in0(N__22778),
            .in1(_gnd_net_),
            .in2(N__25612),
            .in3(N__18640),
            .lcout(),
            .ltout(n4_adj_1750_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_4_25_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_4_25_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i3_4_lut_LC_4_25_1  (
            .in0(N__25640),
            .in1(N__14958),
            .in2(N__14949),
            .in3(N__18858),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i52_LC_4_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i52_LC_4_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i52_LC_4_25_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i52_LC_4_25_2  (
            .in0(N__15327),
            .in1(N__17501),
            .in2(_gnd_net_),
            .in3(N__19064),
            .lcout(data_in_field_51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i53_LC_4_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i53_LC_4_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i53_LC_4_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_frame_0___i53_LC_4_25_3  (
            .in0(N__25262),
            .in1(N__19126),
            .in2(_gnd_net_),
            .in3(N__15315),
            .lcout(data_in_field_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_650_LC_4_25_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_650_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_650_LC_4_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_650_LC_4_25_4  (
            .in0(N__22777),
            .in1(N__22604),
            .in2(N__25611),
            .in3(N__28009),
            .lcout(\c0.n8831 ),
            .ltout(\c0.n8831_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_656_LC_4_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_656_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_656_LC_4_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_656_LC_4_25_5  (
            .in0(N__15160),
            .in1(N__15292),
            .in2(N__15270),
            .in3(N__16434),
            .lcout(\c0.n4183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i9_LC_4_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i9_LC_4_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i9_LC_4_25_6 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_in_frame_0___i9_LC_4_25_6  (
            .in0(N__15262),
            .in1(N__23451),
            .in2(N__28019),
            .in3(N__19063),
            .lcout(\c0.data_in_field_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i56_LC_4_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i56_LC_4_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i56_LC_4_25_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0___i56_LC_4_25_7  (
            .in0(N__19062),
            .in1(N__15231),
            .in2(_gnd_net_),
            .in3(N__17671),
            .lcout(data_in_field_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i36_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i36_LC_4_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i36_LC_4_26_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i36_LC_4_26_0  (
            .in0(N__15178),
            .in1(N__29624),
            .in2(_gnd_net_),
            .in3(N__15216),
            .lcout(data_in_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_554_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_554_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_554_LC_4_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_554_LC_4_26_1  (
            .in0(N__24442),
            .in1(N__15414),
            .in2(_gnd_net_),
            .in3(N__22728),
            .lcout(\c0.n4556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_609_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_609_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_609_LC_4_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_609_LC_4_26_2  (
            .in0(N__18606),
            .in1(N__15161),
            .in2(N__15144),
            .in3(N__17153),
            .lcout(),
            .ltout(\c0.n10_adj_1640_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_4_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_4_26_3  (
            .in0(N__22675),
            .in1(N__16412),
            .in2(N__15477),
            .in3(N__15474),
            .lcout(\c0.n8933 ),
            .ltout(\c0.n8933_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_4_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_LC_4_26_4  (
            .in0(_gnd_net_),
            .in1(N__21410),
            .in2(N__15462),
            .in3(N__15491),
            .lcout(),
            .ltout(\c0.n8314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_538_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_538_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_538_LC_4_26_5 .LUT_INIT=16'b1111111111111001;
    LogicCell40 \c0.i8_4_lut_adj_538_LC_4_26_5  (
            .in0(N__24441),
            .in1(N__15459),
            .in2(N__15444),
            .in3(N__27233),
            .lcout(\c0.n23_adj_1608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i146_LC_4_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i146_LC_4_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i146_LC_4_26_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_frame_0___i146_LC_4_26_6  (
            .in0(N__15415),
            .in1(_gnd_net_),
            .in2(N__21044),
            .in3(N__28772),
            .lcout(data_in_field_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_555_LC_4_27_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_555_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_555_LC_4_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_555_LC_4_27_0  (
            .in0(N__21233),
            .in1(N__15386),
            .in2(N__15568),
            .in3(N__17125),
            .lcout(\c0.n8974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_645_LC_4_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_645_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_645_LC_4_27_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_645_LC_4_27_1  (
            .in0(N__24781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22468),
            .lcout(\c0.n8861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_526_LC_4_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_526_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_526_LC_4_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_526_LC_4_27_2  (
            .in0(_gnd_net_),
            .in1(N__22407),
            .in2(_gnd_net_),
            .in3(N__17124),
            .lcout(\c0.n4452 ),
            .ltout(\c0.n4452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_4_27_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_4_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_4_27_3  (
            .in0(N__23762),
            .in1(N__15360),
            .in2(N__15354),
            .in3(N__17393),
            .lcout(\c0.n8906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_702_LC_4_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_702_LC_4_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_702_LC_4_27_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_702_LC_4_27_4  (
            .in0(N__21881),
            .in1(_gnd_net_),
            .in2(N__15569),
            .in3(N__24943),
            .lcout(\c0.n4253 ),
            .ltout(\c0.n4253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_531_LC_4_27_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_531_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_531_LC_4_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_531_LC_4_27_5  (
            .in0(N__23845),
            .in1(N__15645),
            .in2(N__15639),
            .in3(N__15635),
            .lcout(\c0.n24_adj_1607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i148_LC_4_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i148_LC_4_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i148_LC_4_27_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i148_LC_4_27_6  (
            .in0(_gnd_net_),
            .in1(N__21155),
            .in2(N__29055),
            .in3(N__15594),
            .lcout(data_in_field_147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35355),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i132_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i132_LC_4_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i132_LC_4_27_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_frame_0___i132_LC_4_27_7  (
            .in0(N__21154),
            .in1(_gnd_net_),
            .in2(N__23775),
            .in3(N__28968),
            .lcout(data_in_field_131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35355),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7950_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7950_LC_4_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7950_LC_4_28_0 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7950_LC_4_28_0  (
            .in0(N__32007),
            .in1(N__33189),
            .in2(N__15570),
            .in3(N__25741),
            .lcout(\c0.n9650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_4_lut_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_4_lut_LC_4_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_4_lut_LC_4_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_2_lut_4_lut_LC_4_28_1  (
            .in0(N__26690),
            .in1(N__17541),
            .in2(N__21126),
            .in3(N__17593),
            .lcout(\c0.n16_adj_1598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_734_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_734_LC_4_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_734_LC_4_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_734_LC_4_28_2  (
            .in0(N__17540),
            .in1(N__17594),
            .in2(_gnd_net_),
            .in3(N__26689),
            .lcout(\c0.n8980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i60_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i60_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i60_LC_4_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i60_LC_4_28_3  (
            .in0(N__26728),
            .in1(N__17542),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(data_in_field_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_633_LC_4_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_633_LC_4_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_633_LC_4_28_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_633_LC_4_28_4  (
            .in0(N__19910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25740),
            .lcout(),
            .ltout(\c0.n6_adj_1645_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_634_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_634_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_634_LC_4_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_634_LC_4_28_5  (
            .in0(N__15518),
            .in1(N__21690),
            .in2(N__15498),
            .in3(N__15495),
            .lcout(\c0.n8788 ),
            .ltout(\c0.n8788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_638_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_638_LC_4_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_638_LC_4_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_638_LC_4_28_6  (
            .in0(N__27269),
            .in1(N__32508),
            .in2(N__15756),
            .in3(N__25553),
            .lcout(\c0.n14_adj_1648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_523_LC_4_29_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_523_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_523_LC_4_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_523_LC_4_29_0  (
            .in0(N__26291),
            .in1(N__26031),
            .in2(N__15747),
            .in3(N__21821),
            .lcout(),
            .ltout(\c0.n24_adj_1600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_4_29_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_4_29_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_4_29_1  (
            .in0(N__15726),
            .in1(N__26556),
            .in2(N__15729),
            .in3(N__24860),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_LC_4_29_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_LC_4_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_LC_4_29_2  (
            .in0(N__25718),
            .in1(N__21880),
            .in2(_gnd_net_),
            .in3(N__24948),
            .lcout(\c0.n18_adj_1603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_605_LC_4_29_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_605_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_605_LC_4_29_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_605_LC_4_29_3  (
            .in0(_gnd_net_),
            .in1(N__22467),
            .in2(_gnd_net_),
            .in3(N__15719),
            .lcout(\c0.tx2_transmit_N_1334 ),
            .ltout(\c0.tx2_transmit_N_1334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_524_LC_4_29_4 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_524_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_524_LC_4_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_524_LC_4_29_4  (
            .in0(N__28344),
            .in1(N__22749),
            .in2(N__15702),
            .in3(N__24903),
            .lcout(),
            .ltout(\c0.n22_adj_1601_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i165_LC_4_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i165_LC_4_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i165_LC_4_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i165_LC_4_29_5  (
            .in0(N__15699),
            .in1(N__18009),
            .in2(N__15690),
            .in3(N__15687),
            .lcout(\c0.data_in_frame_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35370),
            .ce(N__28997),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_4_30_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_4_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_4_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_4_30_0  (
            .in0(N__15801),
            .in1(N__19927),
            .in2(N__21966),
            .in3(N__15879),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i116_LC_4_30_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i116_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i116_LC_4_30_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i116_LC_4_30_1  (
            .in0(N__19439),
            .in1(N__15668),
            .in2(_gnd_net_),
            .in3(N__28985),
            .lcout(data_in_field_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_648_LC_4_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_648_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_648_LC_4_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_648_LC_4_30_2  (
            .in0(_gnd_net_),
            .in1(N__19473),
            .in2(_gnd_net_),
            .in3(N__25276),
            .lcout(),
            .ltout(\c0.n4574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_558_LC_4_30_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_558_LC_4_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_558_LC_4_30_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_558_LC_4_30_3  (
            .in0(N__25808),
            .in1(N__21787),
            .in2(N__15882),
            .in3(N__26345),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_4_30_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_4_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_4_30_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_4_30_4  (
            .in0(_gnd_net_),
            .in1(N__17435),
            .in2(_gnd_net_),
            .in3(N__15878),
            .lcout(\c0.n24_adj_1615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i105_LC_4_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i105_LC_4_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i105_LC_4_30_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i105_LC_4_30_5  (
            .in0(N__19474),
            .in1(N__20675),
            .in2(_gnd_net_),
            .in3(N__28984),
            .lcout(data_in_field_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_539_LC_4_30_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_539_LC_4_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_539_LC_4_30_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_539_LC_4_30_7  (
            .in0(_gnd_net_),
            .in1(N__26206),
            .in2(_gnd_net_),
            .in3(N__27879),
            .lcout(\c0.n8909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_613_LC_4_31_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_613_LC_4_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_613_LC_4_31_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_613_LC_4_31_0  (
            .in0(_gnd_net_),
            .in1(N__21432),
            .in2(_gnd_net_),
            .in3(N__15846),
            .lcout(\c0.n8945 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_570_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_570_LC_4_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_570_LC_4_31_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_570_LC_4_31_1  (
            .in0(_gnd_net_),
            .in1(N__24183),
            .in2(_gnd_net_),
            .in3(N__24299),
            .lcout(\c0.n8825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_552_LC_4_31_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_552_LC_4_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_552_LC_4_31_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_552_LC_4_31_3  (
            .in0(N__21891),
            .in1(_gnd_net_),
            .in2(N__20750),
            .in3(N__21730),
            .lcout(\c0.n4333 ),
            .ltout(\c0.n4333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_729_LC_4_31_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_729_LC_4_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_729_LC_4_31_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_729_LC_4_31_4  (
            .in0(N__24300),
            .in1(_gnd_net_),
            .in2(N__15795),
            .in3(N__27328),
            .lcout(\c0.n8998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_5 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_4_31_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_4_31_5  (
            .in0(N__26938),
            .in1(N__15769),
            .in2(_gnd_net_),
            .in3(N__15792),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_559_LC_4_31_6 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_559_LC_4_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_559_LC_4_31_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_559_LC_4_31_6  (
            .in0(N__31685),
            .in1(N__15963),
            .in2(N__23916),
            .in3(N__15957),
            .lcout(\c0.n38_adj_1616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_LC_4_31_7 .C_ON=1'b0;
    defparam \c0.i8_3_lut_LC_4_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_LC_4_31_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i8_3_lut_LC_4_31_7  (
            .in0(N__21554),
            .in1(N__27098),
            .in2(_gnd_net_),
            .in3(N__21731),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_0 .LUT_INIT=16'b1011000111110000;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_4_32_0  (
            .in0(N__26943),
            .in1(N__15951),
            .in2(N__20495),
            .in3(N__15906),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_4_32_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_4_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_4_32_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_4_32_1  (
            .in0(N__15900),
            .in1(N__22872),
            .in2(N__16107),
            .in3(N__16171),
            .lcout(),
            .ltout(\c0.tx2.n9716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n9716_bdd_4_lut_LC_4_32_2 .C_ON=1'b0;
    defparam \c0.tx2.n9716_bdd_4_lut_LC_4_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n9716_bdd_4_lut_LC_4_32_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.tx2.n9716_bdd_4_lut_LC_4_32_2  (
            .in0(N__25365),
            .in1(N__20010),
            .in2(N__15894),
            .in3(N__16095),
            .lcout(\c0.tx2.n9719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_4_32_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_4_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_4_32_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_4_32_3  (
            .in0(N__16177),
            .in1(N__16145),
            .in2(_gnd_net_),
            .in3(N__16127),
            .lcout(r_Bit_Index_0_adj_1743),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_4_lut_LC_4_32_4.C_ON=1'b0;
    defparam i13_4_lut_4_lut_LC_4_32_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_4_lut_LC_4_32_4.LUT_INIT=16'b0010000001010101;
    LogicCell40 i13_4_lut_4_lut_LC_4_32_4 (
            .in0(N__30789),
            .in1(N__30647),
            .in2(N__30579),
            .in3(N__30723),
            .lcout(),
            .ltout(n4691_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_4_32_5  (
            .in0(N__30648),
            .in1(N__29254),
            .in2(N__15885),
            .in3(N__30790),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam i7769_2_lut_3_lut_LC_4_32_6.C_ON=1'b0;
    defparam i7769_2_lut_3_lut_LC_4_32_6.SEQ_MODE=4'b0000;
    defparam i7769_2_lut_3_lut_LC_4_32_6.LUT_INIT=16'b1101110111111111;
    LogicCell40 i7769_2_lut_3_lut_LC_4_32_6 (
            .in0(N__30788),
            .in1(N__30646),
            .in2(_gnd_net_),
            .in3(N__30722),
            .lcout(n8761),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_32_7 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_4_32_7  (
            .in0(N__16178),
            .in1(N__16146),
            .in2(N__16108),
            .in3(N__16128),
            .lcout(r_Bit_Index_1_adj_1742),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i122_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i122_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i122_LC_5_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i122_LC_5_17_2  (
            .in0(N__29883),
            .in1(N__16005),
            .in2(_gnd_net_),
            .in3(N__16061),
            .lcout(data_in_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i132_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i132_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i132_LC_5_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i132_LC_5_18_1  (
            .in0(N__29953),
            .in1(N__18210),
            .in2(_gnd_net_),
            .in3(N__18230),
            .lcout(data_in_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i141_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i141_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i141_LC_5_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i141_LC_5_18_2  (
            .in0(N__29884),
            .in1(N__16275),
            .in2(_gnd_net_),
            .in3(N__16316),
            .lcout(data_in_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i37_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i37_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i37_LC_5_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i37_LC_5_18_6  (
            .in0(N__29885),
            .in1(N__16900),
            .in2(_gnd_net_),
            .in3(N__16049),
            .lcout(data_in_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i130_LC_5_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i130_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i130_LC_5_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i130_LC_5_18_7  (
            .in0(N__16017),
            .in1(N__29886),
            .in2(_gnd_net_),
            .in3(N__16004),
            .lcout(data_in_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i120_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i120_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i120_LC_5_19_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i120_LC_5_19_0  (
            .in0(N__15981),
            .in1(N__29645),
            .in2(_gnd_net_),
            .in3(N__15992),
            .lcout(data_in_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i128_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i128_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i128_LC_5_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i128_LC_5_19_1  (
            .in0(N__15972),
            .in1(N__29649),
            .in2(_gnd_net_),
            .in3(N__15980),
            .lcout(data_in_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i136_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i136_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i136_LC_5_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i136_LC_5_19_2  (
            .in0(N__29647),
            .in1(N__16296),
            .in2(_gnd_net_),
            .in3(N__15971),
            .lcout(data_in_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i125_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i125_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i125_LC_5_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i125_LC_5_19_4  (
            .in0(N__16305),
            .in1(N__29646),
            .in2(_gnd_net_),
            .in3(N__16328),
            .lcout(data_in_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i133_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i133_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i133_LC_5_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i133_LC_5_19_5  (
            .in0(N__29643),
            .in1(N__16317),
            .in2(_gnd_net_),
            .in3(N__16304),
            .lcout(data_in_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i144_LC_5_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i144_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i144_LC_5_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i144_LC_5_19_6  (
            .in0(N__29648),
            .in1(N__20226),
            .in2(_gnd_net_),
            .in3(N__16295),
            .lcout(data_in_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i149_LC_5_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i149_LC_5_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i149_LC_5_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i149_LC_5_19_7  (
            .in0(N__29644),
            .in1(N__16287),
            .in2(_gnd_net_),
            .in3(N__16274),
            .lcout(data_in_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_5_21_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_5_21_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i22_LC_5_21_0  (
            .in0(N__16544),
            .in1(N__29795),
            .in2(_gnd_net_),
            .in3(N__16254),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i47_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i47_LC_5_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i47_LC_5_21_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i47_LC_5_21_1  (
            .in0(N__16596),
            .in1(_gnd_net_),
            .in2(N__29965),
            .in3(N__16219),
            .lcout(data_in_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i39_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i39_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i39_LC_5_21_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i39_LC_5_21_2  (
            .in0(N__16220),
            .in1(N__29796),
            .in2(_gnd_net_),
            .in3(N__16195),
            .lcout(data_in_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_5_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_5_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i29_LC_5_21_3  (
            .in0(N__29793),
            .in1(N__16907),
            .in2(_gnd_net_),
            .in3(N__18578),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i55_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i55_LC_5_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i55_LC_5_21_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i55_LC_5_21_4  (
            .in0(N__16562),
            .in1(N__29800),
            .in2(_gnd_net_),
            .in3(N__16595),
            .lcout(data_in_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_54_i1_3_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_54_i1_3_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_54_i1_3_lut_LC_5_21_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_54_i1_3_lut_LC_5_21_5  (
            .in0(N__16594),
            .in1(N__20879),
            .in2(_gnd_net_),
            .in3(N__23542),
            .lcout(n1889),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i63_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i63_LC_5_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i63_LC_5_21_6 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \c0.data_in_0___i63_LC_5_21_6  (
            .in0(N__16584),
            .in1(N__29801),
            .in2(N__16566),
            .in3(_gnd_net_),
            .lcout(data_in_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_5_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i30_LC_5_21_7  (
            .in0(N__29794),
            .in1(N__18289),
            .in2(_gnd_net_),
            .in3(N__16543),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i31_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i31_LC_5_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i31_LC_5_22_0 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \c0.data_in_frame_0___i31_LC_5_22_0  (
            .in0(N__16461),
            .in1(N__23553),
            .in2(N__16524),
            .in3(N__19119),
            .lcout(\c0.data_in_field_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_690_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_690_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_690_LC_5_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_690_LC_5_22_1  (
            .in0(N__22672),
            .in1(N__16616),
            .in2(N__16411),
            .in3(N__28042),
            .lcout(\c0.n8843 ),
            .ltout(\c0.n8843_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_621_LC_5_22_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_621_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_621_LC_5_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_621_LC_5_22_2  (
            .in0(N__18743),
            .in1(N__18677),
            .in2(N__16503),
            .in3(N__16489),
            .lcout(\c0.n4151 ),
            .ltout(\c0.n4151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_623_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_623_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_623_LC_5_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_623_LC_5_22_3  (
            .in0(N__21430),
            .in1(N__27989),
            .in2(N__16464),
            .in3(N__16459),
            .lcout(\c0.n8852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7945_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7945_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7945_LC_5_22_4 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7945_LC_5_22_4  (
            .in0(N__16460),
            .in1(N__32013),
            .in2(N__33032),
            .in3(N__16443),
            .lcout(),
            .ltout(\c0.n9638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9638_bdd_4_lut_LC_5_22_5 .C_ON=1'b0;
    defparam \c0.n9638_bdd_4_lut_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9638_bdd_4_lut_LC_5_22_5 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9638_bdd_4_lut_LC_5_22_5  (
            .in0(N__16404),
            .in1(N__32955),
            .in2(N__16383),
            .in3(N__16380),
            .lcout(\c0.n9132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i17_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i17_LC_5_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i17_LC_5_22_6 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \c0.data_in_frame_0___i17_LC_5_22_6  (
            .in0(N__28043),
            .in1(N__23554),
            .in2(N__16884),
            .in3(N__19118),
            .lcout(\c0.data_in_field_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i29_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i29_LC_5_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i29_LC_5_22_7 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \c0.data_in_frame_0___i29_LC_5_22_7  (
            .in0(N__19117),
            .in1(N__18577),
            .in2(N__23565),
            .in3(N__18744),
            .lcout(\c0.data_in_field_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7910_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7910_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7910_LC_5_23_0 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7910_LC_5_23_0  (
            .in0(N__32957),
            .in1(N__32012),
            .in2(N__21735),
            .in3(N__22147),
            .lcout(\c0.n9602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7840_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7840_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7840_LC_5_23_1 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7840_LC_5_23_1  (
            .in0(N__32011),
            .in1(N__16848),
            .in2(N__16817),
            .in3(N__32956),
            .lcout(\c0.n9512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \c0.data_in_frame_0___i18_LC_5_23_2  (
            .in0(N__16764),
            .in1(N__23501),
            .in2(N__19130),
            .in3(N__17304),
            .lcout(\c0.data_in_field_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_616_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_616_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_616_LC_5_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_616_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(N__16945),
            .in2(_gnd_net_),
            .in3(N__16614),
            .lcout(\c0.n4492 ),
            .ltout(\c0.n4492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_617_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_617_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_617_LC_5_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_617_LC_5_23_4  (
            .in0(N__16716),
            .in1(N__16698),
            .in2(N__16686),
            .in3(N__22991),
            .lcout(\c0.n8948 ),
            .ltout(\c0.n8948_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_525_LC_5_23_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_525_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_525_LC_5_23_5 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i4_4_lut_adj_525_LC_5_23_5  (
            .in0(N__22146),
            .in1(N__25019),
            .in2(N__16683),
            .in3(N__16676),
            .lcout(\c0.n19_adj_1602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i2_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i2_LC_5_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i2_LC_5_23_6 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \c0.data_in_frame_0___i2_LC_5_23_6  (
            .in0(N__16615),
            .in1(N__23502),
            .in2(N__19131),
            .in3(N__16650),
            .lcout(\c0.data_in_field_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i16_LC_5_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i16_LC_5_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i16_LC_5_23_7 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \c0.data_in_frame_0___i16_LC_5_23_7  (
            .in0(N__16980),
            .in1(N__16946),
            .in2(N__23552),
            .in3(N__19074),
            .lcout(\c0.data_in_field_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i43_LC_5_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i43_LC_5_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i43_LC_5_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0___i43_LC_5_24_0  (
            .in0(N__19056),
            .in1(N__22923),
            .in2(_gnd_net_),
            .in3(N__18676),
            .lcout(data_in_field_42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_48_i1_3_lut_LC_5_24_1 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_48_i1_3_lut_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_48_i1_3_lut_LC_5_24_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.mux_358_Mux_48_i1_3_lut_LC_5_24_1  (
            .in0(N__23506),
            .in1(_gnd_net_),
            .in2(N__20561),
            .in3(N__24128),
            .lcout(),
            .ltout(n1895_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i49_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i49_LC_5_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i49_LC_5_24_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_in_frame_0___i49_LC_5_24_2  (
            .in0(N__19058),
            .in1(_gnd_net_),
            .in2(N__16932),
            .in3(N__19213),
            .lcout(data_in_field_48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i55_LC_5_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i55_LC_5_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i55_LC_5_24_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i55_LC_5_24_3  (
            .in0(N__16929),
            .in1(N__24437),
            .in2(_gnd_net_),
            .in3(N__19061),
            .lcout(data_in_field_54),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i47_LC_5_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i47_LC_5_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i47_LC_5_24_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0___i47_LC_5_24_4  (
            .in0(N__19057),
            .in1(N__16920),
            .in2(_gnd_net_),
            .in3(N__22671),
            .lcout(data_in_field_46),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i37_LC_5_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i37_LC_5_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i37_LC_5_24_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.data_in_frame_0___i37_LC_5_24_5  (
            .in0(N__23507),
            .in1(N__16908),
            .in2(N__22804),
            .in3(N__19059),
            .lcout(data_in_field_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i41_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i41_LC_5_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i41_LC_5_24_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0___i41_LC_5_24_6  (
            .in0(N__19055),
            .in1(N__20643),
            .in2(_gnd_net_),
            .in3(N__18641),
            .lcout(data_in_field_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i51_LC_5_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i51_LC_5_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i51_LC_5_24_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i51_LC_5_24_7  (
            .in0(N__23202),
            .in1(N__26814),
            .in2(_gnd_net_),
            .in3(N__19060),
            .lcout(data_in_field_50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7830_LC_5_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7830_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7830_LC_5_25_0 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7830_LC_5_25_0  (
            .in0(N__32883),
            .in1(N__26816),
            .in2(N__32035),
            .in3(N__24033),
            .lcout(),
            .ltout(\c0.n9506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9506_bdd_4_lut_LC_5_25_1 .C_ON=1'b0;
    defparam \c0.n9506_bdd_4_lut_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9506_bdd_4_lut_LC_5_25_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9506_bdd_4_lut_LC_5_25_1  (
            .in0(N__32890),
            .in1(N__18675),
            .in2(N__17073),
            .in3(N__17070),
            .lcout(\c0.n9195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_516_LC_5_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_516_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_516_LC_5_25_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_516_LC_5_25_2  (
            .in0(N__22779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17664),
            .lcout(),
            .ltout(\c0.n4_adj_1592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_522_LC_5_25_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_522_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_522_LC_5_25_3 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i6_4_lut_adj_522_LC_5_25_3  (
            .in0(N__26815),
            .in1(N__27119),
            .in2(N__17034),
            .in3(N__17031),
            .lcout(\c0.n21_adj_1599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i81_LC_5_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i81_LC_5_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i81_LC_5_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i81_LC_5_25_4  (
            .in0(N__24129),
            .in1(N__27930),
            .in2(_gnd_net_),
            .in3(N__28673),
            .lcout(data_in_field_80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_5_25_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_5_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_LC_5_25_5  (
            .in0(N__17136),
            .in1(N__17013),
            .in2(N__16995),
            .in3(N__16986),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i57_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i57_LC_5_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i57_LC_5_26_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i57_LC_5_26_0  (
            .in0(N__20921),
            .in1(_gnd_net_),
            .in2(N__28749),
            .in3(N__24213),
            .lcout(data_in_field_56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i140_LC_5_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i140_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i140_LC_5_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i140_LC_5_26_1  (
            .in0(N__26739),
            .in1(N__17394),
            .in2(_gnd_net_),
            .in3(N__28578),
            .lcout(data_in_field_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i95_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i95_LC_5_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i95_LC_5_26_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i95_LC_5_26_2  (
            .in0(N__19365),
            .in1(_gnd_net_),
            .in2(N__28751),
            .in3(N__22523),
            .lcout(data_in_field_94),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_512_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_512_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_512_LC_5_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_512_LC_5_26_3  (
            .in0(N__23012),
            .in1(N__17235),
            .in2(N__17217),
            .in3(N__17205),
            .lcout(),
            .ltout(\c0.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_5_26_4 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_5_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_LC_5_26_4  (
            .in0(_gnd_net_),
            .in1(N__17190),
            .in2(N__17178),
            .in3(N__17175),
            .lcout(),
            .ltout(\c0.n8421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_529_LC_5_26_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_529_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_529_LC_5_26_5 .LUT_INIT=16'b1111111011111101;
    LogicCell40 \c0.i9_4_lut_adj_529_LC_5_26_5  (
            .in0(N__25250),
            .in1(N__17163),
            .in2(N__17157),
            .in3(N__17154),
            .lcout(\c0.n24_adj_1605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i78_LC_5_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i78_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i78_LC_5_26_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0___i78_LC_5_26_6  (
            .in0(N__22411),
            .in1(_gnd_net_),
            .in2(N__28750),
            .in3(N__21278),
            .lcout(data_in_field_77),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i93_LC_5_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i93_LC_5_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i93_LC_5_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i93_LC_5_26_7  (
            .in0(N__29108),
            .in1(N__24944),
            .in2(_gnd_net_),
            .in3(N__28585),
            .lcout(data_in_field_92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i76_LC_5_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i76_LC_5_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i76_LC_5_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i76_LC_5_27_0  (
            .in0(N__19552),
            .in1(N__17126),
            .in2(_gnd_net_),
            .in3(N__28665),
            .lcout(data_in_field_75),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i79_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i79_LC_5_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i79_LC_5_27_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i79_LC_5_27_1  (
            .in0(_gnd_net_),
            .in1(N__22304),
            .in2(N__28854),
            .in3(N__26381),
            .lcout(data_in_field_78),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i94_LC_5_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i94_LC_5_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i94_LC_5_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i94_LC_5_27_2  (
            .in0(N__21464),
            .in1(N__22000),
            .in2(_gnd_net_),
            .in3(N__28672),
            .lcout(data_in_field_93),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i68_LC_5_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i68_LC_5_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i68_LC_5_27_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i68_LC_5_27_3  (
            .in0(N__21156),
            .in1(_gnd_net_),
            .in2(N__28853),
            .in3(N__17097),
            .lcout(data_in_field_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i120_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i120_LC_5_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i120_LC_5_27_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i120_LC_5_27_4  (
            .in0(N__19722),
            .in1(N__25745),
            .in2(_gnd_net_),
            .in3(N__28658),
            .lcout(data_in_field_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i63_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i63_LC_5_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i63_LC_5_27_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i63_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(N__19354),
            .in2(N__28852),
            .in3(N__22715),
            .lcout(data_in_field_62),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_647_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_647_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_647_LC_5_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_647_LC_5_27_6  (
            .in0(N__17340),
            .in1(N__17331),
            .in2(N__27621),
            .in3(N__19781),
            .lcout(\c0.n8939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i92_LC_5_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i92_LC_5_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i92_LC_5_27_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i92_LC_5_27_7  (
            .in0(N__26721),
            .in1(_gnd_net_),
            .in2(N__28855),
            .in3(N__21873),
            .lcout(data_in_field_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_727_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_727_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_727_LC_5_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_727_LC_5_28_0  (
            .in0(N__25220),
            .in1(N__21225),
            .in2(_gnd_net_),
            .in3(N__17703),
            .lcout(\c0.n8992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_5_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_5_28_1  (
            .in0(N__22562),
            .in1(N__21807),
            .in2(N__17325),
            .in3(N__17311),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i86_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i86_LC_5_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i86_LC_5_28_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i86_LC_5_28_2  (
            .in0(N__19676),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__28885),
            .lcout(data_in_field_85),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i61_LC_5_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i61_LC_5_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i61_LC_5_28_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i61_LC_5_28_3  (
            .in0(_gnd_net_),
            .in1(N__29097),
            .in2(N__29011),
            .in3(N__21774),
            .lcout(data_in_field_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i142_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i142_LC_5_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i142_LC_5_28_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i142_LC_5_28_4  (
            .in0(N__21459),
            .in1(N__19920),
            .in2(_gnd_net_),
            .in3(N__28881),
            .lcout(data_in_field_141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_622_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_622_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_622_LC_5_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_622_LC_5_28_5  (
            .in0(N__23851),
            .in1(N__20739),
            .in2(N__21750),
            .in3(N__17261),
            .lcout(\c0.n19_adj_1643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i127_LC_5_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i127_LC_5_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i127_LC_5_28_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i127_LC_5_28_6  (
            .in0(N__19353),
            .in1(N__22563),
            .in2(_gnd_net_),
            .in3(N__28877),
            .lcout(data_in_field_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i138_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i138_LC_5_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i138_LC_5_28_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0___i138_LC_5_28_7  (
            .in0(N__17704),
            .in1(_gnd_net_),
            .in2(N__29010),
            .in3(N__21661),
            .lcout(data_in_field_137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_644_LC_5_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_644_LC_5_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_644_LC_5_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_644_LC_5_29_0  (
            .in0(N__17602),
            .in1(N__31419),
            .in2(N__17550),
            .in3(N__21623),
            .lcout(\c0.n22_adj_1617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i73_LC_5_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i73_LC_5_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i73_LC_5_29_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i73_LC_5_29_1  (
            .in0(_gnd_net_),
            .in1(N__20671),
            .in2(N__29014),
            .in3(N__27886),
            .lcout(data_in_field_72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i137_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i137_LC_5_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i137_LC_5_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i137_LC_5_29_2  (
            .in0(N__20916),
            .in1(N__26212),
            .in2(_gnd_net_),
            .in3(N__28892),
            .lcout(data_in_field_136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_604_LC_5_29_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_604_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_604_LC_5_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_604_LC_5_29_3  (
            .in0(N__17643),
            .in1(N__17885),
            .in2(N__20749),
            .in3(N__17510),
            .lcout(\c0.n4302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i80_LC_5_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i80_LC_5_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i80_LC_5_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i80_LC_5_29_4  (
            .in0(N__19501),
            .in1(N__17436),
            .in2(_gnd_net_),
            .in3(N__28896),
            .lcout(data_in_field_79),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_726_LC_5_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_726_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_726_LC_5_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_726_LC_5_29_5  (
            .in0(N__23849),
            .in1(N__27784),
            .in2(N__17402),
            .in3(N__17357),
            .lcout(\c0.n8782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_709_LC_5_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_709_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_709_LC_5_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_709_LC_5_29_6  (
            .in0(N__27785),
            .in1(N__23850),
            .in2(_gnd_net_),
            .in3(N__22516),
            .lcout(\c0.n8977 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i112_LC_5_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i112_LC_5_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i112_LC_5_29_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i112_LC_5_29_7  (
            .in0(_gnd_net_),
            .in1(N__19500),
            .in2(N__29013),
            .in3(N__17755),
            .lcout(data_in_field_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_5_30_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_5_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_5_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_718_LC_5_30_0  (
            .in0(N__25334),
            .in1(N__25219),
            .in2(N__19782),
            .in3(N__22327),
            .lcout(\c0.n4525 ),
            .ltout(\c0.n4525_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_557_LC_5_30_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_557_LC_5_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_557_LC_5_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_557_LC_5_30_1  (
            .in0(N__19677),
            .in1(N__17913),
            .in2(N__17736),
            .in3(N__22570),
            .lcout(\c0.n8924 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_589_LC_5_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_589_LC_5_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_589_LC_5_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_589_LC_5_30_2  (
            .in0(_gnd_net_),
            .in1(N__17733),
            .in2(_gnd_net_),
            .in3(N__17705),
            .lcout(\c0.n8874 ),
            .ltout(\c0.n8874_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_560_LC_5_30_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_560_LC_5_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_560_LC_5_30_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_560_LC_5_30_3  (
            .in0(N__22245),
            .in1(N__27137),
            .in2(N__17682),
            .in3(N__25722),
            .lcout(\c0.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_602_LC_5_30_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_602_LC_5_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_602_LC_5_30_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_602_LC_5_30_4  (
            .in0(_gnd_net_),
            .in1(N__24390),
            .in2(_gnd_net_),
            .in3(N__17678),
            .lcout(\c0.n6_adj_1636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i134_LC_5_30_5  (
            .in0(N__19304),
            .in1(N__32586),
            .in2(_gnd_net_),
            .in3(N__29057),
            .lcout(data_in_field_133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_701_LC_5_30_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_701_LC_5_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_701_LC_5_30_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_701_LC_5_30_6  (
            .in0(N__19475),
            .in1(N__25277),
            .in2(_gnd_net_),
            .in3(N__27045),
            .lcout(\c0.n8989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i70_LC_5_30_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i70_LC_5_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i70_LC_5_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i70_LC_5_30_7  (
            .in0(N__24391),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__29058),
            .lcout(data_in_field_69),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_528_LC_5_31_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_528_LC_5_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_528_LC_5_31_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_528_LC_5_31_0  (
            .in0(_gnd_net_),
            .in1(N__17912),
            .in2(_gnd_net_),
            .in3(N__21928),
            .lcout(),
            .ltout(\c0.n6_adj_1604_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_530_LC_5_31_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_530_LC_5_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_530_LC_5_31_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_530_LC_5_31_1  (
            .in0(N__24047),
            .in1(N__22729),
            .in2(N__18012),
            .in3(N__27429),
            .lcout(\c0.n8983 ),
            .ltout(\c0.n8983_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_5_31_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_5_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_5_31_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_5_31_2  (
            .in0(N__17997),
            .in1(N__17985),
            .in2(N__17976),
            .in3(N__17973),
            .lcout(\c0.n26_adj_1606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_556_LC_5_31_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_556_LC_5_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_556_LC_5_31_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_556_LC_5_31_3  (
            .in0(N__17954),
            .in1(N__25139),
            .in2(N__26462),
            .in3(N__32121),
            .lcout(\c0.n4203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_532_LC_5_31_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_532_LC_5_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_532_LC_5_31_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_532_LC_5_31_4  (
            .in0(N__17898),
            .in1(N__26115),
            .in2(N__20583),
            .in3(N__17886),
            .lcout(),
            .ltout(\c0.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i164_LC_5_31_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i164_LC_5_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i164_LC_5_31_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i164_LC_5_31_5  (
            .in0(N__17874),
            .in1(N__17862),
            .in2(N__17856),
            .in3(N__17853),
            .lcout(\c0.data_in_frame_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(N__29021),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_561_LC_5_32_0 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_561_LC_5_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_561_LC_5_32_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_561_LC_5_32_0  (
            .in0(N__24365),
            .in1(N__17828),
            .in2(N__17805),
            .in3(N__17790),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1509_2_lut_LC_5_32_1 .C_ON=1'b0;
    defparam \c0.i1509_2_lut_LC_5_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1509_2_lut_LC_5_32_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1509_2_lut_LC_5_32_1  (
            .in0(_gnd_net_),
            .in1(N__32045),
            .in2(_gnd_net_),
            .in3(N__33138),
            .lcout(\c0.n3056 ),
            .ltout(\c0.n3056_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_5_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_5_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_5_32_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_5_32_2  (
            .in0(N__17778),
            .in1(N__18036),
            .in2(N__18114),
            .in3(N__31263),
            .lcout(\c0.n22_adj_1676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i160_LC_5_32_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i160_LC_5_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i160_LC_5_32_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i160_LC_5_32_3  (
            .in0(N__24999),
            .in1(N__18099),
            .in2(N__18093),
            .in3(N__18081),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35398),
            .ce(N__29072),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7960_LC_5_32_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7960_LC_5_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7960_LC_5_32_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7960_LC_5_32_4  (
            .in0(N__25213),
            .in1(N__33148),
            .in2(N__18075),
            .in3(N__32046),
            .lcout(),
            .ltout(\c0.n9662_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9662_bdd_4_lut_LC_5_32_5 .C_ON=1'b0;
    defparam \c0.n9662_bdd_4_lut_LC_5_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9662_bdd_4_lut_LC_5_32_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9662_bdd_4_lut_LC_5_32_5  (
            .in0(N__33149),
            .in1(N__18066),
            .in2(N__18039),
            .in3(N__21555),
            .lcout(\c0.n9665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i84_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i84_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i84_LC_6_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i84_LC_6_18_0  (
            .in0(N__29975),
            .in1(N__20070),
            .in2(_gnd_net_),
            .in3(N__18140),
            .lcout(data_in_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i110_LC_6_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i110_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i110_LC_6_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i110_LC_6_18_1  (
            .in0(N__29966),
            .in1(N__19973),
            .in2(_gnd_net_),
            .in3(N__19953),
            .lcout(data_in_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i100_LC_6_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i100_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i100_LC_6_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i100_LC_6_18_2  (
            .in0(N__18030),
            .in1(N__29969),
            .in2(_gnd_net_),
            .in3(N__20081),
            .lcout(data_in_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i108_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i108_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i108_LC_6_18_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i108_LC_6_18_3  (
            .in0(N__18021),
            .in1(N__29976),
            .in2(_gnd_net_),
            .in3(N__18029),
            .lcout(data_in_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i116_LC_6_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i116_LC_6_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i116_LC_6_18_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i116_LC_6_18_4  (
            .in0(N__18219),
            .in1(N__29970),
            .in2(_gnd_net_),
            .in3(N__18020),
            .lcout(data_in_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i124_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i124_LC_6_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i124_LC_6_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i124_LC_6_18_5  (
            .in0(N__29967),
            .in1(N__18231),
            .in2(_gnd_net_),
            .in3(N__18218),
            .lcout(data_in_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i140_LC_6_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i140_LC_6_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i140_LC_6_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i140_LC_6_18_7  (
            .in0(N__29968),
            .in1(N__18198),
            .in2(_gnd_net_),
            .in3(N__18209),
            .lcout(data_in_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i148_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i148_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i148_LC_6_19_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i148_LC_6_19_0  (
            .in0(N__18186),
            .in1(N__29652),
            .in2(_gnd_net_),
            .in3(N__18197),
            .lcout(data_in_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i156_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i156_LC_6_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i156_LC_6_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i156_LC_6_19_1  (
            .in0(N__18177),
            .in1(N__29654),
            .in2(_gnd_net_),
            .in3(N__18185),
            .lcout(data_in_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i164_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i164_LC_6_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i164_LC_6_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i164_LC_6_19_2  (
            .in0(N__29656),
            .in1(N__20271),
            .in2(_gnd_net_),
            .in3(N__18176),
            .lcout(data_in_20_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i150_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i150_LC_6_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i150_LC_6_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i150_LC_6_19_3  (
            .in0(N__18168),
            .in1(N__29653),
            .in2(_gnd_net_),
            .in3(N__20165),
            .lcout(data_in_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i158_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i158_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i158_LC_6_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i158_LC_6_19_4  (
            .in0(N__29655),
            .in1(N__18324),
            .in2(_gnd_net_),
            .in3(N__18167),
            .lcout(data_in_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i143_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i143_LC_6_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i143_LC_6_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i143_LC_6_19_5  (
            .in0(N__29651),
            .in1(N__20145),
            .in2(_gnd_net_),
            .in3(N__18155),
            .lcout(data_in_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_31_i4_2_lut_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.rx.equal_31_i4_2_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_31_i4_2_lut_LC_6_20_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.equal_31_i4_2_lut_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__27552),
            .in2(_gnd_net_),
            .in3(N__25874),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i76_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i76_LC_6_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i76_LC_6_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i76_LC_6_20_6  (
            .in0(N__29924),
            .in1(N__18125),
            .in2(_gnd_net_),
            .in3(N__18144),
            .lcout(data_in_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i166_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i166_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i166_LC_6_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i166_LC_6_20_7  (
            .in0(N__29923),
            .in1(N__20351),
            .in2(_gnd_net_),
            .in3(N__18323),
            .lcout(data_in_20_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_45_i1_3_lut_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_45_i1_3_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_45_i1_3_lut_LC_6_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_358_Mux_45_i1_3_lut_LC_6_21_0  (
            .in0(N__21274),
            .in1(N__18310),
            .in2(_gnd_net_),
            .in3(N__23543),
            .lcout(n1898),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i46_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i46_LC_6_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i46_LC_6_21_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i46_LC_6_21_1  (
            .in0(N__18311),
            .in1(N__29803),
            .in2(_gnd_net_),
            .in3(N__18270),
            .lcout(data_in_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i38_LC_6_21_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i38_LC_6_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i38_LC_6_21_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i38_LC_6_21_2  (
            .in0(N__29802),
            .in1(N__18312),
            .in2(_gnd_net_),
            .in3(N__18290),
            .lcout(data_in_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i54_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i54_LC_6_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i54_LC_6_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i54_LC_6_21_3  (
            .in0(N__29838),
            .in1(N__18258),
            .in2(_gnd_net_),
            .in3(N__18269),
            .lcout(data_in_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_53_i1_3_lut_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_53_i1_3_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_53_i1_3_lut_LC_6_21_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_53_i1_3_lut_LC_6_21_4  (
            .in0(N__18268),
            .in1(N__19887),
            .in2(_gnd_net_),
            .in3(N__23544),
            .lcout(n1890),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i62_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i62_LC_6_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i62_LC_6_21_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i62_LC_6_21_5  (
            .in0(N__18249),
            .in1(N__29804),
            .in2(_gnd_net_),
            .in3(N__18257),
            .lcout(data_in_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i70_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i70_LC_6_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i70_LC_6_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i70_LC_6_21_6  (
            .in0(N__18240),
            .in1(N__29837),
            .in2(_gnd_net_),
            .in3(N__18248),
            .lcout(data_in_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i78_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i78_LC_6_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i78_LC_6_21_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i78_LC_6_21_7  (
            .in0(N__29839),
            .in1(N__18239),
            .in2(_gnd_net_),
            .in3(N__20001),
            .lcout(data_in_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i113_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i113_LC_6_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i113_LC_6_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i113_LC_6_22_0  (
            .in0(N__18393),
            .in1(N__29983),
            .in2(_gnd_net_),
            .in3(N__18404),
            .lcout(data_in_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i121_LC_6_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i121_LC_6_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i121_LC_6_22_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i121_LC_6_22_1  (
            .in0(N__29980),
            .in1(N__18354),
            .in2(_gnd_net_),
            .in3(N__18392),
            .lcout(data_in_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i135_LC_6_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i135_LC_6_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i135_LC_6_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i135_LC_6_22_2  (
            .in0(N__24657),
            .in1(N__25784),
            .in2(_gnd_net_),
            .in3(N__29012),
            .lcout(data_in_field_134),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_6_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_6_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_6_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i19_LC_6_22_3  (
            .in0(N__29982),
            .in1(N__18544),
            .in2(_gnd_net_),
            .in3(N__18375),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i153_LC_6_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i153_LC_6_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i153_LC_6_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i153_LC_6_22_4  (
            .in0(N__18341),
            .in1(N__29984),
            .in2(_gnd_net_),
            .in3(N__29147),
            .lcout(data_in_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i129_LC_6_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i129_LC_6_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i129_LC_6_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i129_LC_6_22_5  (
            .in0(N__29981),
            .in1(N__18483),
            .in2(_gnd_net_),
            .in3(N__18353),
            .lcout(data_in_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i161_LC_6_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i161_LC_6_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i161_LC_6_22_6 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \c0.data_in_0___i161_LC_6_22_6  (
            .in0(N__20247),
            .in1(N__29985),
            .in2(N__18345),
            .in3(_gnd_net_),
            .lcout(data_in_20_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i46_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i46_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i46_LC_6_23_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i46_LC_6_23_0  (
            .in0(N__18333),
            .in1(N__18850),
            .in2(_gnd_net_),
            .in3(N__19148),
            .lcout(data_in_field_45),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8029_LC_6_23_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8029_LC_6_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8029_LC_6_23_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_8029_LC_6_23_1  (
            .in0(N__31910),
            .in1(N__32871),
            .in2(N__19215),
            .in3(N__24223),
            .lcout(),
            .ltout(\c0.n9746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9746_bdd_4_lut_LC_6_23_2 .C_ON=1'b0;
    defparam \c0.n9746_bdd_4_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.n9746_bdd_4_lut_LC_6_23_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9746_bdd_4_lut_LC_6_23_2  (
            .in0(N__18635),
            .in1(N__32872),
            .in2(N__18720),
            .in3(N__18717),
            .lcout(\c0.n9228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_686_LC_6_23_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_686_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_686_LC_6_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_686_LC_6_23_3  (
            .in0(N__18801),
            .in1(N__18668),
            .in2(_gnd_net_),
            .in3(N__18634),
            .lcout(\c0.n4208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_6_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_6_23_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i21_LC_6_23_4  (
            .in0(N__18582),
            .in1(N__18507),
            .in2(_gnd_net_),
            .in3(N__29873),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_6_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i27_LC_6_23_5  (
            .in0(N__29871),
            .in1(N__26978),
            .in2(_gnd_net_),
            .in3(N__18543),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_6_23_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_6_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_6_23_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i13_LC_6_23_6  (
            .in0(N__19181),
            .in1(N__18508),
            .in2(_gnd_net_),
            .in3(N__29872),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i137_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i137_LC_6_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i137_LC_6_23_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i137_LC_6_23_7  (
            .in0(N__29870),
            .in1(N__29136),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(data_in_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_689_LC_6_24_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_689_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_689_LC_6_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_689_LC_6_24_0  (
            .in0(N__33303),
            .in1(N__25034),
            .in2(N__26541),
            .in3(N__27926),
            .lcout(\c0.n8960 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_6_24_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i5_LC_6_24_1  (
            .in0(N__30032),
            .in1(N__18439),
            .in2(_gnd_net_),
            .in3(N__19180),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i54_LC_6_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i54_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i54_LC_6_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i54_LC_6_24_2  (
            .in0(N__22151),
            .in1(N__18420),
            .in2(_gnd_net_),
            .in3(N__19113),
            .lcout(data_in_field_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i131_LC_6_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i131_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i131_LC_6_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i131_LC_6_24_3  (
            .in0(N__23714),
            .in1(N__26532),
            .in2(_gnd_net_),
            .in3(N__28752),
            .lcout(data_in_field_130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i13_LC_6_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i13_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i13_LC_6_24_4 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \c0.data_in_frame_0___i13_LC_6_24_4  (
            .in0(N__19179),
            .in1(N__23508),
            .in2(N__18812),
            .in3(N__19112),
            .lcout(\c0.data_in_field_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9602_bdd_4_lut_LC_6_24_5 .C_ON=1'b0;
    defparam \c0.n9602_bdd_4_lut_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9602_bdd_4_lut_LC_6_24_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9602_bdd_4_lut_LC_6_24_5  (
            .in0(N__32789),
            .in1(N__18849),
            .in2(N__18822),
            .in3(N__25613),
            .lcout(\c0.n9150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_586_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_586_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_586_LC_6_24_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_586_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(N__19206),
            .in2(_gnd_net_),
            .in3(N__18802),
            .lcout(\c0.n9019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_665_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_665_LC_6_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_665_LC_6_24_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_665_LC_6_24_7  (
            .in0(_gnd_net_),
            .in1(N__18757),
            .in2(_gnd_net_),
            .in3(N__22208),
            .lcout(\c0.n8813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i59_LC_6_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i59_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i59_LC_6_25_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i59_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__23944),
            .in2(N__28748),
            .in3(N__24040),
            .lcout(data_in_field_58),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_551_LC_6_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_551_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_551_LC_6_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_551_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__26484),
            .in2(_gnd_net_),
            .in3(N__26813),
            .lcout(\c0.n8828 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i150_LC_6_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i150_LC_6_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i150_LC_6_25_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i150_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__19305),
            .in2(N__28747),
            .in3(N__19769),
            .lcout(data_in_field_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i139_LC_6_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i139_LC_6_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i139_LC_6_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i139_LC_6_25_3  (
            .in0(N__23943),
            .in1(N__26485),
            .in2(_gnd_net_),
            .in3(N__28567),
            .lcout(data_in_field_138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i125_LC_6_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i125_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i125_LC_6_25_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i125_LC_6_25_4  (
            .in0(_gnd_net_),
            .in1(N__29107),
            .in2(N__28745),
            .in3(N__24281),
            .lcout(data_in_field_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i109_LC_6_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i109_LC_6_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i109_LC_6_25_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i109_LC_6_25_5  (
            .in0(N__21506),
            .in1(N__24887),
            .in2(_gnd_net_),
            .in3(N__28563),
            .lcout(data_in_field_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i143_LC_6_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i143_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i143_LC_6_25_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i143_LC_6_25_6  (
            .in0(_gnd_net_),
            .in1(N__19361),
            .in2(N__28746),
            .in3(N__26441),
            .lcout(data_in_field_142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i65_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i65_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i65_LC_6_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i65_LC_6_25_7  (
            .in0(N__27843),
            .in1(N__25987),
            .in2(_gnd_net_),
            .in3(N__28577),
            .lcout(data_in_field_64),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam i7420_4_lut_LC_6_26_0.C_ON=1'b0;
    defparam i7420_4_lut_LC_6_26_0.SEQ_MODE=4'b0000;
    defparam i7420_4_lut_LC_6_26_0.LUT_INIT=16'b1111010001010000;
    LogicCell40 i7420_4_lut_LC_6_26_0 (
            .in0(N__30269),
            .in1(N__30296),
            .in2(N__30360),
            .in3(N__30323),
            .lcout(n9091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7421_4_lut_LC_6_26_1.C_ON=1'b0;
    defparam i7421_4_lut_LC_6_26_1.SEQ_MODE=4'b0000;
    defparam i7421_4_lut_LC_6_26_1.LUT_INIT=16'b1111111010001010;
    LogicCell40 i7421_4_lut_LC_6_26_1 (
            .in0(N__30297),
            .in1(N__30270),
            .in2(N__30327),
            .in3(N__30359),
            .lcout(),
            .ltout(n9092_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7422_3_lut_LC_6_26_2.C_ON=1'b0;
    defparam i7422_3_lut_LC_6_26_2.SEQ_MODE=4'b0000;
    defparam i7422_3_lut_LC_6_26_2.LUT_INIT=16'b0000111101010101;
    LogicCell40 i7422_3_lut_LC_6_26_2 (
            .in0(N__19251),
            .in1(_gnd_net_),
            .in2(N__19245),
            .in3(N__30243),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_6_26_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_6_26_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_6_26_3  (
            .in0(N__31086),
            .in1(N__27447),
            .in2(N__31032),
            .in3(N__30972),
            .lcout(r_SM_Main_2_adj_1734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35364),
            .ce(),
            .sr(N__19227));
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_6_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_6_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_699_LC_6_26_4  (
            .in0(N__26380),
            .in1(N__25480),
            .in2(_gnd_net_),
            .in3(N__19214),
            .lcout(\c0.n8883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_3_lut_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.i20_3_lut_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20_3_lut_LC_6_26_5 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \c0.i20_3_lut_LC_6_26_5  (
            .in0(N__23662),
            .in1(N__23401),
            .in2(_gnd_net_),
            .in3(N__20774),
            .lcout(\c0.n4897 ),
            .ltout(\c0.n4897_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3607_2_lut_3_lut_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.i3607_2_lut_3_lut_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3607_2_lut_3_lut_LC_6_26_6 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \c0.i3607_2_lut_3_lut_LC_6_26_6  (
            .in0(N__23402),
            .in1(_gnd_net_),
            .in2(N__19323),
            .in3(N__23663),
            .lcout(\c0.n5154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7744_3_lut_LC_6_26_7 .C_ON=1'b0;
    defparam \c0.i7744_3_lut_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7744_3_lut_LC_6_26_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i7744_3_lut_LC_6_26_7  (
            .in0(N__23661),
            .in1(N__23400),
            .in2(_gnd_net_),
            .in3(N__20775),
            .lcout(n4806),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i0_LC_6_27_0.C_ON=1'b1;
    defparam rand_data_422__i0_LC_6_27_0.SEQ_MODE=4'b1000;
    defparam rand_data_422__i0_LC_6_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i0_LC_6_27_0 (
            .in0(_gnd_net_),
            .in1(N__25976),
            .in2(_gnd_net_),
            .in3(N__19320),
            .lcout(rand_data_0),
            .ltout(),
            .carryin(bfn_6_27_0_),
            .carryout(n8155),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i1_LC_6_27_1.C_ON=1'b1;
    defparam rand_data_422__i1_LC_6_27_1.SEQ_MODE=4'b1000;
    defparam rand_data_422__i1_LC_6_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i1_LC_6_27_1 (
            .in0(_gnd_net_),
            .in1(N__21018),
            .in2(_gnd_net_),
            .in3(N__19317),
            .lcout(rand_data_1),
            .ltout(),
            .carryin(n8155),
            .carryout(n8156),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i2_LC_6_27_2.C_ON=1'b1;
    defparam rand_data_422__i2_LC_6_27_2.SEQ_MODE=4'b1000;
    defparam rand_data_422__i2_LC_6_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i2_LC_6_27_2 (
            .in0(_gnd_net_),
            .in1(N__23706),
            .in2(_gnd_net_),
            .in3(N__19314),
            .lcout(rand_data_2),
            .ltout(),
            .carryin(n8156),
            .carryout(n8157),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i3_LC_6_27_3.C_ON=1'b1;
    defparam rand_data_422__i3_LC_6_27_3.SEQ_MODE=4'b1000;
    defparam rand_data_422__i3_LC_6_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i3_LC_6_27_3 (
            .in0(_gnd_net_),
            .in1(N__21144),
            .in2(_gnd_net_),
            .in3(N__19311),
            .lcout(rand_data_3),
            .ltout(),
            .carryin(n8157),
            .carryout(n8158),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i4_LC_6_27_4.C_ON=1'b1;
    defparam rand_data_422__i4_LC_6_27_4.SEQ_MODE=4'b1000;
    defparam rand_data_422__i4_LC_6_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i4_LC_6_27_4 (
            .in0(_gnd_net_),
            .in1(N__21179),
            .in2(_gnd_net_),
            .in3(N__19308),
            .lcout(rand_data_4),
            .ltout(),
            .carryin(n8158),
            .carryout(n8159),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i5_LC_6_27_5.C_ON=1'b1;
    defparam rand_data_422__i5_LC_6_27_5.SEQ_MODE=4'b1000;
    defparam rand_data_422__i5_LC_6_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i5_LC_6_27_5 (
            .in0(_gnd_net_),
            .in1(N__19272),
            .in2(_gnd_net_),
            .in3(N__19257),
            .lcout(rand_data_5),
            .ltout(),
            .carryin(n8159),
            .carryout(n8160),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i6_LC_6_27_6.C_ON=1'b1;
    defparam rand_data_422__i6_LC_6_27_6.SEQ_MODE=4'b1000;
    defparam rand_data_422__i6_LC_6_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i6_LC_6_27_6 (
            .in0(_gnd_net_),
            .in1(N__24629),
            .in2(_gnd_net_),
            .in3(N__19254),
            .lcout(rand_data_6),
            .ltout(),
            .carryin(n8160),
            .carryout(n8161),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i7_LC_6_27_7.C_ON=1'b1;
    defparam rand_data_422__i7_LC_6_27_7.SEQ_MODE=4'b1000;
    defparam rand_data_422__i7_LC_6_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i7_LC_6_27_7 (
            .in0(_gnd_net_),
            .in1(N__21063),
            .in2(_gnd_net_),
            .in3(N__19386),
            .lcout(rand_data_7),
            .ltout(),
            .carryin(n8161),
            .carryout(n8162),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i8_LC_6_28_0.C_ON=1'b1;
    defparam rand_data_422__i8_LC_6_28_0.SEQ_MODE=4'b1000;
    defparam rand_data_422__i8_LC_6_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i8_LC_6_28_0 (
            .in0(_gnd_net_),
            .in1(N__20903),
            .in2(_gnd_net_),
            .in3(N__19383),
            .lcout(rand_data_8),
            .ltout(),
            .carryin(bfn_6_28_0_),
            .carryout(n8163),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i9_LC_6_28_1.C_ON=1'b1;
    defparam rand_data_422__i9_LC_6_28_1.SEQ_MODE=4'b1000;
    defparam rand_data_422__i9_LC_6_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i9_LC_6_28_1 (
            .in0(_gnd_net_),
            .in1(N__21650),
            .in2(_gnd_net_),
            .in3(N__19380),
            .lcout(rand_data_9),
            .ltout(),
            .carryin(n8163),
            .carryout(n8164),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i10_LC_6_28_2.C_ON=1'b1;
    defparam rand_data_422__i10_LC_6_28_2.SEQ_MODE=4'b1000;
    defparam rand_data_422__i10_LC_6_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i10_LC_6_28_2 (
            .in0(_gnd_net_),
            .in1(N__23932),
            .in2(_gnd_net_),
            .in3(N__19377),
            .lcout(rand_data_10),
            .ltout(),
            .carryin(n8164),
            .carryout(n8165),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i11_LC_6_28_3.C_ON=1'b1;
    defparam rand_data_422__i11_LC_6_28_3.SEQ_MODE=4'b1000;
    defparam rand_data_422__i11_LC_6_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i11_LC_6_28_3 (
            .in0(_gnd_net_),
            .in1(N__26717),
            .in2(_gnd_net_),
            .in3(N__19374),
            .lcout(rand_data_11),
            .ltout(),
            .carryin(n8165),
            .carryout(n8166),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i12_LC_6_28_4.C_ON=1'b1;
    defparam rand_data_422__i12_LC_6_28_4.SEQ_MODE=4'b1000;
    defparam rand_data_422__i12_LC_6_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i12_LC_6_28_4 (
            .in0(_gnd_net_),
            .in1(N__29096),
            .in2(_gnd_net_),
            .in3(N__19371),
            .lcout(rand_data_12),
            .ltout(),
            .carryin(n8166),
            .carryout(n8167),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i13_LC_6_28_5.C_ON=1'b1;
    defparam rand_data_422__i13_LC_6_28_5.SEQ_MODE=4'b1000;
    defparam rand_data_422__i13_LC_6_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i13_LC_6_28_5 (
            .in0(_gnd_net_),
            .in1(N__21458),
            .in2(_gnd_net_),
            .in3(N__19368),
            .lcout(rand_data_13),
            .ltout(),
            .carryin(n8167),
            .carryout(n8168),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i14_LC_6_28_6.C_ON=1'b1;
    defparam rand_data_422__i14_LC_6_28_6.SEQ_MODE=4'b1000;
    defparam rand_data_422__i14_LC_6_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i14_LC_6_28_6 (
            .in0(_gnd_net_),
            .in1(N__19352),
            .in2(_gnd_net_),
            .in3(N__19329),
            .lcout(rand_data_14),
            .ltout(),
            .carryin(n8168),
            .carryout(n8169),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i15_LC_6_28_7.C_ON=1'b1;
    defparam rand_data_422__i15_LC_6_28_7.SEQ_MODE=4'b1000;
    defparam rand_data_422__i15_LC_6_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i15_LC_6_28_7 (
            .in0(_gnd_net_),
            .in1(N__21576),
            .in2(_gnd_net_),
            .in3(N__19326),
            .lcout(rand_data_15),
            .ltout(),
            .carryin(n8169),
            .carryout(n8170),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i16_LC_6_29_0.C_ON=1'b1;
    defparam rand_data_422__i16_LC_6_29_0.SEQ_MODE=4'b1000;
    defparam rand_data_422__i16_LC_6_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i16_LC_6_29_0 (
            .in0(_gnd_net_),
            .in1(N__24106),
            .in2(_gnd_net_),
            .in3(N__19449),
            .lcout(rand_data_16),
            .ltout(),
            .carryin(bfn_6_29_0_),
            .carryout(n8171),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i17_LC_6_29_1.C_ON=1'b1;
    defparam rand_data_422__i17_LC_6_29_1.SEQ_MODE=4'b1000;
    defparam rand_data_422__i17_LC_6_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i17_LC_6_29_1 (
            .in0(_gnd_net_),
            .in1(N__19839),
            .in2(_gnd_net_),
            .in3(N__19446),
            .lcout(rand_data_17),
            .ltout(),
            .carryin(n8171),
            .carryout(n8172),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i18_LC_6_29_2.C_ON=1'b1;
    defparam rand_data_422__i18_LC_6_29_2.SEQ_MODE=4'b1000;
    defparam rand_data_422__i18_LC_6_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i18_LC_6_29_2 (
            .in0(_gnd_net_),
            .in1(N__26126),
            .in2(_gnd_net_),
            .in3(N__19443),
            .lcout(rand_data_18),
            .ltout(),
            .carryin(n8172),
            .carryout(n8173),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i19_LC_6_29_3.C_ON=1'b1;
    defparam rand_data_422__i19_LC_6_29_3.SEQ_MODE=4'b1000;
    defparam rand_data_422__i19_LC_6_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i19_LC_6_29_3 (
            .in0(_gnd_net_),
            .in1(N__19420),
            .in2(_gnd_net_),
            .in3(N__19404),
            .lcout(rand_data_19),
            .ltout(),
            .carryin(n8173),
            .carryout(n8174),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i20_LC_6_29_4.C_ON=1'b1;
    defparam rand_data_422__i20_LC_6_29_4.SEQ_MODE=4'b1000;
    defparam rand_data_422__i20_LC_6_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i20_LC_6_29_4 (
            .in0(_gnd_net_),
            .in1(N__24313),
            .in2(_gnd_net_),
            .in3(N__19401),
            .lcout(rand_data_20),
            .ltout(),
            .carryin(n8174),
            .carryout(n8175),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i21_LC_6_29_5.C_ON=1'b1;
    defparam rand_data_422__i21_LC_6_29_5.SEQ_MODE=4'b1000;
    defparam rand_data_422__i21_LC_6_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i21_LC_6_29_5 (
            .in0(_gnd_net_),
            .in1(N__19875),
            .in2(_gnd_net_),
            .in3(N__19398),
            .lcout(rand_data_21),
            .ltout(),
            .carryin(n8175),
            .carryout(n8176),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i22_LC_6_29_6.C_ON=1'b1;
    defparam rand_data_422__i22_LC_6_29_6.SEQ_MODE=4'b1000;
    defparam rand_data_422__i22_LC_6_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i22_LC_6_29_6 (
            .in0(_gnd_net_),
            .in1(N__20848),
            .in2(_gnd_net_),
            .in3(N__19395),
            .lcout(rand_data_22),
            .ltout(),
            .carryin(n8176),
            .carryout(n8177),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i23_LC_6_29_7.C_ON=1'b1;
    defparam rand_data_422__i23_LC_6_29_7.SEQ_MODE=4'b1000;
    defparam rand_data_422__i23_LC_6_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i23_LC_6_29_7 (
            .in0(_gnd_net_),
            .in1(N__19704),
            .in2(_gnd_net_),
            .in3(N__19392),
            .lcout(rand_data_23),
            .ltout(),
            .carryin(n8177),
            .carryout(n8178),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i24_LC_6_30_0.C_ON=1'b1;
    defparam rand_data_422__i24_LC_6_30_0.SEQ_MODE=4'b1000;
    defparam rand_data_422__i24_LC_6_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i24_LC_6_30_0 (
            .in0(_gnd_net_),
            .in1(N__20664),
            .in2(_gnd_net_),
            .in3(N__19389),
            .lcout(rand_data_24),
            .ltout(),
            .carryin(bfn_6_30_0_),
            .carryout(n8179),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i25_LC_6_30_1.C_ON=1'b1;
    defparam rand_data_422__i25_LC_6_30_1.SEQ_MODE=4'b1000;
    defparam rand_data_422__i25_LC_6_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i25_LC_6_30_1 (
            .in0(_gnd_net_),
            .in1(N__19588),
            .in2(_gnd_net_),
            .in3(N__19572),
            .lcout(rand_data_25),
            .ltout(),
            .carryin(n8179),
            .carryout(n8180),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i26_LC_6_30_2.C_ON=1'b1;
    defparam rand_data_422__i26_LC_6_30_2.SEQ_MODE=4'b1000;
    defparam rand_data_422__i26_LC_6_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i26_LC_6_30_2 (
            .in0(_gnd_net_),
            .in1(N__24070),
            .in2(_gnd_net_),
            .in3(N__19569),
            .lcout(rand_data_26),
            .ltout(),
            .carryin(n8180),
            .carryout(n8181),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i27_LC_6_30_3.C_ON=1'b1;
    defparam rand_data_422__i27_LC_6_30_3.SEQ_MODE=4'b1000;
    defparam rand_data_422__i27_LC_6_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i27_LC_6_30_3 (
            .in0(_gnd_net_),
            .in1(N__19539),
            .in2(_gnd_net_),
            .in3(N__19521),
            .lcout(rand_data_27),
            .ltout(),
            .carryin(n8181),
            .carryout(n8182),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i28_LC_6_30_4.C_ON=1'b1;
    defparam rand_data_422__i28_LC_6_30_4.SEQ_MODE=4'b1000;
    defparam rand_data_422__i28_LC_6_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i28_LC_6_30_4 (
            .in0(_gnd_net_),
            .in1(N__21486),
            .in2(_gnd_net_),
            .in3(N__19518),
            .lcout(rand_data_28),
            .ltout(),
            .carryin(n8182),
            .carryout(n8183),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i29_LC_6_30_5.C_ON=1'b1;
    defparam rand_data_422__i29_LC_6_30_5.SEQ_MODE=4'b1000;
    defparam rand_data_422__i29_LC_6_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i29_LC_6_30_5 (
            .in0(_gnd_net_),
            .in1(N__21258),
            .in2(_gnd_net_),
            .in3(N__19515),
            .lcout(rand_data_29),
            .ltout(),
            .carryin(n8183),
            .carryout(n8184),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i30_LC_6_30_6.C_ON=1'b1;
    defparam rand_data_422__i30_LC_6_30_6.SEQ_MODE=4'b1000;
    defparam rand_data_422__i30_LC_6_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i30_LC_6_30_6 (
            .in0(_gnd_net_),
            .in1(N__22284),
            .in2(_gnd_net_),
            .in3(N__19512),
            .lcout(rand_data_30),
            .ltout(),
            .carryin(n8184),
            .carryout(n8185),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_422__i31_LC_6_30_7.C_ON=1'b0;
    defparam rand_data_422__i31_LC_6_30_7.SEQ_MODE=4'b1000;
    defparam rand_data_422__i31_LC_6_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_422__i31_LC_6_30_7 (
            .in0(_gnd_net_),
            .in1(N__19502),
            .in2(_gnd_net_),
            .in3(N__19509),
            .lcout(rand_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8019_LC_6_31_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8019_LC_6_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8019_LC_6_31_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_8019_LC_6_31_0  (
            .in0(N__22326),
            .in1(N__27041),
            .in2(N__33014),
            .in3(N__32015),
            .lcout(),
            .ltout(\c0.n9734_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9734_bdd_4_lut_LC_6_31_1 .C_ON=1'b0;
    defparam \c0.n9734_bdd_4_lut_LC_6_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9734_bdd_4_lut_LC_6_31_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9734_bdd_4_lut_LC_6_31_1  (
            .in0(N__19479),
            .in1(N__32918),
            .in2(N__19452),
            .in3(N__27672),
            .lcout(\c0.n9234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_533_LC_6_31_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_533_LC_6_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_533_LC_6_31_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_533_LC_6_31_2  (
            .in0(N__19928),
            .in1(N__22058),
            .in2(_gnd_net_),
            .in3(N__19800),
            .lcout(\c0.n9013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i121_LC_6_31_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i121_LC_6_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i121_LC_6_31_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i121_LC_6_31_3  (
            .in0(N__22329),
            .in1(N__20920),
            .in2(_gnd_net_),
            .in3(N__29019),
            .lcout(data_in_field_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i118_LC_6_31_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i118_LC_6_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i118_LC_6_31_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i118_LC_6_31_4  (
            .in0(_gnd_net_),
            .in1(N__19886),
            .in2(N__29065),
            .in3(N__19631),
            .lcout(data_in_field_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i114_LC_6_31_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i114_LC_6_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i114_LC_6_31_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i114_LC_6_31_5  (
            .in0(N__19801),
            .in1(N__19852),
            .in2(_gnd_net_),
            .in3(N__29015),
            .lcout(data_in_field_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1290_2_lut_3_lut_LC_6_31_6 .C_ON=1'b0;
    defparam \c0.i1290_2_lut_3_lut_LC_6_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1290_2_lut_3_lut_LC_6_31_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1290_2_lut_3_lut_LC_6_31_6  (
            .in0(N__19771),
            .in1(N__25214),
            .in2(_gnd_net_),
            .in3(N__25338),
            .lcout(\c0.n1893_adj_1635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i88_LC_6_31_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i88_LC_6_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i88_LC_6_31_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i88_LC_6_31_7  (
            .in0(N__19715),
            .in1(N__21929),
            .in2(_gnd_net_),
            .in3(N__29020),
            .lcout(data_in_field_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7905_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7905_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7905_LC_6_32_0 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7905_LC_6_32_0  (
            .in0(N__19685),
            .in1(N__32052),
            .in2(N__33098),
            .in3(N__22022),
            .lcout(),
            .ltout(\c0.n9596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9596_bdd_4_lut_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.n9596_bdd_4_lut_LC_6_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9596_bdd_4_lut_LC_6_32_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n9596_bdd_4_lut_LC_6_32_1  (
            .in0(N__22418),
            .in1(N__24398),
            .in2(N__19638),
            .in3(N__33028),
            .lcout(\c0.n9153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7900_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7900_LC_6_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7900_LC_6_32_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7900_LC_6_32_2  (
            .in0(N__33029),
            .in1(N__19627),
            .in2(N__24559),
            .in3(N__32053),
            .lcout(),
            .ltout(\c0.n9590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9590_bdd_4_lut_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.n9590_bdd_4_lut_LC_6_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9590_bdd_4_lut_LC_6_32_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n9590_bdd_4_lut_LC_6_32_3  (
            .in0(N__24188),
            .in1(N__21232),
            .in2(N__20055),
            .in3(N__33030),
            .lcout(),
            .ltout(\c0.n9156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7915_LC_6_32_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7915_LC_6_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7915_LC_6_32_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7915_LC_6_32_4  (
            .in0(N__20052),
            .in1(N__31604),
            .in2(N__20046),
            .in3(N__31243),
            .lcout(),
            .ltout(\c0.n9584_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9584_bdd_4_lut_LC_6_32_5 .C_ON=1'b0;
    defparam \c0.n9584_bdd_4_lut_LC_6_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9584_bdd_4_lut_LC_6_32_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9584_bdd_4_lut_LC_6_32_5  (
            .in0(N__31605),
            .in1(N__21291),
            .in2(N__20043),
            .in3(N__20040),
            .lcout(),
            .ltout(\c0.n9587_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_6_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_6_32_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_6_32_6  (
            .in0(N__32383),
            .in1(N__20028),
            .in2(N__20013),
            .in3(N__31606),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35406),
            .ce(N__32229),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i86_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i86_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i86_LC_7_18_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i86_LC_7_18_0  (
            .in0(N__19983),
            .in1(N__29974),
            .in2(_gnd_net_),
            .in3(N__19994),
            .lcout(data_in_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i94_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i94_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i94_LC_7_18_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i94_LC_7_18_1  (
            .in0(N__19962),
            .in1(N__29979),
            .in2(_gnd_net_),
            .in3(N__19982),
            .lcout(data_in_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i102_LC_7_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i102_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i102_LC_7_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i102_LC_7_18_2  (
            .in0(N__29977),
            .in1(N__19974),
            .in2(_gnd_net_),
            .in3(N__19961),
            .lcout(data_in_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i118_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i118_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i118_LC_7_18_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i118_LC_7_18_4  (
            .in0(N__19941),
            .in1(N__29972),
            .in2(_gnd_net_),
            .in3(N__19952),
            .lcout(data_in_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i126_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i126_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i126_LC_7_18_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i126_LC_7_18_5  (
            .in0(N__20175),
            .in1(N__29978),
            .in2(_gnd_net_),
            .in3(N__19940),
            .lcout(data_in_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i134_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i134_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i134_LC_7_18_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i134_LC_7_18_6  (
            .in0(N__20154),
            .in1(N__29973),
            .in2(_gnd_net_),
            .in3(N__20174),
            .lcout(data_in_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i142_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i142_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i142_LC_7_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i142_LC_7_18_7  (
            .in0(N__29971),
            .in1(N__20166),
            .in2(_gnd_net_),
            .in3(N__20153),
            .lcout(data_in_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i151_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i151_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i151_LC_7_19_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i151_LC_7_19_0  (
            .in0(N__20259),
            .in1(_gnd_net_),
            .in2(N__29988),
            .in3(N__20144),
            .lcout(data_in_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i146_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i146_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i146_LC_7_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i146_LC_7_19_1  (
            .in0(N__20115),
            .in1(N__29874),
            .in2(_gnd_net_),
            .in3(N__20126),
            .lcout(data_in_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i154_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i154_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i154_LC_7_19_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i154_LC_7_19_2  (
            .in0(N__20106),
            .in1(_gnd_net_),
            .in2(N__29989),
            .in3(N__20114),
            .lcout(data_in_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i162_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i162_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i162_LC_7_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i162_LC_7_19_3  (
            .in0(N__20190),
            .in1(N__29875),
            .in2(_gnd_net_),
            .in3(N__20105),
            .lcout(data_in_20_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_19_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_7_19_4  (
            .in0(N__20282),
            .in1(N__28167),
            .in2(N__20097),
            .in3(N__20337),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i163_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i163_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i163_LC_7_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i163_LC_7_19_7  (
            .in0(N__29882),
            .in1(N__20093),
            .in2(_gnd_net_),
            .in3(N__23078),
            .lcout(data_in_20_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i92_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i92_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i92_LC_7_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i92_LC_7_20_0  (
            .in0(N__29926),
            .in1(N__20085),
            .in2(_gnd_net_),
            .in3(N__20066),
            .lcout(data_in_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_7_20_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_7_20_1  (
            .in0(N__20270),
            .in1(N__28159),
            .in2(N__20289),
            .in3(N__20366),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i159_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i159_LC_7_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i159_LC_7_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i159_LC_7_20_2  (
            .in0(N__20208),
            .in1(N__29927),
            .in2(_gnd_net_),
            .in3(N__20258),
            .lcout(data_in_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_20_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_20_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_7_20_3  (
            .in0(N__20199),
            .in1(N__28157),
            .in2(N__20246),
            .in3(N__20336),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i152_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i152_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i152_LC_7_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i152_LC_7_20_4  (
            .in0(N__29925),
            .in1(N__20379),
            .in2(_gnd_net_),
            .in3(N__20219),
            .lcout(data_in_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i167_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i167_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i167_LC_7_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i167_LC_7_20_5  (
            .in0(N__29928),
            .in1(N__20430),
            .in2(_gnd_net_),
            .in3(N__20207),
            .lcout(data_in_20_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_32_i4_2_lut_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.rx.equal_32_i4_2_lut_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_32_i4_2_lut_LC_7_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.equal_32_i4_2_lut_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__27551),
            .in2(_gnd_net_),
            .in3(N__25873),
            .lcout(n4_adj_1725),
            .ltout(n4_adj_1725_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_20_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_7_20_7  (
            .in0(N__20189),
            .in1(N__28158),
            .in2(N__20193),
            .in3(N__20365),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_506_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_506_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_506_LC_7_21_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_adj_506_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__25926),
            .in2(_gnd_net_),
            .in3(N__27473),
            .lcout(n4044),
            .ltout(n4044_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_7_21_2 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_7_21_2  (
            .in0(N__23058),
            .in1(N__20397),
            .in2(N__20178),
            .in3(N__28156),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_21_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_7_21_3  (
            .in0(N__20335),
            .in1(N__20429),
            .in2(N__28166),
            .in3(N__23057),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_21_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_7_21_4  (
            .in0(N__25823),
            .in1(N__28151),
            .in2(N__20414),
            .in3(N__20334),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i168_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i168_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i168_LC_7_21_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i168_LC_7_21_5  (
            .in0(N__20396),
            .in1(_gnd_net_),
            .in2(N__29987),
            .in3(N__20387),
            .lcout(data_in_20_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i160_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i160_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i160_LC_7_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i160_LC_7_21_6  (
            .in0(N__20388),
            .in1(N__29866),
            .in2(_gnd_net_),
            .in3(N__20378),
            .lcout(data_in_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_7_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_7_21_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_7_21_7  (
            .in0(N__28152),
            .in1(N__25824),
            .in2(N__20352),
            .in3(N__20367),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_7_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__25925),
            .in2(_gnd_net_),
            .in3(N__27474),
            .lcout(n4049),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_566_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_566_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_566_LC_7_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_566_LC_7_22_4  (
            .in0(N__26623),
            .in1(N__25128),
            .in2(N__27330),
            .in3(N__26500),
            .lcout(\c0.n28_adj_1619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7805_LC_7_22_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7805_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7805_LC_7_22_7 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7805_LC_7_22_7  (
            .in0(N__32870),
            .in1(N__31952),
            .in2(N__22057),
            .in3(N__22382),
            .lcout(\c0.n9476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_2056_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.tx2_transmit_2056_LC_7_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_2056_LC_7_23_0 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \c0.tx2_transmit_2056_LC_7_23_0  (
            .in0(N__23667),
            .in1(N__23524),
            .in2(N__20700),
            .in3(N__20789),
            .lcout(\c0.r_SM_Main_2_N_1483_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7965_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7965_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7965_LC_7_23_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7965_LC_7_23_2  (
            .in0(N__25303),
            .in1(N__32806),
            .in2(N__22935),
            .in3(N__31897),
            .lcout(\c0.n9668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_40_i1_3_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_40_i1_3_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_40_i1_3_lut_LC_7_23_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.mux_358_Mux_40_i1_3_lut_LC_7_23_3  (
            .in0(N__20518),
            .in1(N__20676),
            .in2(N__23559),
            .in3(_gnd_net_),
            .lcout(n1903),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i130_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i130_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i130_LC_7_23_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_frame_0___i130_LC_7_23_4  (
            .in0(N__20605),
            .in1(_gnd_net_),
            .in2(N__21045),
            .in3(N__28998),
            .lcout(data_in_field_129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_610_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_610_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_610_LC_7_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_610_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__20604),
            .in2(_gnd_net_),
            .in3(N__26060),
            .lcout(\c0.n8791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i145_LC_7_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i145_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i145_LC_7_23_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i145_LC_7_23_6  (
            .in0(N__26061),
            .in1(N__25998),
            .in2(_gnd_net_),
            .in3(N__28999),
            .lcout(data_in_field_144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i41_LC_7_23_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i41_LC_7_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i41_LC_7_23_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i41_LC_7_23_7  (
            .in0(N__20519),
            .in1(N__29387),
            .in2(_gnd_net_),
            .in3(N__20562),
            .lcout(data_in_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_676_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_676_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_676_LC_7_24_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_676_LC_7_24_0  (
            .in0(N__20978),
            .in1(N__20993),
            .in2(N__20961),
            .in3(N__22818),
            .lcout(\c0.n19_adj_1665 ),
            .ltout(\c0.n19_adj_1665_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7763_2_lut_3_lut_LC_7_24_1 .C_ON=1'b0;
    defparam \c0.i7763_2_lut_3_lut_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7763_2_lut_3_lut_LC_7_24_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \c0.i7763_2_lut_3_lut_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(N__20505),
            .in3(N__20501),
            .lcout(\c0.tx2_transmit_N_1444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5656_2_lut_3_lut_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.i5656_2_lut_3_lut_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5656_2_lut_3_lut_LC_7_24_2 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \c0.i5656_2_lut_3_lut_LC_7_24_2  (
            .in0(N__20502),
            .in1(_gnd_net_),
            .in2(N__20456),
            .in3(N__20436),
            .lcout(\c0.n7194 ),
            .ltout(\c0.n7194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_4_lut_adj_733_LC_7_24_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_4_lut_adj_733_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_4_lut_adj_733_LC_7_24_3 .LUT_INIT=16'b0110001001110011;
    LogicCell40 \c0.i1_4_lut_4_lut_adj_733_LC_7_24_3  (
            .in0(N__23520),
            .in1(N__23659),
            .in2(N__20832),
            .in3(N__20829),
            .lcout(n4839),
            .ltout(n4839_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state__i2_LC_7_24_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state__i2_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state__i2_LC_7_24_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.FRAME_MATCHER_state__i2_LC_7_24_4  (
            .in0(N__23660),
            .in1(N__23589),
            .in2(N__20793),
            .in3(N__20790),
            .lcout(FRAME_MATCHER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i66_LC_7_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i66_LC_7_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i66_LC_7_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i66_LC_7_24_5  (
            .in0(N__21040),
            .in1(N__20718),
            .in2(_gnd_net_),
            .in3(N__28873),
            .lcout(data_in_field_65),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i151_LC_7_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i151_LC_7_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i151_LC_7_24_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i151_LC_7_24_6  (
            .in0(N__24655),
            .in1(_gnd_net_),
            .in2(N__29008),
            .in3(N__25318),
            .lcout(data_in_field_150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i119_LC_7_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i119_LC_7_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i119_LC_7_24_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_frame_0___i119_LC_7_24_7  (
            .in0(N__20880),
            .in1(_gnd_net_),
            .in2(N__24010),
            .in3(N__28869),
            .lcout(data_in_field_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_425__i0_LC_7_25_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i0_LC_7_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i0_LC_7_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i0_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__20696),
            .in2(N__31971),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(\c0.n8113 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i1_LC_7_25_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i1_LC_7_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i1_LC_7_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i1_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__32790),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n8113 ),
            .carryout(\c0.n8114 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i2_LC_7_25_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i2_LC_7_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i2_LC_7_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i2_LC_7_25_2  (
            .in0(_gnd_net_),
            .in1(N__31178),
            .in2(_gnd_net_),
            .in3(N__20682),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(\c0.n8114 ),
            .carryout(\c0.n8115 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i3_LC_7_25_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i3_LC_7_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i3_LC_7_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i3_LC_7_25_3  (
            .in0(_gnd_net_),
            .in1(N__31532),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(\c0.n8115 ),
            .carryout(\c0.n8116 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i4_LC_7_25_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i4_LC_7_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i4_LC_7_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i4_LC_7_25_4  (
            .in0(_gnd_net_),
            .in1(N__32319),
            .in2(_gnd_net_),
            .in3(N__20997),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(\c0.n8116 ),
            .carryout(\c0.n8117 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i5_LC_7_25_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i5_LC_7_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i5_LC_7_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i5_LC_7_25_5  (
            .in0(_gnd_net_),
            .in1(N__20994),
            .in2(_gnd_net_),
            .in3(N__20982),
            .lcout(\c0.byte_transmit_counter2_5 ),
            .ltout(),
            .carryin(\c0.n8117 ),
            .carryout(\c0.n8118 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i6_LC_7_25_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_425__i6_LC_7_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i6_LC_7_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i6_LC_7_25_6  (
            .in0(_gnd_net_),
            .in1(N__20979),
            .in2(_gnd_net_),
            .in3(N__20967),
            .lcout(\c0.byte_transmit_counter2_6 ),
            .ltout(),
            .carryin(\c0.n8118 ),
            .carryout(\c0.n8119 ),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.byte_transmit_counter2_425__i7_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_425__i7_LC_7_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_425__i7_LC_7_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_425__i7_LC_7_25_7  (
            .in0(_gnd_net_),
            .in1(N__20960),
            .in2(_gnd_net_),
            .in3(N__20964),
            .lcout(\c0.byte_transmit_counter2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(N__20946),
            .sr(N__20934));
    defparam \c0.data_in_frame_0___i83_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i83_LC_7_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i83_LC_7_26_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i83_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(N__26146),
            .in2(N__28743),
            .in3(N__32158),
            .lcout(data_in_field_82),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i89_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i89_LC_7_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i89_LC_7_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i89_LC_7_26_1  (
            .in0(N__20922),
            .in1(N__28381),
            .in2(_gnd_net_),
            .in3(N__28558),
            .lcout(data_in_field_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i133_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i133_LC_7_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i133_LC_7_26_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i133_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(N__21182),
            .in2(N__28742),
            .in3(N__33302),
            .lcout(data_in_field_132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i87_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i87_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i87_LC_7_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i87_LC_7_26_3  (
            .in0(N__20875),
            .in1(N__25118),
            .in2(_gnd_net_),
            .in3(N__28557),
            .lcout(data_in_field_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i96_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i96_LC_7_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i96_LC_7_26_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i96_LC_7_26_4  (
            .in0(N__21584),
            .in1(_gnd_net_),
            .in2(N__28744),
            .in3(N__27703),
            .lcout(data_in_field_95),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i100_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i100_LC_7_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i100_LC_7_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i100_LC_7_26_5  (
            .in0(N__21153),
            .in1(N__23824),
            .in2(_gnd_net_),
            .in3(N__28550),
            .lcout(data_in_field_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_577_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_577_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_577_LC_7_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_577_LC_7_26_6  (
            .in0(N__21125),
            .in1(N__23898),
            .in2(N__22128),
            .in3(N__23145),
            .lcout(\c0.n21_adj_1624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i91_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i91_LC_7_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i91_LC_7_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i91_LC_7_26_7  (
            .in0(N__23951),
            .in1(N__32104),
            .in2(_gnd_net_),
            .in3(N__28559),
            .lcout(data_in_field_90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i104_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i104_LC_7_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i104_LC_7_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i104_LC_7_27_0  (
            .in0(N__21075),
            .in1(N__32538),
            .in2(_gnd_net_),
            .in3(N__28643),
            .lcout(data_in_field_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i99_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i99_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i99_LC_7_27_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i99_LC_7_27_1  (
            .in0(N__23707),
            .in1(_gnd_net_),
            .in2(N__28851),
            .in3(N__31462),
            .lcout(data_in_field_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i101_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i101_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i101_LC_7_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i101_LC_7_27_2  (
            .in0(N__21180),
            .in1(N__24845),
            .in2(_gnd_net_),
            .in3(N__28642),
            .lcout(data_in_field_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i69_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i69_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i69_LC_7_27_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i69_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(N__21181),
            .in2(N__28850),
            .in3(N__25511),
            .lcout(data_in_field_68),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i129_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i129_LC_7_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i129_LC_7_27_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i129_LC_7_27_4  (
            .in0(N__25977),
            .in1(N__26179),
            .in2(_gnd_net_),
            .in3(N__28647),
            .lcout(data_in_field_128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i126_LC_7_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i126_LC_7_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i126_LC_7_27_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i126_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(N__21463),
            .in2(N__28848),
            .in3(N__24539),
            .lcout(data_in_field_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i98_LC_7_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i98_LC_7_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i98_LC_7_27_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i98_LC_7_27_6  (
            .in0(N__21019),
            .in1(N__27763),
            .in2(_gnd_net_),
            .in3(N__28654),
            .lcout(data_in_field_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i144_LC_7_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i144_LC_7_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i144_LC_7_27_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i144_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__21577),
            .in2(N__28849),
            .in3(N__21537),
            .lcout(data_in_field_143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_626_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_626_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_626_LC_7_28_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_626_LC_7_28_0  (
            .in0(N__21528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26172),
            .lcout(\c0.n4288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i77_LC_7_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i77_LC_7_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i77_LC_7_28_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i77_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__21505),
            .in2(N__29007),
            .in3(N__25476),
            .lcout(data_in_field_76),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i62_LC_7_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i62_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i62_LC_7_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i62_LC_7_28_2  (
            .in0(N__21465),
            .in1(N__21717),
            .in2(_gnd_net_),
            .in3(N__28863),
            .lcout(data_in_field_61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7920_LC_7_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7920_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7920_LC_7_28_3 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7920_LC_7_28_3  (
            .in0(N__21431),
            .in1(N__32016),
            .in2(N__33024),
            .in3(N__21374),
            .lcout(),
            .ltout(\c0.n9608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9608_bdd_4_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.n9608_bdd_4_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.n9608_bdd_4_lut_LC_7_28_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9608_bdd_4_lut_LC_7_28_4  (
            .in0(N__32946),
            .in1(N__22223),
            .in2(N__21330),
            .in3(N__21327),
            .lcout(\c0.n9147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i110_LC_7_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i110_LC_7_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i110_LC_7_28_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i110_LC_7_28_5  (
            .in0(N__21279),
            .in1(_gnd_net_),
            .in2(N__29005),
            .in3(N__21218),
            .lcout(data_in_field_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i107_LC_7_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i107_LC_7_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i107_LC_7_28_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i107_LC_7_28_6  (
            .in0(N__24082),
            .in1(N__31414),
            .in2(_gnd_net_),
            .in3(N__28856),
            .lcout(data_in_field_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i149_LC_7_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i149_LC_7_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i149_LC_7_28_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_frame_0___i149_LC_7_28_7  (
            .in0(N__21183),
            .in1(_gnd_net_),
            .in2(N__29006),
            .in3(N__32497),
            .lcout(data_in_field_148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_515_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_515_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_515_LC_7_29_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_515_LC_7_29_0  (
            .in0(N__21794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24249),
            .lcout(\c0.n8942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i58_LC_7_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i58_LC_7_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i58_LC_7_29_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_frame_0___i58_LC_7_29_1  (
            .in0(N__22056),
            .in1(_gnd_net_),
            .in2(N__21662),
            .in3(N__28868),
            .lcout(data_in_field_57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_698_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_698_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_698_LC_7_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_698_LC_7_29_2  (
            .in0(N__24959),
            .in1(N__22023),
            .in2(_gnd_net_),
            .in3(N__22531),
            .lcout(\c0.n4390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_730_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_730_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_730_LC_7_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_730_LC_7_29_3  (
            .in0(N__21942),
            .in1(N__21892),
            .in2(N__21828),
            .in3(N__21675),
            .lcout(\c0.n4197 ),
            .ltout(\c0.n4197_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_545_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_545_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_545_LC_7_29_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_545_LC_7_29_4  (
            .in0(N__21795),
            .in1(_gnd_net_),
            .in2(N__21753),
            .in3(_gnd_net_),
            .lcout(\c0.n8834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_619_LC_7_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_619_LC_7_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_619_LC_7_29_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_619_LC_7_29_5  (
            .in0(_gnd_net_),
            .in1(N__31407),
            .in2(_gnd_net_),
            .in3(N__21611),
            .lcout(\c0.n4399 ),
            .ltout(\c0.n4399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_541_LC_7_29_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_541_LC_7_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_541_LC_7_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_541_LC_7_29_6  (
            .in0(N__21718),
            .in1(N__25454),
            .in2(N__21693),
            .in3(N__21686),
            .lcout(\c0.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i122_LC_7_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i122_LC_7_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i122_LC_7_29_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i122_LC_7_29_7  (
            .in0(N__21654),
            .in1(N__21612),
            .in2(_gnd_net_),
            .in3(N__28867),
            .lcout(data_in_field_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9572_bdd_4_lut_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.n9572_bdd_4_lut_LC_7_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.n9572_bdd_4_lut_LC_7_30_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n9572_bdd_4_lut_LC_7_30_0  (
            .in0(N__32945),
            .in1(N__22475),
            .in2(N__22809),
            .in3(N__22431),
            .lcout(\c0.n9165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_707_LC_7_30_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_707_LC_7_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_707_LC_7_30_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_707_LC_7_30_1  (
            .in0(N__22157),
            .in1(N__25512),
            .in2(N__22422),
            .in3(N__22383),
            .lcout(\c0.n8887 ),
            .ltout(\c0.n8887_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_705_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_705_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_705_LC_7_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_705_LC_7_30_2  (
            .in0(N__22262),
            .in1(N__32598),
            .in2(N__22332),
            .in3(N__22328),
            .lcout(\c0.n8893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i111_LC_7_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i111_LC_7_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i111_LC_7_30_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i111_LC_7_30_3  (
            .in0(N__27308),
            .in1(N__22294),
            .in2(_gnd_net_),
            .in3(N__29056),
            .lcout(data_in_field_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_632_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_632_LC_7_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_632_LC_7_30_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_632_LC_7_30_4  (
            .in0(N__22263),
            .in1(N__22238),
            .in2(_gnd_net_),
            .in3(N__32599),
            .lcout(),
            .ltout(\c0.n4240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_7_30_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_7_30_5  (
            .in0(N__22164),
            .in1(N__26628),
            .in2(N__22227),
            .in3(N__22224),
            .lcout(\c0.n44_adj_1609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_553_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_553_LC_7_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_553_LC_7_30_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_553_LC_7_30_6  (
            .in0(_gnd_net_),
            .in1(N__27307),
            .in2(_gnd_net_),
            .in3(N__24298),
            .lcout(\c0.n4553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_630_LC_7_30_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_630_LC_7_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_630_LC_7_30_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_630_LC_7_30_7  (
            .in0(N__22158),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25513),
            .lcout(\c0.n8964 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_7_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_7_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_7_31_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_7_31_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22116),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35407),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_7_31_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_7_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_7_31_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_3_lut_LC_7_31_2  (
            .in0(N__31569),
            .in1(N__32348),
            .in2(_gnd_net_),
            .in3(N__31179),
            .lcout(\c0.n18_adj_1666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_652_LC_7_31_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_652_LC_7_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_652_LC_7_31_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_652_LC_7_31_3  (
            .in0(N__24003),
            .in1(N__22574),
            .in2(N__22737),
            .in3(N__22805),
            .lcout(\c0.n8810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1042_2_lut_LC_7_31_5 .C_ON=1'b0;
    defparam \c0.i1042_2_lut_LC_7_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1042_2_lut_LC_7_31_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1042_2_lut_LC_7_31_5  (
            .in0(_gnd_net_),
            .in1(N__25218),
            .in2(_gnd_net_),
            .in3(N__25339),
            .lcout(\c0.n1645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7935_LC_7_31_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7935_LC_7_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7935_LC_7_31_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7935_LC_7_31_6  (
            .in0(N__24450),
            .in1(N__32947),
            .in2(N__22736),
            .in3(N__32030),
            .lcout(),
            .ltout(\c0.n9632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9632_bdd_4_lut_LC_7_31_7 .C_ON=1'b0;
    defparam \c0.n9632_bdd_4_lut_LC_7_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.n9632_bdd_4_lut_LC_7_31_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9632_bdd_4_lut_LC_7_31_7  (
            .in0(N__32948),
            .in1(N__22686),
            .in2(N__22626),
            .in3(N__22623),
            .lcout(\c0.n9135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7925_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7925_LC_7_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7925_LC_7_32_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7925_LC_7_32_0  (
            .in0(N__32054),
            .in1(N__24011),
            .in2(N__22575),
            .in3(N__32848),
            .lcout(),
            .ltout(\c0.n9620_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9620_bdd_4_lut_LC_7_32_1 .C_ON=1'b0;
    defparam \c0.n9620_bdd_4_lut_LC_7_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9620_bdd_4_lut_LC_7_32_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9620_bdd_4_lut_LC_7_32_1  (
            .in0(N__32849),
            .in1(N__24604),
            .in2(N__22536),
            .in3(N__27327),
            .lcout(\c0.n9141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7930_LC_7_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7930_LC_7_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7930_LC_7_32_2 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7930_LC_7_32_2  (
            .in0(N__32055),
            .in1(N__32850),
            .in2(N__25138),
            .in3(N__22533),
            .lcout(),
            .ltout(\c0.n9626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9626_bdd_4_lut_LC_7_32_3 .C_ON=1'b0;
    defparam \c0.n9626_bdd_4_lut_LC_7_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9626_bdd_4_lut_LC_7_32_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9626_bdd_4_lut_LC_7_32_3  (
            .in0(N__32851),
            .in1(N__26404),
            .in2(N__22479),
            .in3(N__27081),
            .lcout(),
            .ltout(\c0.n9138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7940_LC_7_32_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7940_LC_7_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7940_LC_7_32_4 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7940_LC_7_32_4  (
            .in0(N__31570),
            .in1(N__22911),
            .in2(N__22905),
            .in3(N__31192),
            .lcout(),
            .ltout(\c0.n9614_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9614_bdd_4_lut_LC_7_32_5 .C_ON=1'b0;
    defparam \c0.n9614_bdd_4_lut_LC_7_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9614_bdd_4_lut_LC_7_32_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n9614_bdd_4_lut_LC_7_32_5  (
            .in0(N__22902),
            .in1(N__22884),
            .in2(N__22878),
            .in3(N__31571),
            .lcout(),
            .ltout(\c0.n9617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_7_32_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_7_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_7_32_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_7_32_6  (
            .in0(N__31572),
            .in1(N__31107),
            .in2(N__22875),
            .in3(N__32349),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35411),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i83_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i83_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i83_LC_9_20_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i83_LC_9_20_0  (
            .in0(N__22863),
            .in1(_gnd_net_),
            .in2(N__30034),
            .in3(N__23165),
            .lcout(data_in_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i91_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i91_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i91_LC_9_20_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i91_LC_9_20_1  (
            .in0(N__22854),
            .in1(N__30008),
            .in2(_gnd_net_),
            .in3(N__22862),
            .lcout(data_in_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i99_LC_9_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i99_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i99_LC_9_20_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i99_LC_9_20_2  (
            .in0(N__22845),
            .in1(_gnd_net_),
            .in2(N__30035),
            .in3(N__22853),
            .lcout(data_in_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i107_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i107_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i107_LC_9_20_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i107_LC_9_20_3  (
            .in0(N__22836),
            .in1(N__30006),
            .in2(_gnd_net_),
            .in3(N__22844),
            .lcout(data_in_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i115_LC_9_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i115_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i115_LC_9_20_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i115_LC_9_20_4  (
            .in0(N__22827),
            .in1(_gnd_net_),
            .in2(N__30033),
            .in3(N__22835),
            .lcout(data_in_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i123_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i123_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i123_LC_9_20_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i123_LC_9_20_5  (
            .in0(N__23115),
            .in1(N__30007),
            .in2(_gnd_net_),
            .in3(N__22826),
            .lcout(data_in_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i131_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i131_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i131_LC_9_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i131_LC_9_20_6  (
            .in0(N__30005),
            .in1(N__23097),
            .in2(_gnd_net_),
            .in3(N__23114),
            .lcout(data_in_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i147_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i147_LC_9_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i147_LC_9_21_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i147_LC_9_21_0  (
            .in0(N__29990),
            .in1(N__23105),
            .in2(_gnd_net_),
            .in3(N__23067),
            .lcout(data_in_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i139_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i139_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i139_LC_9_21_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i139_LC_9_21_1  (
            .in0(N__23106),
            .in1(N__29992),
            .in2(_gnd_net_),
            .in3(N__23096),
            .lcout(data_in_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i155_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i155_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i155_LC_9_21_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i155_LC_9_21_6  (
            .in0(N__29991),
            .in1(N__23085),
            .in2(_gnd_net_),
            .in3(N__23066),
            .lcout(data_in_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5633_2_lut_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.rx.i5633_2_lut_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5633_2_lut_LC_9_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i5633_2_lut_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__27529),
            .in2(_gnd_net_),
            .in3(N__25863),
            .lcout(n7171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9668_bdd_4_lut_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.n9668_bdd_4_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9668_bdd_4_lut_LC_9_23_1 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n9668_bdd_4_lut_LC_9_23_1  (
            .in0(N__23043),
            .in1(N__26457),
            .in2(N__25809),
            .in3(N__32978),
            .lcout(\c0.n9671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_567_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_567_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_567_LC_9_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_567_LC_9_23_2  (
            .in0(N__23034),
            .in1(N__23016),
            .in2(N__26313),
            .in3(N__22995),
            .lcout(),
            .ltout(\c0.n29_adj_1620_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i159_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i159_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i159_LC_9_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i159_LC_9_23_3  (
            .in0(N__22950),
            .in1(N__23964),
            .in2(N__22938),
            .in3(N__23685),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35366),
            .ce(N__29009),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_42_i1_3_lut_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_42_i1_3_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_42_i1_3_lut_LC_9_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.mux_358_Mux_42_i1_3_lut_LC_9_24_0  (
            .in0(N__24089),
            .in1(N__26995),
            .in2(_gnd_net_),
            .in3(N__23551),
            .lcout(n1901),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i43_LC_9_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i43_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i43_LC_9_24_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i43_LC_9_24_1  (
            .in0(N__26996),
            .in1(_gnd_net_),
            .in2(N__30030),
            .in3(N__23577),
            .lcout(data_in_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7655_2_lut_1_lut_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.i7655_2_lut_1_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7655_2_lut_1_lut_LC_9_24_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.i7655_2_lut_1_lut_LC_9_24_2  (
            .in0(N__23669),
            .in1(N__23550),
            .in2(_gnd_net_),
            .in3(N__23609),
            .lcout(n9262),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i51_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i51_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i51_LC_9_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i51_LC_9_24_3  (
            .in0(N__29993),
            .in1(N__23190),
            .in2(_gnd_net_),
            .in3(N__23576),
            .lcout(data_in_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_358_Mux_50_i1_3_lut_LC_9_24_4 .C_ON=1'b0;
    defparam \c0.mux_358_Mux_50_i1_3_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_358_Mux_50_i1_3_lut_LC_9_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_358_Mux_50_i1_3_lut_LC_9_24_4  (
            .in0(N__23575),
            .in1(N__26147),
            .in2(_gnd_net_),
            .in3(N__23549),
            .lcout(n1893),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i59_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i59_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i59_LC_9_24_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i59_LC_9_24_5  (
            .in0(N__23181),
            .in1(_gnd_net_),
            .in2(N__30031),
            .in3(N__23189),
            .lcout(data_in_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i67_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i67_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i67_LC_9_24_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i67_LC_9_24_6  (
            .in0(N__23154),
            .in1(N__29995),
            .in2(_gnd_net_),
            .in3(N__23180),
            .lcout(data_in_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i75_LC_9_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i75_LC_9_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i75_LC_9_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i75_LC_9_24_7  (
            .in0(N__29994),
            .in1(N__23153),
            .in2(_gnd_net_),
            .in3(N__23172),
            .lcout(data_in_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_724_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_724_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_724_LC_9_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_724_LC_9_25_0  (
            .in0(N__24888),
            .in1(N__26654),
            .in2(N__23787),
            .in3(N__23144),
            .lcout(\c0.n4562 ),
            .ltout(\c0.n4562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_582_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_582_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_582_LC_9_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_582_LC_9_25_1  (
            .in0(N__26004),
            .in1(N__26267),
            .in2(N__23118),
            .in3(N__26750),
            .lcout(\c0.n8837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_654_LC_9_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_654_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_654_LC_9_25_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_654_LC_9_25_3  (
            .in0(N__32116),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26605),
            .lcout(),
            .ltout(\c0.n4235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_549_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_549_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_549_LC_9_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_549_LC_9_25_4  (
            .in0(N__23877),
            .in1(N__27390),
            .in2(N__23862),
            .in3(N__23859),
            .lcout(\c0.n25_adj_1614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_618_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_618_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_618_LC_9_25_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_618_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__27932),
            .in2(_gnd_net_),
            .in3(N__26219),
            .lcout(\c0.n4365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_649_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_649_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_649_LC_9_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_649_LC_9_25_6  (
            .in0(N__27787),
            .in1(N__24184),
            .in2(N__23853),
            .in3(N__24291),
            .lcout(\c0.n4534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_725_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_725_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_725_LC_9_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_725_LC_9_25_7  (
            .in0(N__26655),
            .in1(N__23786),
            .in2(_gnd_net_),
            .in3(N__24889),
            .lcout(\c0.n8846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i71_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i71_LC_9_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i71_LC_9_26_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0___i71_LC_9_26_0  (
            .in0(N__27067),
            .in1(_gnd_net_),
            .in2(N__29053),
            .in3(N__24656),
            .lcout(data_in_field_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i67_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i67_LC_9_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i67_LC_9_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i67_LC_9_26_1  (
            .in0(N__23721),
            .in1(N__31722),
            .in2(_gnd_net_),
            .in3(N__28957),
            .lcout(data_in_field_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i147_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i147_LC_9_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i147_LC_9_26_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i147_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__23720),
            .in2(N__29052),
            .in3(N__26606),
            .lcout(data_in_field_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_565_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_565_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_565_LC_9_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_565_LC_9_26_3  (
            .in0(N__28320),
            .in1(N__32447),
            .in2(N__24459),
            .in3(N__23894),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_721_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_721_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_721_LC_9_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_721_LC_9_26_4  (
            .in0(N__27066),
            .in1(N__27704),
            .in2(_gnd_net_),
            .in3(N__27411),
            .lcout(\c0.n8918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i75_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i75_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i75_LC_9_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i75_LC_9_26_5  (
            .in0(N__24090),
            .in1(N__31673),
            .in2(_gnd_net_),
            .in3(N__28961),
            .lcout(data_in_field_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_568_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_568_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_568_LC_9_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_568_LC_9_26_6  (
            .in0(N__24048),
            .in1(N__24012),
            .in2(N__23973),
            .in3(N__28388),
            .lcout(\c0.n27_adj_1621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i123_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i123_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i123_LC_9_26_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i123_LC_9_26_7  (
            .in0(N__27412),
            .in1(N__23952),
            .in2(_gnd_net_),
            .in3(N__28953),
            .lcout(data_in_field_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_571_LC_9_27_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_571_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_571_LC_9_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_571_LC_9_27_1  (
            .in0(N__33314),
            .in1(N__24579),
            .in2(_gnd_net_),
            .in3(N__27896),
            .lcout(\c0.n4473 ),
            .ltout(\c0.n4473_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_573_LC_9_27_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_573_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_573_LC_9_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_573_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__27659),
            .in2(N__23901),
            .in3(N__26769),
            .lcout(\c0.n9010 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_597_LC_9_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_597_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_597_LC_9_27_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_597_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__31460),
            .in2(_gnd_net_),
            .in3(N__24846),
            .lcout(\c0.n4511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_719_LC_9_27_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_719_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_719_LC_9_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_719_LC_9_27_4  (
            .in0(N__31461),
            .in1(N__25804),
            .in2(N__24987),
            .in3(N__32513),
            .lcout(\c0.n4244 ),
            .ltout(\c0.n4244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_738_LC_9_27_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_738_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_738_LC_9_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_738_LC_9_27_5  (
            .in0(N__28343),
            .in1(N__33247),
            .in2(N__23880),
            .in3(N__24224),
            .lcout(\c0.n8995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i103_LC_9_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i103_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i103_LC_9_27_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i103_LC_9_27_6  (
            .in0(N__24580),
            .in1(N__24654),
            .in2(_gnd_net_),
            .in3(N__28924),
            .lcout(data_in_field_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_716_LC_9_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_716_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_716_LC_9_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_716_LC_9_27_7  (
            .in0(N__24549),
            .in1(N__24504),
            .in2(_gnd_net_),
            .in3(N__24984),
            .lcout(\c0.n18_adj_1618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_615_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_615_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_615_LC_9_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_615_LC_9_28_0  (
            .in0(N__25523),
            .in1(N__24449),
            .in2(_gnd_net_),
            .in3(N__24402),
            .lcout(\c0.n8912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_9_28_1 .C_ON=1'b0;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_3_lut_4_lut_LC_9_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_2_lut_3_lut_4_lut_LC_9_28_1  (
            .in0(N__24372),
            .in1(N__31678),
            .in2(N__33257),
            .in3(N__28398),
            .lcout(\c0.n16_adj_1591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i117_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i117_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i117_LC_9_28_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i117_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__24331),
            .in2(N__29071),
            .in3(N__24242),
            .lcout(data_in_field_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i85_LC_9_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i85_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i85_LC_9_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i85_LC_9_28_3  (
            .in0(N__24332),
            .in1(N__24986),
            .in2(_gnd_net_),
            .in3(N__29046),
            .lcout(data_in_field_84),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7875_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7875_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7875_LC_9_28_4 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7875_LC_9_28_4  (
            .in0(N__24292),
            .in1(N__24240),
            .in2(N__33204),
            .in3(N__31975),
            .lcout(\c0.n9560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_585_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_585_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_585_LC_9_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_585_LC_9_28_5  (
            .in0(N__24241),
            .in1(N__24225),
            .in2(N__24189),
            .in3(N__24985),
            .lcout(\c0.n16_adj_1629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i113_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i113_LC_9_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i113_LC_9_28_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i113_LC_9_28_7  (
            .in0(N__24127),
            .in1(N__27033),
            .in2(_gnd_net_),
            .in3(N__29042),
            .lcout(data_in_field_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_562_LC_9_29_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_562_LC_9_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_562_LC_9_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_562_LC_9_29_0  (
            .in0(N__24800),
            .in1(N__25059),
            .in2(N__25044),
            .in3(N__25023),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7880_LC_9_29_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7880_LC_9_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7880_LC_9_29_3 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7880_LC_9_29_3  (
            .in0(N__24980),
            .in1(N__31976),
            .in2(N__33135),
            .in3(N__24958),
            .lcout(\c0.n9566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_612_LC_9_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_612_LC_9_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_612_LC_9_29_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_612_LC_9_29_4  (
            .in0(_gnd_net_),
            .in1(N__26108),
            .in2(_gnd_net_),
            .in3(N__26186),
            .lcout(\c0.n8954 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9560_bdd_4_lut_LC_9_29_6 .C_ON=1'b0;
    defparam \c0.n9560_bdd_4_lut_LC_9_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.n9560_bdd_4_lut_LC_9_29_6 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \c0.n9560_bdd_4_lut_LC_9_29_6  (
            .in0(N__24909),
            .in1(N__24902),
            .in2(N__33136),
            .in3(N__24856),
            .lcout(\c0.n9171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_587_LC_9_29_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_587_LC_9_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_587_LC_9_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_587_LC_9_29_7  (
            .in0(N__24813),
            .in1(N__24801),
            .in2(N__25079),
            .in3(N__24789),
            .lcout(\c0.n17_adj_1630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7975_LC_9_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7975_LC_9_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7975_LC_9_30_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7975_LC_9_30_0  (
            .in0(N__32988),
            .in1(N__32509),
            .in2(N__24684),
            .in3(N__32037),
            .lcout(\c0.n9680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i157_LC_9_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i157_LC_9_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i157_LC_9_30_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i157_LC_9_30_3  (
            .in0(N__26030),
            .in1(N__24729),
            .in2(N__24720),
            .in3(N__24690),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35412),
            .ce(N__29073),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_9_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_9_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_9_30_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_9_30_4  (
            .in0(N__31343),
            .in1(N__32631),
            .in2(N__24675),
            .in3(N__31255),
            .lcout(\c0.n22_adj_1679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9566_bdd_4_lut_LC_9_31_1 .C_ON=1'b0;
    defparam \c0.n9566_bdd_4_lut_LC_9_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9566_bdd_4_lut_LC_9_31_1 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n9566_bdd_4_lut_LC_9_31_1  (
            .in0(N__33023),
            .in1(N__25527),
            .in2(N__25482),
            .in3(N__25437),
            .lcout(),
            .ltout(\c0.n9168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7890_LC_9_31_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7890_LC_9_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7890_LC_9_31_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7890_LC_9_31_2  (
            .in0(N__25428),
            .in1(N__31614),
            .in2(N__25419),
            .in3(N__31242),
            .lcout(\c0.n9554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9554_bdd_4_lut_LC_9_31_5 .C_ON=1'b0;
    defparam \c0.n9554_bdd_4_lut_LC_9_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9554_bdd_4_lut_LC_9_31_5 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n9554_bdd_4_lut_LC_9_31_5  (
            .in0(N__31615),
            .in1(N__25416),
            .in2(N__25404),
            .in3(N__25383),
            .lcout(),
            .ltout(\c0.n9557_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_9_31_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_9_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_9_31_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_9_31_6  (
            .in0(N__25377),
            .in1(N__31616),
            .in2(N__25368),
            .in3(N__32382),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35417),
            .ce(N__32277),
            .sr(_gnd_net_));
    defparam \c0.rx.i7410_3_lut_4_lut_LC_9_32_0 .C_ON=1'b0;
    defparam \c0.rx.i7410_3_lut_4_lut_LC_9_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7410_3_lut_4_lut_LC_9_32_0 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \c0.rx.i7410_3_lut_4_lut_LC_9_32_0  (
            .in0(N__27518),
            .in1(N__30792),
            .in2(N__27570),
            .in3(N__25947),
            .lcout(n5185),
            .ltout(n5185_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_9_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_9_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_9_32_1 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_9_32_1  (
            .in0(N__25950),
            .in1(N__27519),
            .in2(N__25350),
            .in3(N__27568),
            .lcout(r_Bit_Index_2_adj_1731),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i7406_4_lut_LC_9_32_2 .C_ON=1'b0;
    defparam \c0.rx.i7406_4_lut_LC_9_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7406_4_lut_LC_9_32_2 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \c0.rx.i7406_4_lut_LC_9_32_2  (
            .in0(N__30567),
            .in1(N__30724),
            .in2(N__30657),
            .in3(N__30791),
            .lcout(n9077),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_722_LC_9_32_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_722_LC_9_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_722_LC_9_32_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_722_LC_9_32_3  (
            .in0(N__25347),
            .in1(N__25278),
            .in2(N__25224),
            .in3(N__25140),
            .lcout(\c0.n8915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_9_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_9_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_9_32_4 .LUT_INIT=16'b1000100000101000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_9_32_4  (
            .in0(N__25935),
            .in1(N__25843),
            .in2(N__25906),
            .in3(N__25949),
            .lcout(r_Bit_Index_1_adj_1732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i635_2_lut_LC_9_32_5 .C_ON=1'b0;
    defparam \c0.rx.i635_2_lut_LC_9_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i635_2_lut_LC_9_32_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i635_2_lut_LC_9_32_5  (
            .in0(N__25842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25895),
            .lcout(n2185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_9_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_9_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_9_32_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_9_32_7  (
            .in0(N__25948),
            .in1(N__25896),
            .in2(_gnd_net_),
            .in3(N__25934),
            .lcout(r_Bit_Index_0_adj_1733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_29_i4_2_lut_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.rx.equal_29_i4_2_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_29_i4_2_lut_LC_10_22_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.equal_29_i4_2_lut_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__27544),
            .in2(_gnd_net_),
            .in3(N__25875),
            .lcout(n4_adj_1724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_653_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_653_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_653_LC_10_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_653_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__25791),
            .in2(_gnd_net_),
            .in3(N__32514),
            .lcout(\c0.n8770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_3_lut_LC_10_24_3 .C_ON=1'b0;
    defparam \c0.i3_2_lut_3_lut_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_3_lut_LC_10_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_2_lut_3_lut_LC_10_24_3  (
            .in0(N__32117),
            .in1(N__26612),
            .in2(_gnd_net_),
            .in3(N__25752),
            .lcout(\c0.n16_adj_1657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_657_LC_10_24_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_657_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_657_LC_10_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_657_LC_10_24_5  (
            .in0(N__25711),
            .in1(N__25686),
            .in2(N__25673),
            .in3(N__25647),
            .lcout(),
            .ltout(\c0.n22_adj_1655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_659_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_659_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_659_LC_10_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_659_LC_10_24_6  (
            .in0(N__25623),
            .in1(N__31731),
            .in2(N__25617),
            .in3(N__25614),
            .lcout(\c0.n24_adj_1658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i153_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i153_LC_10_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i153_LC_10_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i153_LC_10_25_1  (
            .in0(N__28319),
            .in1(N__25572),
            .in2(N__25566),
            .in3(N__25542),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(N__29047),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7855_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7855_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7855_LC_10_25_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7855_LC_10_25_2  (
            .in0(N__26080),
            .in1(N__32884),
            .in2(N__32036),
            .in3(N__26229),
            .lcout(),
            .ltout(\c0.n9536_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9536_bdd_4_lut_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.n9536_bdd_4_lut_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9536_bdd_4_lut_LC_10_25_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n9536_bdd_4_lut_LC_10_25_3  (
            .in0(N__32885),
            .in1(N__26223),
            .in2(N__26190),
            .in3(N__26187),
            .lcout(),
            .ltout(\c0.n9539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_25_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_25_4  (
            .in0(N__27195),
            .in1(N__31383),
            .in2(N__26154),
            .in3(N__31203),
            .lcout(\c0.n22_adj_1661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i115_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i115_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i115_LC_10_26_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i115_LC_10_26_0  (
            .in0(N__26096),
            .in1(N__26151),
            .in2(_gnd_net_),
            .in3(N__28962),
            .lcout(data_in_field_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7820_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7820_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7820_LC_10_26_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7820_LC_10_26_1  (
            .in0(N__27410),
            .in1(N__26095),
            .in2(N__33090),
            .in3(N__31993),
            .lcout(\c0.n9494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_584_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_584_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_584_LC_10_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_584_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(N__26079),
            .in2(_gnd_net_),
            .in3(N__26501),
            .lcout(\c0.n8971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_581_LC_10_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_581_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_581_LC_10_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_581_LC_10_26_3  (
            .in0(_gnd_net_),
            .in1(N__26592),
            .in2(_gnd_net_),
            .in3(N__32160),
            .lcout(\c0.n6_adj_1628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i97_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i97_LC_10_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i97_LC_10_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0___i97_LC_10_26_4  (
            .in0(N__27647),
            .in1(N__25997),
            .in2(_gnd_net_),
            .in3(N__28966),
            .lcout(data_in_field_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_595_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_595_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_595_LC_10_26_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_595_LC_10_26_5  (
            .in0(_gnd_net_),
            .in1(N__31712),
            .in2(_gnd_net_),
            .in3(N__27646),
            .lcout(),
            .ltout(\c0.n8840_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_599_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_599_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_599_LC_10_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_599_LC_10_26_6  (
            .in0(N__26554),
            .in1(N__26783),
            .in2(N__26772),
            .in3(N__26768),
            .lcout(\c0.n4309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i124_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i124_LC_10_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i124_LC_10_26_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_frame_0___i124_LC_10_26_7  (
            .in0(_gnd_net_),
            .in1(N__26738),
            .in2(N__29054),
            .in3(N__26659),
            .lcout(data_in_field_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7989_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7989_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7989_LC_10_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7989_LC_10_27_0  (
            .in0(N__26591),
            .in1(N__33018),
            .in2(N__26238),
            .in3(N__31977),
            .lcout(),
            .ltout(\c0.n9698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9698_bdd_4_lut_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.n9698_bdd_4_lut_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n9698_bdd_4_lut_LC_10_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n9698_bdd_4_lut_LC_10_27_1  (
            .in0(N__33019),
            .in1(N__26555),
            .in2(N__26508),
            .in3(N__26505),
            .lcout(),
            .ltout(\c0.n9701_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_10_27_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_10_27_2  (
            .in0(N__31379),
            .in1(N__27009),
            .in2(N__26466),
            .in3(N__31233),
            .lcout(\c0.n22_adj_1681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_713_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_713_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_713_LC_10_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_713_LC_10_27_3  (
            .in0(N__26463),
            .in1(N__32171),
            .in2(N__26408),
            .in3(N__26346),
            .lcout(\c0.n8819 ),
            .ltout(\c0.n8819_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_624_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_624_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_624_LC_10_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_624_LC_10_27_4  (
            .in0(N__26303),
            .in1(N__26292),
            .in2(N__26274),
            .in3(N__26271),
            .lcout(),
            .ltout(\c0.n21_adj_1644_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i155_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i155_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i155_LC_10_27_5 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.data_in_frame_0___i155_LC_10_27_5  (
            .in0(N__27489),
            .in1(_gnd_net_),
            .in2(N__26256),
            .in3(N__26253),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(N__29048),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_547_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_547_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_547_LC_10_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_547_LC_10_28_0  (
            .in0(N__27372),
            .in1(N__32554),
            .in2(N__27345),
            .in3(N__27329),
            .lcout(\c0.n26_adj_1613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_548_LC_10_28_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_548_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_548_LC_10_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_548_LC_10_28_2  (
            .in0(N__27276),
            .in1(N__27162),
            .in2(N__27270),
            .in3(N__27240),
            .lcout(),
            .ltout(\c0.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i161_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i161_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i161_LC_10_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_frame_0___i161_LC_10_28_3  (
            .in0(N__27222),
            .in1(N__27213),
            .in2(N__27207),
            .in3(N__27204),
            .lcout(\c0.data_in_frame_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(N__29030),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_535_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_535_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_535_LC_10_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_535_LC_10_28_4  (
            .in0(N__27176),
            .in1(N__27161),
            .in2(N__27147),
            .in3(N__27123),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i163_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i163_LC_10_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i163_LC_10_28_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_in_frame_0___i163_LC_10_28_5  (
            .in0(N__27102),
            .in1(N__27077),
            .in2(N__27048),
            .in3(N__27034),
            .lcout(\c0.data_in_frame_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(N__29030),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i35_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i35_LC_10_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i35_LC_10_29_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i35_LC_10_29_1  (
            .in0(N__29842),
            .in1(N__26959),
            .in2(_gnd_net_),
            .in3(N__27003),
            .lcout(data_in_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35408),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i6_1_lut_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.tx2.i6_1_lut_LC_10_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i6_1_lut_LC_10_29_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.i6_1_lut_LC_10_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26942),
            .lcout(\c0.tx2.n4880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_620_LC_10_29_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_620_LC_10_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_620_LC_10_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_620_LC_10_29_7  (
            .in0(N__27614),
            .in1(N__26853),
            .in2(N__26838),
            .in3(N__26823),
            .lcout(\c0.n20_adj_1642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_10_30_0.C_ON=1'b0;
    defparam i5_4_lut_LC_10_30_0.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_10_30_0.LUT_INIT=16'b0000000000100000;
    LogicCell40 i5_4_lut_LC_10_30_0 (
            .in0(N__30450),
            .in1(N__31016),
            .in2(N__30530),
            .in3(N__30489),
            .lcout(),
            .ltout(n12_adj_1753_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7695_4_lut_LC_10_30_1.C_ON=1'b0;
    defparam i7695_4_lut_LC_10_30_1.SEQ_MODE=4'b0000;
    defparam i7695_4_lut_LC_10_30_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 i7695_4_lut_LC_10_30_1 (
            .in0(N__30965),
            .in1(N__31074),
            .in2(N__27480),
            .in3(N__30411),
            .lcout(n9246),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_10_30_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.rx.i1_4_lut_LC_10_30_2  (
            .in0(N__31073),
            .in1(N__27440),
            .in2(N__31021),
            .in3(N__30964),
            .lcout(r_SM_Main_2_N_1537_2),
            .ltout(r_SM_Main_2_N_1537_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_10_30_3 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_10_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_10_30_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.rx.i2_4_lut_LC_10_30_3  (
            .in0(N__30641),
            .in1(N__30721),
            .in2(N__27477),
            .in3(N__30786),
            .lcout(\c0.rx.n4090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5849_3_lut_LC_10_30_5 .C_ON=1'b0;
    defparam \c0.rx.i5849_3_lut_LC_10_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5849_3_lut_LC_10_30_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.rx.i5849_3_lut_LC_10_30_5  (
            .in0(N__30488),
            .in1(N__30410),
            .in2(_gnd_net_),
            .in3(N__30449),
            .lcout(\c0.rx.n7393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_10_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_10_30_6 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_10_30_6  (
            .in0(N__31012),
            .in1(N__30909),
            .in2(N__30876),
            .in3(N__30978),
            .lcout(r_Clock_Count_7_adj_1727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35413),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_590_LC_10_30_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_590_LC_10_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_590_LC_10_30_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_590_LC_10_30_7  (
            .in0(_gnd_net_),
            .in1(N__27720),
            .in2(_gnd_net_),
            .in3(N__27425),
            .lcout(\c0.n4537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i6_4_lut_LC_10_31_0 .C_ON=1'b0;
    defparam \c0.rx.i6_4_lut_LC_10_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i6_4_lut_LC_10_31_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.rx.i6_4_lut_LC_10_31_0  (
            .in0(N__30491),
            .in1(N__30451),
            .in2(N__27594),
            .in3(N__30963),
            .lcout(\c0.rx.r_SM_Main_2_N_1543_0 ),
            .ltout(\c0.rx.r_SM_Main_2_N_1543_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_10_31_1 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_10_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_10_31_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \c0.rx.i2_2_lut_LC_10_31_1  (
            .in0(N__28163),
            .in1(_gnd_net_),
            .in2(N__27375),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n6_adj_1751_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_10_31_2.C_ON=1'b0;
    defparam i1_4_lut_LC_10_31_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_10_31_2.LUT_INIT=16'b1100110011101100;
    LogicCell40 i1_4_lut_LC_10_31_2 (
            .in0(N__30714),
            .in1(N__30658),
            .in2(N__27798),
            .in3(N__30783),
            .lcout(n30),
            .ltout(n30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_10_31_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_10_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_10_31_3 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_10_31_3  (
            .in0(N__30504),
            .in1(N__30523),
            .in2(N__27795),
            .in3(N__30873),
            .lcout(r_Clock_Count_0_adj_1730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35418),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_643_LC_10_31_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_643_LC_10_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_643_LC_10_31_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_643_LC_10_31_6  (
            .in0(N__27786),
            .in1(N__27727),
            .in2(_gnd_net_),
            .in3(N__27671),
            .lcout(\c0.n4296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5_4_lut_LC_10_31_7 .C_ON=1'b0;
    defparam \c0.rx.i5_4_lut_LC_10_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5_4_lut_LC_10_31_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.rx.i5_4_lut_LC_10_31_7  (
            .in0(N__31072),
            .in1(N__30522),
            .in2(N__31022),
            .in3(N__30412),
            .lcout(\c0.rx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_10_32_0 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_10_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_10_32_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_10_32_0  (
            .in0(N__34112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_10_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_10_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_10_32_1 .LUT_INIT=16'b1011111101010101;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_10_32_1  (
            .in0(N__30720),
            .in1(N__27569),
            .in2(N__27535),
            .in3(N__30569),
            .lcout(),
            .ltout(n7415_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_10_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_10_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_10_32_2 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_10_32_2  (
            .in0(N__30659),
            .in1(N__30784),
            .in2(N__27495),
            .in3(N__28173),
            .lcout(r_SM_Main_0_adj_1736),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35424),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i7714_2_lut_LC_10_32_3 .C_ON=1'b0;
    defparam \c0.rx.i7714_2_lut_LC_10_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7714_2_lut_LC_10_32_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i7714_2_lut_LC_10_32_3  (
            .in0(_gnd_net_),
            .in1(N__30719),
            .in2(_gnd_net_),
            .in3(N__30568),
            .lcout(),
            .ltout(n9301_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_10_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_10_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_10_32_4 .LUT_INIT=16'b0000010000010101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_10_32_4  (
            .in0(N__30660),
            .in1(N__30785),
            .in2(N__27492),
            .in3(N__28089),
            .lcout(r_SM_Main_1_adj_1735),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35424),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_10_32_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_10_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_10_32_6 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_10_32_6  (
            .in0(N__28098),
            .in1(_gnd_net_),
            .in2(N__30728),
            .in3(N__28164),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i7683_3_lut_LC_10_32_7 .C_ON=1'b0;
    defparam \c0.rx.i7683_3_lut_LC_10_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7683_3_lut_LC_10_32_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.rx.i7683_3_lut_LC_10_32_7  (
            .in0(N__28165),
            .in1(N__28097),
            .in2(_gnd_net_),
            .in3(N__30715),
            .lcout(n9300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7790_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7790_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7790_LC_11_24_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7790_LC_11_24_3  (
            .in0(N__32044),
            .in1(N__28083),
            .in2(N__33150),
            .in3(N__28053),
            .lcout(),
            .ltout(\c0.n9446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9446_bdd_4_lut_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.n9446_bdd_4_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.n9446_bdd_4_lut_LC_11_24_4 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n9446_bdd_4_lut_LC_11_24_4  (
            .in0(N__28023),
            .in1(N__27993),
            .in2(N__27957),
            .in3(N__33095),
            .lcout(),
            .ltout(\c0.n9449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9728_bdd_4_lut_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.n9728_bdd_4_lut_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9728_bdd_4_lut_LC_11_24_5 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n9728_bdd_4_lut_LC_11_24_5  (
            .in0(N__27954),
            .in1(N__27804),
            .in2(N__27939),
            .in3(N__31583),
            .lcout(\c0.n9731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8024_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8024_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_8024_LC_11_25_2 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_8024_LC_11_25_2  (
            .in0(N__27931),
            .in1(N__28395),
            .in2(N__32987),
            .in3(N__31967),
            .lcout(),
            .ltout(\c0.n9740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9740_bdd_4_lut_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.n9740_bdd_4_lut_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9740_bdd_4_lut_LC_11_25_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n9740_bdd_4_lut_LC_11_25_3  (
            .in0(N__27897),
            .in1(N__32889),
            .in2(N__27858),
            .in3(N__27855),
            .lcout(),
            .ltout(\c0.n9231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_11_25_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_11_25_4  (
            .in0(N__27822),
            .in1(N__31551),
            .in2(N__27807),
            .in3(N__31193),
            .lcout(\c0.n9728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_11_25_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_11_25_5  (
            .in0(N__31552),
            .in1(N__32344),
            .in2(N__30072),
            .in3(N__30060),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(N__32271),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i145_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i145_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i145_LC_11_26_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i145_LC_11_26_1  (
            .in0(N__29841),
            .in1(N__29126),
            .in2(_gnd_net_),
            .in3(N__29157),
            .lcout(data_in_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i141_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i141_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i141_LC_11_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0___i141_LC_11_26_2  (
            .in0(N__29115),
            .in1(N__33234),
            .in2(_gnd_net_),
            .in3(N__28967),
            .lcout(data_in_field_140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_537_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_537_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_537_LC_11_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_537_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__31674),
            .in2(_gnd_net_),
            .in3(N__28396),
            .lcout(\c0.n4292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_646_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_646_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_646_LC_11_26_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_646_LC_11_26_4  (
            .in0(N__32164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33233),
            .lcout(\c0.n8957 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_688_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_688_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_688_LC_11_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_688_LC_11_26_6  (
            .in0(_gnd_net_),
            .in1(N__28301),
            .in2(_gnd_net_),
            .in3(N__28248),
            .lcout(\c0.n8871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i0_LC_11_27_0.C_ON=1'b1;
    defparam blink_counter_423__i0_LC_11_27_0.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i0_LC_11_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i0_LC_11_27_0 (
            .in0(_gnd_net_),
            .in1(N__28191),
            .in2(_gnd_net_),
            .in3(N__28185),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_11_27_0_),
            .carryout(n8130),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i1_LC_11_27_1.C_ON=1'b1;
    defparam blink_counter_423__i1_LC_11_27_1.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i1_LC_11_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i1_LC_11_27_1 (
            .in0(_gnd_net_),
            .in1(N__28182),
            .in2(_gnd_net_),
            .in3(N__28176),
            .lcout(n25_adj_1722),
            .ltout(),
            .carryin(n8130),
            .carryout(n8131),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i2_LC_11_27_2.C_ON=1'b1;
    defparam blink_counter_423__i2_LC_11_27_2.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i2_LC_11_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i2_LC_11_27_2 (
            .in0(_gnd_net_),
            .in1(N__30153),
            .in2(_gnd_net_),
            .in3(N__30147),
            .lcout(n24),
            .ltout(),
            .carryin(n8131),
            .carryout(n8132),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i3_LC_11_27_3.C_ON=1'b1;
    defparam blink_counter_423__i3_LC_11_27_3.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i3_LC_11_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i3_LC_11_27_3 (
            .in0(_gnd_net_),
            .in1(N__30144),
            .in2(_gnd_net_),
            .in3(N__30138),
            .lcout(n23),
            .ltout(),
            .carryin(n8132),
            .carryout(n8133),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i4_LC_11_27_4.C_ON=1'b1;
    defparam blink_counter_423__i4_LC_11_27_4.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i4_LC_11_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i4_LC_11_27_4 (
            .in0(_gnd_net_),
            .in1(N__30135),
            .in2(_gnd_net_),
            .in3(N__30129),
            .lcout(n22),
            .ltout(),
            .carryin(n8133),
            .carryout(n8134),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i5_LC_11_27_5.C_ON=1'b1;
    defparam blink_counter_423__i5_LC_11_27_5.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i5_LC_11_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i5_LC_11_27_5 (
            .in0(_gnd_net_),
            .in1(N__30126),
            .in2(_gnd_net_),
            .in3(N__30120),
            .lcout(n21),
            .ltout(),
            .carryin(n8134),
            .carryout(n8135),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i6_LC_11_27_6.C_ON=1'b1;
    defparam blink_counter_423__i6_LC_11_27_6.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i6_LC_11_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i6_LC_11_27_6 (
            .in0(_gnd_net_),
            .in1(N__30117),
            .in2(_gnd_net_),
            .in3(N__30111),
            .lcout(n20),
            .ltout(),
            .carryin(n8135),
            .carryout(n8136),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i7_LC_11_27_7.C_ON=1'b1;
    defparam blink_counter_423__i7_LC_11_27_7.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i7_LC_11_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i7_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(N__30108),
            .in2(_gnd_net_),
            .in3(N__30102),
            .lcout(n19),
            .ltout(),
            .carryin(n8136),
            .carryout(n8137),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i8_LC_11_28_0.C_ON=1'b1;
    defparam blink_counter_423__i8_LC_11_28_0.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i8_LC_11_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i8_LC_11_28_0 (
            .in0(_gnd_net_),
            .in1(N__30099),
            .in2(_gnd_net_),
            .in3(N__30093),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_11_28_0_),
            .carryout(n8138),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i9_LC_11_28_1.C_ON=1'b1;
    defparam blink_counter_423__i9_LC_11_28_1.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i9_LC_11_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i9_LC_11_28_1 (
            .in0(_gnd_net_),
            .in1(N__30090),
            .in2(_gnd_net_),
            .in3(N__30084),
            .lcout(n17),
            .ltout(),
            .carryin(n8138),
            .carryout(n8139),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i10_LC_11_28_2.C_ON=1'b1;
    defparam blink_counter_423__i10_LC_11_28_2.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i10_LC_11_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i10_LC_11_28_2 (
            .in0(_gnd_net_),
            .in1(N__30081),
            .in2(_gnd_net_),
            .in3(N__30075),
            .lcout(n16),
            .ltout(),
            .carryin(n8139),
            .carryout(n8140),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i11_LC_11_28_3.C_ON=1'b1;
    defparam blink_counter_423__i11_LC_11_28_3.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i11_LC_11_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i11_LC_11_28_3 (
            .in0(_gnd_net_),
            .in1(N__30225),
            .in2(_gnd_net_),
            .in3(N__30219),
            .lcout(n15),
            .ltout(),
            .carryin(n8140),
            .carryout(n8141),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i12_LC_11_28_4.C_ON=1'b1;
    defparam blink_counter_423__i12_LC_11_28_4.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i12_LC_11_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i12_LC_11_28_4 (
            .in0(_gnd_net_),
            .in1(N__30216),
            .in2(_gnd_net_),
            .in3(N__30210),
            .lcout(n14),
            .ltout(),
            .carryin(n8141),
            .carryout(n8142),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i13_LC_11_28_5.C_ON=1'b1;
    defparam blink_counter_423__i13_LC_11_28_5.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i13_LC_11_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i13_LC_11_28_5 (
            .in0(_gnd_net_),
            .in1(N__30207),
            .in2(_gnd_net_),
            .in3(N__30201),
            .lcout(n13),
            .ltout(),
            .carryin(n8142),
            .carryout(n8143),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i14_LC_11_28_6.C_ON=1'b1;
    defparam blink_counter_423__i14_LC_11_28_6.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i14_LC_11_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i14_LC_11_28_6 (
            .in0(_gnd_net_),
            .in1(N__30198),
            .in2(_gnd_net_),
            .in3(N__30192),
            .lcout(n12),
            .ltout(),
            .carryin(n8143),
            .carryout(n8144),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i15_LC_11_28_7.C_ON=1'b1;
    defparam blink_counter_423__i15_LC_11_28_7.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i15_LC_11_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i15_LC_11_28_7 (
            .in0(_gnd_net_),
            .in1(N__30189),
            .in2(_gnd_net_),
            .in3(N__30183),
            .lcout(n11),
            .ltout(),
            .carryin(n8144),
            .carryout(n8145),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i16_LC_11_29_0.C_ON=1'b1;
    defparam blink_counter_423__i16_LC_11_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i16_LC_11_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i16_LC_11_29_0 (
            .in0(_gnd_net_),
            .in1(N__30180),
            .in2(_gnd_net_),
            .in3(N__30174),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_11_29_0_),
            .carryout(n8146),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i17_LC_11_29_1.C_ON=1'b1;
    defparam blink_counter_423__i17_LC_11_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i17_LC_11_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i17_LC_11_29_1 (
            .in0(_gnd_net_),
            .in1(N__30171),
            .in2(_gnd_net_),
            .in3(N__30165),
            .lcout(n9),
            .ltout(),
            .carryin(n8146),
            .carryout(n8147),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i18_LC_11_29_2.C_ON=1'b1;
    defparam blink_counter_423__i18_LC_11_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i18_LC_11_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i18_LC_11_29_2 (
            .in0(_gnd_net_),
            .in1(N__30162),
            .in2(_gnd_net_),
            .in3(N__30156),
            .lcout(n8),
            .ltout(),
            .carryin(n8147),
            .carryout(n8148),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i19_LC_11_29_3.C_ON=1'b1;
    defparam blink_counter_423__i19_LC_11_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i19_LC_11_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i19_LC_11_29_3 (
            .in0(_gnd_net_),
            .in1(N__30378),
            .in2(_gnd_net_),
            .in3(N__30372),
            .lcout(n7),
            .ltout(),
            .carryin(n8148),
            .carryout(n8149),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i20_LC_11_29_4.C_ON=1'b1;
    defparam blink_counter_423__i20_LC_11_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i20_LC_11_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i20_LC_11_29_4 (
            .in0(_gnd_net_),
            .in1(N__30369),
            .in2(_gnd_net_),
            .in3(N__30363),
            .lcout(n6),
            .ltout(),
            .carryin(n8149),
            .carryout(n8150),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i21_LC_11_29_5.C_ON=1'b1;
    defparam blink_counter_423__i21_LC_11_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i21_LC_11_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i21_LC_11_29_5 (
            .in0(_gnd_net_),
            .in1(N__30341),
            .in2(_gnd_net_),
            .in3(N__30330),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n8150),
            .carryout(n8151),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i22_LC_11_29_6.C_ON=1'b1;
    defparam blink_counter_423__i22_LC_11_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i22_LC_11_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i22_LC_11_29_6 (
            .in0(_gnd_net_),
            .in1(N__30311),
            .in2(_gnd_net_),
            .in3(N__30300),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n8151),
            .carryout(n8152),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i23_LC_11_29_7.C_ON=1'b1;
    defparam blink_counter_423__i23_LC_11_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i23_LC_11_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i23_LC_11_29_7 (
            .in0(_gnd_net_),
            .in1(N__30284),
            .in2(_gnd_net_),
            .in3(N__30273),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n8152),
            .carryout(n8153),
            .clk(N__35414),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i24_LC_11_30_0.C_ON=1'b1;
    defparam blink_counter_423__i24_LC_11_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i24_LC_11_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i24_LC_11_30_0 (
            .in0(_gnd_net_),
            .in1(N__30260),
            .in2(_gnd_net_),
            .in3(N__30249),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_11_30_0_),
            .carryout(n8154),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_423__i25_LC_11_30_1.C_ON=1'b0;
    defparam blink_counter_423__i25_LC_11_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_423__i25_LC_11_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_423__i25_LC_11_30_1 (
            .in0(_gnd_net_),
            .in1(N__30236),
            .in2(_gnd_net_),
            .in3(N__30246),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_11_30_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_11_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_11_30_2 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_11_30_2  (
            .in0(N__30913),
            .in1(N__31076),
            .in2(N__31044),
            .in3(N__30869),
            .lcout(r_Clock_Count_6_adj_1728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_11_30_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_11_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_11_30_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_11_30_3  (
            .in0(N__30867),
            .in1(N__30911),
            .in2(N__30426),
            .in3(N__30453),
            .lcout(r_Clock_Count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_11_30_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_11_30_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_11_30_4  (
            .in0(N__30910),
            .in1(N__30868),
            .in2(N__30495),
            .in3(N__30465),
            .lcout(r_Clock_Count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam i48_4_lut_LC_11_30_5.C_ON=1'b0;
    defparam i48_4_lut_LC_11_30_5.SEQ_MODE=4'b0000;
    defparam i48_4_lut_LC_11_30_5.LUT_INIT=16'b1110111101000101;
    LogicCell40 i48_4_lut_LC_11_30_5 (
            .in0(N__30787),
            .in1(N__30738),
            .in2(N__30732),
            .in3(N__30537),
            .lcout(n44),
            .ltout(n44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_11_30_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_11_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_11_30_6 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_11_30_6  (
            .in0(N__30912),
            .in1(N__30387),
            .in2(N__30663),
            .in3(N__30414),
            .lcout(r_Clock_Count_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35419),
            .ce(),
            .sr(_gnd_net_));
    defparam i7646_2_lut_LC_11_30_7.C_ON=1'b0;
    defparam i7646_2_lut_LC_11_30_7.SEQ_MODE=4'b0000;
    defparam i7646_2_lut_LC_11_30_7.LUT_INIT=16'b1111111110101010;
    LogicCell40 i7646_2_lut_LC_11_30_7 (
            .in0(N__30642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30563),
            .lcout(n9245),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_11_31_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_11_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_11_31_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30531),
            .in3(N__30498),
            .lcout(n226),
            .ltout(),
            .carryin(bfn_11_31_0_),
            .carryout(\c0.rx.n8098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_11_31_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_11_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_11_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_3_lut_LC_11_31_1  (
            .in0(_gnd_net_),
            .in1(N__30490),
            .in2(_gnd_net_),
            .in3(N__30456),
            .lcout(n225),
            .ltout(),
            .carryin(\c0.rx.n8098 ),
            .carryout(\c0.rx.n8099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_11_31_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_11_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_11_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_4_lut_LC_11_31_2  (
            .in0(_gnd_net_),
            .in1(N__30452),
            .in2(_gnd_net_),
            .in3(N__30417),
            .lcout(n224),
            .ltout(),
            .carryin(\c0.rx.n8099 ),
            .carryout(\c0.rx.n8100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_11_31_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_11_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_11_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_5_lut_LC_11_31_3  (
            .in0(_gnd_net_),
            .in1(N__30413),
            .in2(_gnd_net_),
            .in3(N__30381),
            .lcout(n223),
            .ltout(),
            .carryin(\c0.rx.n8100 ),
            .carryout(\c0.rx.n8101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_11_31_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_11_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_11_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_6_lut_LC_11_31_4  (
            .in0(_gnd_net_),
            .in1(N__30837),
            .in2(_gnd_net_),
            .in3(N__31092),
            .lcout(n222),
            .ltout(),
            .carryin(\c0.rx.n8101 ),
            .carryout(\c0.rx.n8102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_11_31_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_11_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_11_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_7_lut_LC_11_31_5  (
            .in0(_gnd_net_),
            .in1(N__30930),
            .in2(_gnd_net_),
            .in3(N__31089),
            .lcout(n221),
            .ltout(),
            .carryin(\c0.rx.n8102 ),
            .carryout(\c0.rx.n8103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_11_31_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_11_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_11_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_8_lut_LC_11_31_6  (
            .in0(_gnd_net_),
            .in1(N__31075),
            .in2(_gnd_net_),
            .in3(N__31035),
            .lcout(n220),
            .ltout(),
            .carryin(\c0.rx.n8103 ),
            .carryout(\c0.rx.n8104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_11_31_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_11_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_11_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_9_lut_LC_11_31_7  (
            .in0(_gnd_net_),
            .in1(N__31020),
            .in2(_gnd_net_),
            .in3(N__30981),
            .lcout(n219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_505_LC_11_32_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_505_LC_11_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_505_LC_11_32_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_505_LC_11_32_4  (
            .in0(_gnd_net_),
            .in1(N__30928),
            .in2(_gnd_net_),
            .in3(N__30835),
            .lcout(n4084),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_11_32_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_11_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_11_32_5 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_11_32_5  (
            .in0(N__30929),
            .in1(N__30915),
            .in2(N__30942),
            .in3(N__30875),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35429),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_11_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_11_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_11_32_7 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_11_32_7  (
            .in0(N__30836),
            .in1(N__30914),
            .in2(N__30885),
            .in3(N__30874),
            .lcout(r_Clock_Count_4_adj_1729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35429),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9488_bdd_4_lut_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.n9488_bdd_4_lut_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.n9488_bdd_4_lut_LC_12_26_3 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n9488_bdd_4_lut_LC_12_26_3  (
            .in0(N__30822),
            .in1(N__31476),
            .in2(N__30807),
            .in3(N__31585),
            .lcout(),
            .ltout(\c0.n9491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_12_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_12_26_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_12_26_4  (
            .in0(N__31586),
            .in1(N__32403),
            .in2(N__32391),
            .in3(N__32381),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35404),
            .ce(N__32272),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7825_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7825_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_7825_LC_12_26_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_7825_LC_12_26_6  (
            .in0(N__32159),
            .in1(N__33091),
            .in2(N__32120),
            .in3(N__32043),
            .lcout(\c0.n9500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9500_bdd_4_lut_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.n9500_bdd_4_lut_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.n9500_bdd_4_lut_LC_12_27_6 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n9500_bdd_4_lut_LC_12_27_6  (
            .in0(N__33097),
            .in1(N__31732),
            .in2(N__31686),
            .in3(N__31638),
            .lcout(),
            .ltout(\c0.n9198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7835_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7835_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_7835_LC_12_27_7 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_7835_LC_12_27_7  (
            .in0(N__31389),
            .in1(N__31584),
            .in2(N__31479),
            .in3(N__31232),
            .lcout(\c0.n9488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9494_bdd_4_lut_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.n9494_bdd_4_lut_LC_12_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.n9494_bdd_4_lut_LC_12_28_2 .LUT_INIT=16'b1100111011000010;
    LogicCell40 \c0.n9494_bdd_4_lut_LC_12_28_2  (
            .in0(N__31470),
            .in1(N__31431),
            .in2(N__33210),
            .in3(N__31415),
            .lcout(\c0.n9201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_12_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_12_28_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_12_28_7  (
            .in0(N__31360),
            .in1(N__31296),
            .in2(N__31281),
            .in3(N__31259),
            .lcout(\c0.n22_adj_1677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_12_29_3.C_ON=1'b0;
    defparam i1_2_lut_LC_12_29_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_12_29_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_LC_12_29_3 (
            .in0(_gnd_net_),
            .in1(N__34031),
            .in2(_gnd_net_),
            .in3(N__33985),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_29_5 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_4_lut_LC_12_29_5 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \c0.tx.i1_3_lut_4_lut_LC_12_29_5  (
            .in0(N__33986),
            .in1(N__35638),
            .in2(N__34440),
            .in3(N__34032),
            .lcout(n5062),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_13_25_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_13_25_4  (
            .in0(N__34351),
            .in1(N__33673),
            .in2(N__35814),
            .in3(N__33420),
            .lcout(\c0.byte_transmit_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35405),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_2_lut_LC_13_26_0 .C_ON=1'b1;
    defparam \c0.add_2248_2_lut_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_2_lut_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_2_lut_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__33849),
            .in2(N__33836),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_6_7_N_965_0 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\c0.n8083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_3_lut_LC_13_26_1 .C_ON=1'b1;
    defparam \c0.add_2248_3_lut_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_3_lut_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_3_lut_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__33896),
            .in2(_gnd_net_),
            .in3(N__32424),
            .lcout(\c0.data_out_6_7_N_965_1 ),
            .ltout(),
            .carryin(\c0.n8083 ),
            .carryout(\c0.n8084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_4_lut_LC_13_26_2 .C_ON=1'b1;
    defparam \c0.add_2248_4_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_4_lut_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_4_lut_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__33700),
            .in2(_gnd_net_),
            .in3(N__32421),
            .lcout(\c0.data_out_6_7_N_965_2 ),
            .ltout(),
            .carryin(\c0.n8084 ),
            .carryout(\c0.n8085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_5_lut_LC_13_26_3 .C_ON=1'b1;
    defparam \c0.add_2248_5_lut_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_5_lut_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_5_lut_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__33660),
            .in2(_gnd_net_),
            .in3(N__32418),
            .lcout(\c0.data_out_6_7_N_965_3 ),
            .ltout(),
            .carryin(\c0.n8085 ),
            .carryout(\c0.n8086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_6_lut_LC_13_26_4 .C_ON=1'b1;
    defparam \c0.add_2248_6_lut_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_6_lut_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_6_lut_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__33758),
            .in2(_gnd_net_),
            .in3(N__32415),
            .lcout(\c0.data_out_6_7_N_965_4 ),
            .ltout(),
            .carryin(\c0.n8086 ),
            .carryout(\c0.n8087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_7_lut_LC_13_26_5 .C_ON=1'b1;
    defparam \c0.add_2248_7_lut_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_7_lut_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_7_lut_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__33494),
            .in2(_gnd_net_),
            .in3(N__32412),
            .lcout(data_out_6_7_N_965_5),
            .ltout(),
            .carryin(\c0.n8087 ),
            .carryout(\c0.n8088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_8_lut_LC_13_26_6 .C_ON=1'b1;
    defparam \c0.add_2248_8_lut_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_8_lut_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_8_lut_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__33443),
            .in2(_gnd_net_),
            .in3(N__32409),
            .lcout(\c0.data_out_6_7_N_965_6 ),
            .ltout(),
            .carryin(\c0.n8088 ),
            .carryout(\c0.n8089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2248_9_lut_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.add_2248_9_lut_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2248_9_lut_LC_13_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2248_9_lut_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__33431),
            .in2(_gnd_net_),
            .in3(N__32406),
            .lcout(\c0.data_out_6_7_N_965_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_740_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_740_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_740_LC_13_27_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i1_2_lut_adj_740_LC_13_27_1  (
            .in0(N__33780),
            .in1(N__33675),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n11 ),
            .ltout(\c0.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_691_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_691_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_691_LC_13_27_2 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \c0.i2_4_lut_adj_691_LC_13_27_2  (
            .in0(N__33821),
            .in1(N__33727),
            .in2(N__32619),
            .in3(N__33910),
            .lcout(tx_data_0_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_692_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_692_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_692_LC_13_27_3 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_692_LC_13_27_3  (
            .in0(N__33911),
            .in1(N__33375),
            .in2(N__33842),
            .in3(N__33861),
            .lcout(),
            .ltout(tx_data_3_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_13_27_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_13_27_4  (
            .in0(N__34207),
            .in1(_gnd_net_),
            .in2(N__32616),
            .in3(N__33632),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35415),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_13_27_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_13_27_7  (
            .in0(N__33779),
            .in1(N__33674),
            .in2(_gnd_net_),
            .in3(N__33820),
            .lcout(\c0.n45_adj_1656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_13_28_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_13_28_0  (
            .in0(N__32613),
            .in1(N__34218),
            .in2(_gnd_net_),
            .in3(N__34079),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35420),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7754_4_lut_LC_13_28_1 .C_ON=1'b0;
    defparam \c0.i7754_4_lut_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7754_4_lut_LC_13_28_1 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \c0.i7754_4_lut_LC_13_28_1  (
            .in0(N__33918),
            .in1(N__33724),
            .in2(N__33379),
            .in3(N__33837),
            .lcout(tx_data_7_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_564_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_564_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_564_LC_13_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_564_LC_13_28_2  (
            .in0(N__32607),
            .in1(N__32556),
            .in2(_gnd_net_),
            .in3(N__32507),
            .lcout(\c0.n8986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_696_LC_13_28_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_696_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_696_LC_13_28_3 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \c0.i1_3_lut_adj_696_LC_13_28_3  (
            .in0(N__33917),
            .in1(N__32430),
            .in2(_gnd_net_),
            .in3(N__33725),
            .lcout(tx_data_6_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_4_lut_4_lut_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_4_lut_4_lut_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_4_lut_4_lut_LC_13_28_5 .LUT_INIT=16'b0000000100001010;
    LogicCell40 \c0.i1_4_lut_4_lut_4_lut_LC_13_28_5  (
            .in0(N__33919),
            .in1(N__33726),
            .in2(N__33380),
            .in3(N__33838),
            .lcout(),
            .ltout(tx_data_5_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_28_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(N__34219),
            .in2(N__33384),
            .in3(N__33584),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35420),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_13_29_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_13_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_13_29_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_13_29_0  (
            .in0(N__33843),
            .in1(N__33920),
            .in2(N__33735),
            .in3(N__33381),
            .lcout(),
            .ltout(tx_data_2_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_13_29_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_29_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_13_29_1  (
            .in0(N__33330),
            .in1(_gnd_net_),
            .in2(N__33351),
            .in3(N__34220),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35425),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_13_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_13_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_13_29_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_13_29_3  (
            .in0(N__33348),
            .in1(N__34221),
            .in2(_gnd_net_),
            .in3(N__33339),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35425),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_13_29_4.C_ON=1'b0;
    defparam i13_4_lut_LC_13_29_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_13_29_4.LUT_INIT=16'b0001110000010000;
    LogicCell40 i13_4_lut_LC_13_29_4 (
            .in0(N__34003),
            .in1(N__35631),
            .in2(N__34568),
            .in3(N__34439),
            .lcout(),
            .ltout(n8705_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_13_29_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_13_29_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_13_29_5  (
            .in0(N__35632),
            .in1(_gnd_net_),
            .in2(N__33342),
            .in3(N__34044),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35425),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_7994_LC_13_29_6.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_7994_LC_13_29_6.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_7994_LC_13_29_6.LUT_INIT=16'b1010111111000000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_7994_LC_13_29_6 (
            .in0(N__33338),
            .in1(N__33329),
            .in2(N__33987),
            .in3(N__35630),
            .lcout(n9452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_13_29_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_13_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_13_29_7 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_13_29_7  (
            .in0(N__34034),
            .in1(N__34004),
            .in2(_gnd_net_),
            .in3(N__34043),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35425),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n9680_bdd_4_lut_LC_13_31_5 .C_ON=1'b0;
    defparam \c0.n9680_bdd_4_lut_LC_13_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.n9680_bdd_4_lut_LC_13_31_5 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n9680_bdd_4_lut_LC_13_31_5  (
            .in0(N__33321),
            .in1(N__33273),
            .in2(N__33261),
            .in3(N__33096),
            .lcout(\c0.n9683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.i6_3_lut_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_LC_14_25_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i6_3_lut_LC_14_25_0  (
            .in0(N__34983),
            .in1(N__35850),
            .in2(_gnd_net_),
            .in3(N__34917),
            .lcout(),
            .ltout(\c0.n17_adj_1663_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_671_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_671_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_671_LC_14_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_671_LC_14_25_1  (
            .in0(N__34125),
            .in1(N__34230),
            .in2(N__33453),
            .in3(N__33927),
            .lcout(\c0.n123 ),
            .ltout(\c0.n123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_14_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_14_25_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_14_25_2  (
            .in0(N__35785),
            .in1(N__33770),
            .in2(N__33450),
            .in3(N__33543),
            .lcout(\c0.byte_transmit_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_14_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_14_25_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_14_25_4  (
            .in0(N__33473),
            .in1(N__33719),
            .in2(N__35813),
            .in3(N__33408),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_14_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_14_25_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_14_25_5  (
            .in0(N__34348),
            .in1(N__35786),
            .in2(N__33447),
            .in3(N__33555),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_14_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_14_25_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_14_25_6  (
            .in0(N__33432),
            .in1(N__34349),
            .in2(N__35812),
            .in3(N__33531),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i1_LC_14_25_7 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_14_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_14_25_7 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.UART_TRANSMITTER_state__i1_LC_14_25_7  (
            .in0(N__34350),
            .in1(N__35784),
            .in2(_gnd_net_),
            .in3(N__34283),
            .lcout(UART_TRANSMITTER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_14_26_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \c0.i2_4_lut_LC_14_26_0  (
            .in0(N__33419),
            .in1(N__33482),
            .in2(N__33396),
            .in3(N__33407),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i0_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_14_26_1 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_14_26_1  (
            .in0(N__33469),
            .in1(N__33395),
            .in2(N__35815),
            .in3(N__33835),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35416),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_672_LC_14_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_672_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_672_LC_14_26_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_672_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__33506),
            .in2(_gnd_net_),
            .in3(N__33554),
            .lcout(),
            .ltout(\c0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_673_LC_14_26_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_673_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_673_LC_14_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_673_LC_14_26_3  (
            .in0(N__33542),
            .in1(N__33530),
            .in2(N__33519),
            .in3(N__33516),
            .lcout(\c0.n7814 ),
            .ltout(\c0.n7814_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_674_LC_14_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_674_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_674_LC_14_26_4 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \c0.i1_2_lut_adj_674_LC_14_26_4  (
            .in0(N__34347),
            .in1(_gnd_net_),
            .in2(N__33510),
            .in3(_gnd_net_),
            .lcout(n7204),
            .ltout(n7204_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_14_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_14_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_14_26_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_14_26_5  (
            .in0(N__33507),
            .in1(N__35817),
            .in2(N__33498),
            .in3(N__33495),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35416),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_1995_LC_14_26_6 .C_ON=1'b0;
    defparam \c0.tx_transmit_1995_LC_14_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_1995_LC_14_26_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx_transmit_1995_LC_14_26_6  (
            .in0(N__34547),
            .in1(N__34284),
            .in2(N__35827),
            .in3(N__34158),
            .lcout(\c0.tx_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35416),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_14_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i1_LC_14_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_14_26_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_14_26_7  (
            .in0(N__33483),
            .in1(N__35816),
            .in2(N__33474),
            .in3(N__33913),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35416),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7750_3_lut_4_lut_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.i7750_3_lut_4_lut_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7750_3_lut_4_lut_LC_14_27_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.i7750_3_lut_4_lut_LC_14_27_0  (
            .in0(N__33677),
            .in1(N__33723),
            .in2(N__33921),
            .in3(N__33777),
            .lcout(tx_data_1_N_keep),
            .ltout(tx_data_1_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_14_27_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_14_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_14_27_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__34195),
            .in2(N__33456),
            .in3(N__33599),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35421),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_14_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_14_27_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_663_LC_14_27_2  (
            .in0(N__33676),
            .in1(N__33823),
            .in2(_gnd_net_),
            .in3(N__33776),
            .lcout(),
            .ltout(\c0.n7779_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_693_LC_14_27_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_693_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_693_LC_14_27_3 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \c0.i1_4_lut_adj_693_LC_14_27_3  (
            .in0(N__33912),
            .in1(N__33639),
            .in2(N__33864),
            .in3(N__33860),
            .lcout(tx_data_4_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_737_LC_14_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_737_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_737_LC_14_27_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_737_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__34167),
            .in2(_gnd_net_),
            .in3(N__34153),
            .lcout(\c0.data_out_6__7__N_973 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7693_2_lut_3_lut_4_lut_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.i7693_2_lut_3_lut_4_lut_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7693_2_lut_3_lut_4_lut_LC_14_27_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i7693_2_lut_3_lut_4_lut_LC_14_27_5  (
            .in0(N__33822),
            .in1(N__33778),
            .in2(N__33731),
            .in3(N__33678),
            .lcout(\c0.n9291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_LC_14_27_6.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_LC_14_27_6.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_LC_14_27_6.LUT_INIT=16'b1111010110001000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_LC_14_27_6 (
            .in0(N__33984),
            .in1(N__33633),
            .in2(N__33612),
            .in3(N__35645),
            .lcout(n9710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_14_27_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_14_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_14_27_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_14_27_7  (
            .in0(N__33618),
            .in1(N__34196),
            .in2(_gnd_net_),
            .in3(N__33611),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35421),
            .ce(),
            .sr(_gnd_net_));
    defparam n9710_bdd_4_lut_LC_14_28_1.C_ON=1'b0;
    defparam n9710_bdd_4_lut_LC_14_28_1.SEQ_MODE=4'b0000;
    defparam n9710_bdd_4_lut_LC_14_28_1.LUT_INIT=16'b1111101001000100;
    LogicCell40 n9710_bdd_4_lut_LC_14_28_1 (
            .in0(N__33973),
            .in1(N__33600),
            .in2(N__33585),
            .in3(N__33570),
            .lcout(),
            .ltout(n9713_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i591325_i1_3_lut_LC_14_28_2.C_ON=1'b0;
    defparam i591325_i1_3_lut_LC_14_28_2.SEQ_MODE=4'b0000;
    defparam i591325_i1_3_lut_LC_14_28_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 i591325_i1_3_lut_LC_14_28_2 (
            .in0(N__34033),
            .in1(_gnd_net_),
            .in2(N__33564),
            .in3(N__34065),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_14_28_3 .LUT_INIT=16'b1111110000110011;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_14_28_3  (
            .in0(_gnd_net_),
            .in1(N__34501),
            .in2(N__33561),
            .in3(N__34427),
            .lcout(),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_14_28_4 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_14_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_14_28_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_14_28_4  (
            .in0(_gnd_net_),
            .in1(N__34097),
            .in2(N__33558),
            .in3(N__35538),
            .lcout(tx_o_adj_1726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35426),
            .ce(),
            .sr(_gnd_net_));
    defparam n9452_bdd_4_lut_LC_14_28_6.C_ON=1'b0;
    defparam n9452_bdd_4_lut_LC_14_28_6.SEQ_MODE=4'b0000;
    defparam n9452_bdd_4_lut_LC_14_28_6.LUT_INIT=16'b1010101011011000;
    LogicCell40 n9452_bdd_4_lut_LC_14_28_6 (
            .in0(N__34086),
            .in1(N__34052),
            .in2(N__34080),
            .in3(N__33972),
            .lcout(n9455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_14_28_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_14_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_14_28_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_14_28_7  (
            .in0(N__34053),
            .in1(N__34200),
            .in2(_gnd_net_),
            .in3(N__34059),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35426),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7402_4_lut_LC_14_29_2 .C_ON=1'b0;
    defparam \c0.tx.i7402_4_lut_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7402_4_lut_LC_14_29_2 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \c0.tx.i7402_4_lut_LC_14_29_2  (
            .in0(N__35536),
            .in1(N__35745),
            .in2(N__34500),
            .in3(N__34423),
            .lcout(n9073),
            .ltout(n9073_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_14_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_14_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_14_29_3 .LUT_INIT=16'b1111000100000010;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_14_29_3  (
            .in0(N__34035),
            .in1(N__34008),
            .in2(N__33990),
            .in3(N__33980),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35430),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_14_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_14_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_14_29_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_14_29_4  (
            .in0(N__35537),
            .in1(N__34658),
            .in2(_gnd_net_),
            .in3(N__34638),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35430),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Done_44_LC_14_30_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Done_44_LC_14_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Done_44_LC_14_30_0 .LUT_INIT=16'b1111010111101100;
    LogicCell40 \c0.tx.r_Tx_Done_44_LC_14_30_0  (
            .in0(N__34512),
            .in1(N__34359),
            .in2(N__33936),
            .in3(N__35553),
            .lcout(n3892),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35432),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_669_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_669_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_669_LC_15_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_669_LC_15_25_0  (
            .in0(N__34719),
            .in1(N__34892),
            .in2(N__34854),
            .in3(N__34679),
            .lcout(\c0.n18_adj_1662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5731_2_lut_3_lut_LC_15_25_1 .C_ON=1'b0;
    defparam \c0.i5731_2_lut_3_lut_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5731_2_lut_3_lut_LC_15_25_1 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i5731_2_lut_3_lut_LC_15_25_1  (
            .in0(N__34680),
            .in1(N__34339),
            .in2(_gnd_net_),
            .in3(N__34279),
            .lcout(\c0.n20_adj_1652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5736_2_lut_3_lut_LC_15_25_2 .C_ON=1'b0;
    defparam \c0.i5736_2_lut_3_lut_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5736_2_lut_3_lut_LC_15_25_2 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \c0.i5736_2_lut_3_lut_LC_15_25_2  (
            .in0(N__34282),
            .in1(_gnd_net_),
            .in2(N__34353),
            .in3(N__34893),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5730_2_lut_3_lut_LC_15_25_3 .C_ON=1'b0;
    defparam \c0.i5730_2_lut_3_lut_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5730_2_lut_3_lut_LC_15_25_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i5730_2_lut_3_lut_LC_15_25_3  (
            .in0(N__34698),
            .in1(N__34338),
            .in2(_gnd_net_),
            .in3(N__34278),
            .lcout(\c0.n21_adj_1653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5733_2_lut_3_lut_LC_15_25_4 .C_ON=1'b0;
    defparam \c0.i5733_2_lut_3_lut_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5733_2_lut_3_lut_LC_15_25_4 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \c0.i5733_2_lut_3_lut_LC_15_25_4  (
            .in0(N__34281),
            .in1(_gnd_net_),
            .in2(N__34352),
            .in3(N__34958),
            .lcout(\c0.n18_adj_1650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_670_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_670_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_670_LC_15_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_adj_670_LC_15_25_5  (
            .in0(N__34697),
            .in1(N__34937),
            .in2(N__34959),
            .in3(N__34874),
            .lcout(\c0.n19_adj_1664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5732_2_lut_3_lut_LC_15_25_7 .C_ON=1'b0;
    defparam \c0.i5732_2_lut_3_lut_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5732_2_lut_3_lut_LC_15_25_7 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i5732_2_lut_3_lut_LC_15_25_7  (
            .in0(N__34982),
            .in1(N__34340),
            .in2(_gnd_net_),
            .in3(N__34280),
            .lcout(\c0.n19_adj_1651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5667_2_lut_3_lut_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.i5667_2_lut_3_lut_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5667_2_lut_3_lut_LC_15_26_0 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.i5667_2_lut_3_lut_LC_15_26_0  (
            .in0(N__34272),
            .in1(N__34718),
            .in2(_gnd_net_),
            .in3(N__34332),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_675_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_675_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_675_LC_15_26_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i2_3_lut_adj_675_LC_15_26_1  (
            .in0(N__34543),
            .in1(N__34271),
            .in2(_gnd_net_),
            .in3(N__34157),
            .lcout(\c0.n900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5734_2_lut_3_lut_LC_15_26_2 .C_ON=1'b0;
    defparam \c0.i5734_2_lut_3_lut_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5734_2_lut_3_lut_LC_15_26_2 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.i5734_2_lut_3_lut_LC_15_26_2  (
            .in0(N__34273),
            .in1(N__34938),
            .in2(_gnd_net_),
            .in3(N__34333),
            .lcout(\c0.n17_adj_1649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5738_2_lut_3_lut_LC_15_26_3 .C_ON=1'b0;
    defparam \c0.i5738_2_lut_3_lut_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5738_2_lut_3_lut_LC_15_26_3 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.i5738_2_lut_3_lut_LC_15_26_3  (
            .in0(N__34336),
            .in1(N__34853),
            .in2(_gnd_net_),
            .in3(N__34276),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5739_2_lut_3_lut_LC_15_26_4 .C_ON=1'b0;
    defparam \c0.i5739_2_lut_3_lut_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5739_2_lut_3_lut_LC_15_26_4 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.i5739_2_lut_3_lut_LC_15_26_4  (
            .in0(N__34277),
            .in1(N__35846),
            .in2(_gnd_net_),
            .in3(N__34337),
            .lcout(\c0.n12_adj_1634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5737_2_lut_3_lut_LC_15_26_5 .C_ON=1'b0;
    defparam \c0.i5737_2_lut_3_lut_LC_15_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5737_2_lut_3_lut_LC_15_26_5 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.i5737_2_lut_3_lut_LC_15_26_5  (
            .in0(N__34335),
            .in1(N__34875),
            .in2(_gnd_net_),
            .in3(N__34275),
            .lcout(\c0.n14_adj_1639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5735_2_lut_3_lut_LC_15_26_7 .C_ON=1'b0;
    defparam \c0.i5735_2_lut_3_lut_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5735_2_lut_3_lut_LC_15_26_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.i5735_2_lut_3_lut_LC_15_26_7  (
            .in0(N__34334),
            .in1(N__34916),
            .in2(_gnd_net_),
            .in3(N__34274),
            .lcout(\c0.n16_adj_1641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_668_LC_15_27_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_668_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_668_LC_15_27_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_668_LC_15_27_0  (
            .in0(_gnd_net_),
            .in1(N__34540),
            .in2(_gnd_net_),
            .in3(N__34154),
            .lcout(\c0.n117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_15_27_2 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_15_27_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_4_lut_LC_15_27_2  (
            .in0(N__35534),
            .in1(N__34419),
            .in2(N__34502),
            .in3(N__34541),
            .lcout(n3747),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_1994_LC_15_27_3 .C_ON=1'b0;
    defparam \c0.tx_active_prev_1994_LC_15_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_1994_LC_15_27_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.tx_active_prev_1994_LC_15_27_3  (
            .in0(N__34156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35427),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7727_3_lut_4_lut_4_lut_LC_15_27_4 .C_ON=1'b0;
    defparam \c0.tx.i7727_3_lut_4_lut_4_lut_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7727_3_lut_4_lut_4_lut_LC_15_27_4 .LUT_INIT=16'b1000001110000000;
    LogicCell40 \c0.tx.i7727_3_lut_4_lut_4_lut_LC_15_27_4  (
            .in0(N__35735),
            .in1(N__34420),
            .in2(N__34503),
            .in3(N__34542),
            .lcout(),
            .ltout(n8749_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_15_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_15_27_5 .LUT_INIT=16'b1000101010111010;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_15_27_5  (
            .in0(N__34155),
            .in1(N__35535),
            .in2(N__34161),
            .in3(N__34428),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35427),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7389_2_lut_3_lut_LC_15_28_0 .C_ON=1'b0;
    defparam \c0.tx.i7389_2_lut_3_lut_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7389_2_lut_3_lut_LC_15_28_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.tx.i7389_2_lut_3_lut_LC_15_28_0  (
            .in0(N__35710),
            .in1(N__34410),
            .in2(_gnd_net_),
            .in3(N__35513),
            .lcout(\c0.tx.n9059 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_3_lut_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_3_lut_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_3_lut_LC_15_28_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \c0.tx.i1_2_lut_3_lut_LC_15_28_1  (
            .in0(N__35512),
            .in1(_gnd_net_),
            .in2(N__34429),
            .in3(N__35709),
            .lcout(),
            .ltout(\c0.tx.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_509_LC_15_28_2 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_509_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_509_LC_15_28_2 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \c0.tx.i1_4_lut_adj_509_LC_15_28_2  (
            .in0(N__35683),
            .in1(N__34479),
            .in2(N__34128),
            .in3(N__34578),
            .lcout(\c0.tx.n9027 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_15_28_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_15_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_15_28_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_15_28_3  (
            .in0(N__35516),
            .in1(N__35736),
            .in2(N__34499),
            .in3(N__34426),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35431),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_15_28_4 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_15_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_15_28_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_15_28_4  (
            .in0(N__34425),
            .in1(N__34484),
            .in2(N__35744),
            .in3(N__35515),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35431),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i6328_4_lut_LC_15_28_5 .C_ON=1'b0;
    defparam \c0.tx.i6328_4_lut_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i6328_4_lut_LC_15_28_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.tx.i6328_4_lut_LC_15_28_5  (
            .in0(N__35610),
            .in1(N__34424),
            .in2(N__34572),
            .in3(N__34548),
            .lcout(),
            .ltout(n3151_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_15_28_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_15_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_15_28_6 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_15_28_6  (
            .in0(N__35737),
            .in1(N__34483),
            .in2(N__34515),
            .in3(N__35514),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35431),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_747_LC_15_29_0.C_ON=1'b0;
    defparam i1_2_lut_adj_747_LC_15_29_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_747_LC_15_29_0.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_747_LC_15_29_0 (
            .in0(N__34421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34486),
            .lcout(n11_adj_1752),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_15_29_1 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_15_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_15_29_1 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx.i1_4_lut_LC_15_29_1  (
            .in0(N__34627),
            .in1(N__35572),
            .in2(N__34659),
            .in3(N__34603),
            .lcout(),
            .ltout(\c0.tx.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_508_LC_15_29_2 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_508_LC_15_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_508_LC_15_29_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx.i1_4_lut_adj_508_LC_15_29_2  (
            .in0(N__35596),
            .in1(N__34825),
            .in2(N__34506),
            .in3(N__35452),
            .lcout(\c0.tx.n23 ),
            .ltout(\c0.tx.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7651_2_lut_3_lut_4_lut_LC_15_29_3 .C_ON=1'b0;
    defparam \c0.tx.i7651_2_lut_3_lut_4_lut_LC_15_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7651_2_lut_3_lut_4_lut_LC_15_29_3 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \c0.tx.i7651_2_lut_3_lut_4_lut_LC_15_29_3  (
            .in0(N__34485),
            .in1(N__35689),
            .in2(N__34443),
            .in3(N__34422),
            .lcout(n9259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_15_29_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_15_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_15_29_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_15_29_4  (
            .in0(N__34604),
            .in1(_gnd_net_),
            .in2(N__35556),
            .in3(N__34590),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_15_29_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_15_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_15_29_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_15_29_5  (
            .in0(N__34826),
            .in1(N__35550),
            .in2(_gnd_net_),
            .in3(N__34812),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_510_LC_15_29_6 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_510_LC_15_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_510_LC_15_29_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.tx.i1_2_lut_adj_510_LC_15_29_6  (
            .in0(N__35545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34668),
            .lcout(\c0.tx.n7916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_15_29_7  (
            .in0(N__34628),
            .in1(N__35546),
            .in2(_gnd_net_),
            .in3(N__34614),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35433),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_15_30_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_15_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_15_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_2_lut_LC_15_30_0  (
            .in0(N__34792),
            .in1(N__34751),
            .in2(_gnd_net_),
            .in3(N__34662),
            .lcout(n9249),
            .ltout(),
            .carryin(bfn_15_30_0_),
            .carryout(\c0.tx.n8090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_15_30_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_15_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_15_30_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_3_lut_LC_15_30_1  (
            .in0(N__34796),
            .in1(N__34657),
            .in2(_gnd_net_),
            .in3(N__34632),
            .lcout(\c0.tx.n9290 ),
            .ltout(),
            .carryin(\c0.tx.n8090 ),
            .carryout(\c0.tx.n8091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_15_30_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_15_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_15_30_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_4_lut_LC_15_30_2  (
            .in0(N__34793),
            .in1(N__34629),
            .in2(_gnd_net_),
            .in3(N__34608),
            .lcout(\c0.tx.n9313 ),
            .ltout(),
            .carryin(\c0.tx.n8091 ),
            .carryout(\c0.tx.n8092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_15_30_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_15_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_15_30_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_5_lut_LC_15_30_3  (
            .in0(N__34797),
            .in1(N__34605),
            .in2(_gnd_net_),
            .in3(N__34584),
            .lcout(\c0.tx.n9281 ),
            .ltout(),
            .carryin(\c0.tx.n8092 ),
            .carryout(\c0.tx.n8093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_15_30_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_15_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_15_30_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_6_lut_LC_15_30_4  (
            .in0(N__34794),
            .in1(N__35597),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(n9305),
            .ltout(),
            .carryin(\c0.tx.n8093 ),
            .carryout(\c0.tx.n8094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_15_30_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_15_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_15_30_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_7_lut_LC_15_30_5  (
            .in0(N__34798),
            .in1(N__35573),
            .in2(_gnd_net_),
            .in3(N__34830),
            .lcout(\c0.tx.n9314 ),
            .ltout(),
            .carryin(\c0.tx.n8094 ),
            .carryout(\c0.tx.n8095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_15_30_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_15_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_15_30_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_8_lut_LC_15_30_6  (
            .in0(N__34795),
            .in1(N__34827),
            .in2(_gnd_net_),
            .in3(N__34806),
            .lcout(n9304),
            .ltout(),
            .carryin(\c0.tx.n8095 ),
            .carryout(\c0.tx.n8096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_15_30_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_15_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_15_30_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_9_lut_LC_15_30_7  (
            .in0(N__34799),
            .in1(N__35453),
            .in2(_gnd_net_),
            .in3(N__34803),
            .lcout(n9303),
            .ltout(),
            .carryin(\c0.tx.n8096 ),
            .carryout(\c0.tx.n8097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_15_31_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_15_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_15_31_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_10_lut_LC_15_31_0  (
            .in0(N__34800),
            .in1(N__35681),
            .in2(_gnd_net_),
            .in3(N__34761),
            .lcout(n9266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_15_31_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_15_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_15_31_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_15_31_2  (
            .in0(N__34758),
            .in1(N__34752),
            .in2(_gnd_net_),
            .in3(N__35551),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35435),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_15_31_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_15_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_15_31_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_15_31_6  (
            .in0(N__35682),
            .in1(N__35552),
            .in2(_gnd_net_),
            .in3(N__34740),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35435),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i0_LC_16_25_0 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i0_LC_16_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i0_LC_16_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i0_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__34734),
            .in2(N__34728),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\c0.n8120 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i1_LC_16_25_1 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i1_LC_16_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i1_LC_16_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i1_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__34704),
            .in2(_gnd_net_),
            .in3(N__34689),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n8120 ),
            .carryout(\c0.n8121 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i2_LC_16_25_2 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i2_LC_16_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i2_LC_16_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i2_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__34686),
            .in2(_gnd_net_),
            .in3(N__34671),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n8121 ),
            .carryout(\c0.n8122 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i3_LC_16_25_3 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i3_LC_16_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i3_LC_16_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i3_LC_16_25_3  (
            .in0(_gnd_net_),
            .in1(N__34989),
            .in2(_gnd_net_),
            .in3(N__34968),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n8122 ),
            .carryout(\c0.n8123 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i4_LC_16_25_4 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i4_LC_16_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i4_LC_16_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i4_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(N__34965),
            .in2(_gnd_net_),
            .in3(N__34947),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n8123 ),
            .carryout(\c0.n8124 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i5_LC_16_25_5 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i5_LC_16_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i5_LC_16_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i5_LC_16_25_5  (
            .in0(_gnd_net_),
            .in1(N__34944),
            .in2(_gnd_net_),
            .in3(N__34926),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n8124 ),
            .carryout(\c0.n8125 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i6_LC_16_25_6 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i6_LC_16_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i6_LC_16_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i6_LC_16_25_6  (
            .in0(_gnd_net_),
            .in1(N__34923),
            .in2(_gnd_net_),
            .in3(N__34902),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n8125 ),
            .carryout(\c0.n8126 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i7_LC_16_25_7 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i7_LC_16_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i7_LC_16_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i7_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__34899),
            .in2(_gnd_net_),
            .in3(N__34884),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(\c0.n8126 ),
            .carryout(\c0.n8127 ),
            .clk(N__35422),
            .ce(N__35832),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i8_LC_16_26_0 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i8_LC_16_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i8_LC_16_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i8_LC_16_26_0  (
            .in0(_gnd_net_),
            .in1(N__34881),
            .in2(_gnd_net_),
            .in3(N__34863),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_16_26_0_),
            .carryout(\c0.n8128 ),
            .clk(N__35428),
            .ce(N__35831),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i9_LC_16_26_1 .C_ON=1'b1;
    defparam \c0.delay_counter_424__i9_LC_16_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i9_LC_16_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i9_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__34860),
            .in2(_gnd_net_),
            .in3(N__34839),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(\c0.n8128 ),
            .carryout(\c0.n8129 ),
            .clk(N__35428),
            .ce(N__35831),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_424__i10_LC_16_26_2 .C_ON=1'b0;
    defparam \c0.delay_counter_424__i10_LC_16_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_424__i10_LC_16_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_424__i10_LC_16_26_2  (
            .in0(_gnd_net_),
            .in1(N__34836),
            .in2(_gnd_net_),
            .in3(N__35853),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35428),
            .ce(N__35831),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_16_28_5 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_16_28_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_16_28_5  (
            .in0(_gnd_net_),
            .in1(N__35690),
            .in2(_gnd_net_),
            .in3(N__35711),
            .lcout(r_SM_Main_2_N_1480_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7696_2_lut_3_lut_LC_16_28_6 .C_ON=1'b0;
    defparam \c0.tx.i7696_2_lut_3_lut_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7696_2_lut_3_lut_LC_16_28_6 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \c0.tx.i7696_2_lut_3_lut_LC_16_28_6  (
            .in0(N__35712),
            .in1(_gnd_net_),
            .in2(N__35694),
            .in3(N__35649),
            .lcout(\c0.tx.n9310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_16_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_16_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_16_29_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_16_29_3  (
            .in0(N__35539),
            .in1(N__35598),
            .in2(_gnd_net_),
            .in3(N__35604),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35434),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_16_30_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_16_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_16_30_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_16_30_1  (
            .in0(N__35554),
            .in1(N__35574),
            .in2(_gnd_net_),
            .in3(N__35580),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35436),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_16_30_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_16_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_16_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_16_30_5  (
            .in0(N__35555),
            .in1(N__35454),
            .in2(_gnd_net_),
            .in3(N__35460),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35436),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
