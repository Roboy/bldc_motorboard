// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Sep 12 18:02:55 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    inout PIN_1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    inout PIN_2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    input PIN_12 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    input PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    input PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    input PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire GND_net, VCC_net, LED_c, tx_o, tx2_o, tx_enable, tx2_enable, 
        rx_i;
    wire [25:0]blink_counter;   // verilog/TinyFPGA_B.v(64[14:27])
    
    wire n16346, n16466;
    wire [31:0]rand_data;   // verilog/TinyFPGA_B.v(77[14:23])
    wire [31:0]rand_setpoint;   // verilog/TinyFPGA_B.v(78[14:27])
    
    wire n9390, n10351;
    wire [7:0]byte_transmit_counter;   // coms.v(19[11:32])
    
    wire n10419, n157, n19, n165, n10471, n10420, n10418, n10421, 
        n10358, n164;
    wire [7:0]\data_out[8] ;   // coms.v(21[11:19])
    
    wire n14;
    wire [7:0]\data_out[3] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    
    wire n163;
    wire [14:0]delay_counter;   // coms.v(266[12:25])
    wire [7:0]\UART_TRANSMITTER.state ;   // coms.v(271[13:18])
    
    wire rx_data_ready;
    wire [7:0]rx_data;   // coms.v(378[13:20])
    wire [7:0]\data_in[20] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[19] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[18] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[17] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[16] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[15] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[14] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[13] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[12] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[11] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[10] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[9] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[8] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[7] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[6] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[5] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[4] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[3] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[2] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[1] ;   // coms.v(382[12:19])
    wire [7:0]\data_in[0] ;   // coms.v(382[12:19])
    
    wire n6878;
    wire [7:0]\data_in_frame[10] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[9] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[8] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[7] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[6] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[5] ;   // coms.v(383[12:25])
    wire [7:0]\data_in_frame[1] ;   // coms.v(383[12:25])
    wire [7:0]\data_out_frame2[19] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[18] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[17] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[16] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[15] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[14] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[13] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[12] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[11] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[10] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[9] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[8] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[7] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[6] ;   // coms.v(384[12:27])
    wire [7:0]\data_out_frame2[5] ;   // coms.v(384[12:27])
    
    wire n10625, n10628, n10631, n10632, n10633, n10634, n10635, 
        n10636, n10637, n10638, n7080, n7086;
    wire [31:0]\FRAME_MATCHER.next_state ;   // coms.v(423[11:21])
    
    wire n162, n4980, n10510, n10502, n161, n10509, n10508, data_out_6__6__N_729, 
        n10347, data_out_6__7__N_678, n159, n160, n63, data_out_5__4__N_959, 
        n16998, n116, data_out_5__7__N_931, n15;
    wire [7:0]tx_transmit_N_2239;
    
    wire n17312, n10346, n159_adj_2580, n158, n157_adj_2581, n156, 
        n155, n154, n153, n152, n151, n150, n149, n148, n147, 
        n146, n145, n144, n143, n142, n141, n140, n139, n138, 
        n137, n118, n136, n135, n134, n10415, n16345, n16344, 
        n16326, n16343, n16420, n10245, n16419, n17028, n16418, 
        n16417, n16325, n11, n9796, n9135, n10244, n16416, n16415, 
        n16342, n16341, n13601, n16324, n16414, n16413, n13597, 
        n8, n10474, n9, n4, n16412, n1, n4_adj_2582, n10432, 
        n111;
    wire [7:0]\UART_TRANSMITTER.state_7__N_1749 ;
    
    wire n10483, n133, n6, n16340, n10427, data_out_6__1__N_850, 
        data_out_6__2__N_804, n128, n10426, n10475, n6_adj_2583, n114;
    wire [7:0]i_Tx_Byte;   // verilog/uart_tx.v(18[16:25])
    
    wire tx_active, tx_o_adj_2584, n29, n125, n132, n115, n121, 
        n47, n10416, data_out_10__7__N_114, n13880, n10476, n16864, 
        n10477, n135_adj_2585, n130, n17548, n10194, n131, n17080, 
        n127, n126, n16323, n12123, n17030, n155_adj_2586, n165_adj_2587, 
        n164_adj_2588, n163_adj_2589, n152_adj_2590, n154_adj_2591, 
        n161_adj_2592, n16, n10, n146_adj_2593, n149_adj_2594, n153_adj_2595, 
        n156_adj_2596, n140_adj_2597, n136_adj_2598, n143_adj_2599, 
        n10170, n26, n162_adj_2600, n135_adj_2601, n134_adj_2602, 
        n10166, n139_adj_2603, n6_adj_2604, n16339, n16322, n10597, 
        n16338, n10414, n2560, n2561, n2562, n2563, n2564, n2565, 
        n2566, n2567, n2568, n2570, n2571, n2572, n2573, n2574, 
        n2575, n10488, n10489, n10490, n10491, n10494, n10500, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2593, n2594, n2595, n2596, n2597, n2598, n2599, n10516, 
        n10518, n10519, n10520, n10523, n10525, n10529, n10563, 
        n10564, n10565, n10566, n10567, n10568, n10569, n10570, 
        n10571, n10572, n10573, n10574, n10575, n10576, n10577, 
        n10578, n10579, n10580, n10581, n10582, n10583, n10584, 
        n10585, n10586, n10587, n10588, n10589, n10590, n10591, 
        n10592, n10593, n16321;
    wire [31:0]\FRAME_MATCHER.next_state_31__N_2026 ;
    
    wire n8529, n8_adj_2605, n121_adj_2606, n41, n17356, n119, n96, 
        n16337, n16336, n16335, n17767, n17757, n17856, n10594, 
        n16320, n16404, n16334, n9054, n9100, n17681, n9051, n16403, 
        n16402, n16401, n10160, n17547, n17092, n17737, n17082, 
        n17084, n17366, n160_adj_2607, n8517, n158_adj_2608, n151_adj_2609, 
        n16400, n16333, n10484, n21, n24, n25, n16399, n10428, 
        n10429, n10430, n10431, n10481, n16332, n112, n142_adj_2610, 
        n10603, n10602, n10601, n10600, n10599, n10598, n16398, 
        n16397, n16396, n16395, n16394, n16393, n16392, n16391, 
        n16390, n16442, n17078, n16389, n16441, n16440, n16388, 
        n16439, n17709, n10702, n16485, n16468, n10691, n10683, 
        n10671, n10662, n10659, n10655, n16438, n10652, n10649, 
        n10646, n10645, n10644, n10643, n9652, n9646, n8_adj_2611, 
        n16437, n9631, n16436, n10144, n10142, n10141, n10140, 
        n10139, n10137, n10135, n18104, n10134, n10133, n10132, 
        n10130, n10129, n10128, n10127, n10126, n10604, n18103, 
        n4_adj_2612, n18102, n113, n10125, n18101, n9606, n10124, 
        n10123, n10121, n10119, n10118, n10116, n10114, n10112, 
        n10110, n10109, n10108, n18098, n10106, n18097, n10105, 
        n17054, n10104, n10102, n10101, n16387, n9519, n10100, 
        n16331, n10099, n10095, n10092, n8_adj_2613, n10089, n1396, 
        n134_adj_2614, n10086, n10083, n16386, n16435, n14_adj_2615, 
        n16385, n16434, n9419, n10407, n10353, n9283, n6_adj_2616, 
        n17306, n10364, n10366, n10367, n10369, n10370, n10371, 
        n10372, n10374, n10375, n10377, n10378, n10379, n10380, 
        n10382, n10383, n10385, n10386, n10387, n10044, n10043, 
        n17364, n17585, n16968, n3, n16330, n10360, n16384, n7734, 
        n17481, n9148, n17479, n10357, n8562, n17672, n9380, n10039, 
        n2615, n16433, n10038, n12, n10487, n18054, n8_adj_2617, 
        n16954, n10485, n10034, n4958, n10562, n10561, n4430, 
        n2720, n10033, n10032, n10031, n18032, n13, n16329, n10473, 
        n10505, n10501, n10027, n117, n10026, n10025, n10024, 
        n16432, n10499, n10497, n16383, n18465, n10405, n10404, 
        n10403, n10495, n10478, n10402, n10401, n10400, n10023, 
        n10022, n10560, n16319, n10559, n10558, n10557, n10556, 
        n10555, n10554, n10553, n10552, n10551, n10550, n10549, 
        n10548, n10547, n12_adj_2618, n10546, n18462, n10545, n10544, 
        n10543, n10021, n10542, n10541, n7364;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n16382, n16431, n18010;
    wire [2:0]r_SM_Main_2__N_2323;
    
    wire n16430, n16429, n43, n10019, n10018, n10017, n10016, 
        n22, n16428, r_Rx_Data;
    wire [7:0]r_Clock_Count_adj_2660;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index_adj_2661;   // verilog/uart_rx.v(33[17:28])
    
    wire n10504, n10398, n10399, n10540, n10539, n10538, n10326, 
        n38, n10396, n16427, n221, n222, n223, n224, n225, n226, 
        n10009, n10008, n10005, n10004, n10003, n10002;
    wire [2:0]r_SM_Main_adj_2665;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_2666;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_2667;   // verilog/uart_tx.v(33[16:27])
    
    wire n16426, n10395, n10394, n10393, n9999, n9996, n9993, 
        n9992, n10391, n316, n317, n318, n319, n320, n321, n10537, 
        n10536, n16425, n10535, n10534, n10533, n138_adj_2638, n10532, 
        n10325, n10531, n10438, n10388, n10439, n16381, n10530, 
        n10440, n16380, n9989, n9988, n123, n9987, n9986, n148_adj_2639, 
        n9985, n141_adj_2640, n137_adj_2641, n16424, n120, n9983, 
        n13415, n9982, n18441, n9981, n9980, n17480, n9979, n10506, 
        n17958, n10324, n23, n16932, n8567, n9978, n63_adj_2642, 
        n20, n10472, n144_adj_2643, n150_adj_2644, n17952, n145_adj_2645, 
        n17950, n9977, n147_adj_2646, n10469, n10468, n10467, n10466, 
        n10465, n10464, n10463, n10462, n10461, n10460, n10459, 
        n10458, n10457, n10456, n10455, n10454, n10453, n10452, 
        n10451, n10450, n10449, n10448, n10447, n10446, n10445, 
        n10444, n10443, n10442, n10441, n10528, n18438, n9976, 
        n129, n9972, n110, n124, n8_adj_2647, n10417, n119_adj_2648, 
        n10389, n10352, n17, n10527, n10526, n10507, n10425, n10363, 
        n10524, n10437, n10424, n10436, n10435, n10434, n10423, 
        n10433, n4_adj_2649, n10422, n10323, n10410, n10596, n10411, 
        n10412, n10515, n16423, n10413, n10517, n10595, n3_adj_2650, 
        n10521, n10522, n17855, n16328, n10482, n10406, n10486, 
        n10408, n10492, n10409, n10493, n16327, n10359, n10361, 
        n16422, n19_adj_2651, n9938, n9937, n9935, n10479, n10480, 
        n16421, n13_adj_2652, n10511, n9922, n4_adj_2653, n10397, 
        n10390, n8_adj_2654, n18, n10470, n122, n8488, n10496, 
        n10503, n22_adj_2655, n7, n10498, n10513, n9920, n10512, 
        n9947, n16_adj_2656, n9942, n10514, n16349, n9941, n9940, 
        n9934, n9933, n9932, n16348, n16347;
    
    VCC i2 (.Y(VCC_net));
    SB_IO tx2_output (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx2_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx2_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx2_output.PIN_TYPE = 6'b101001;
    defparam tx2_output.PULLUP = 1'b1;
    defparam tx2_output.NEG_TRIGGER = 1'b0;
    defparam tx2_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO rx_input (.PACKAGE_PIN(PIN_2), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(rx_i)) /* synthesis lattice_noprune=1, syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam rx_input.PIN_TYPE = 6'b000001;
    defparam rx_input.PULLUP = 1'b1;
    defparam rx_input.NEG_TRIGGER = 1'b0;
    defparam rx_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_1), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rand_data_2269_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[20]), 
            .I3(n16338), .O(n145_adj_2645)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33_3_lut (.I0(n18102), .I1(r_Clock_Count[2]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17082));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_22 (.CI(n16338), .I0(GND_net), .I1(rand_data[20]), 
            .CO(n16339));
    SB_CARRY rand_data_2269_add_4_8 (.CI(n16324), .I0(GND_net), .I1(rand_data[6]), 
            .CO(n16325));
    SB_DFF rand_data_2269__i0 (.Q(rand_data[0]), .C(CLK_c), .D(n165_adj_2587));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8143_3_lut (.I0(\data_out_frame2[13] [3]), .I1(rand_data[27]), 
            .I2(n9606), .I3(GND_net), .O(n10559));   // coms.v(428[12] 532[6])
    defparam i8143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8005_3_lut (.I0(\data_in[12] [1]), .I1(\data_in[13] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10421));   // coms.v(402[9] 410[5])
    defparam i8005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8006_3_lut (.I0(\data_in[12] [2]), .I1(\data_in[13] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10422));   // coms.v(402[9] 410[5])
    defparam i8006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8144_3_lut (.I0(\data_out_frame2[13] [4]), .I1(rand_data[28]), 
            .I2(n9606), .I3(GND_net), .O(n10560));   // coms.v(428[12] 532[6])
    defparam i8144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[6]), .I3(r_Bit_Index[1]), .O(n18462));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18462_bdd_4_lut (.I0(n18462), .I1(r_Tx_Data[4]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n18465));
    defparam n18462_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rand_data_2269_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[5]), 
            .I3(n16323), .O(n160_adj_2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8145_3_lut (.I0(\data_out_frame2[13] [5]), .I1(rand_data[29]), 
            .I2(n9606), .I3(GND_net), .O(n10561));   // coms.v(428[12] 532[6])
    defparam i8145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8146_3_lut (.I0(\data_out_frame2[13] [6]), .I1(rand_data[30]), 
            .I2(n9606), .I3(GND_net), .O(n10562));   // coms.v(428[12] 532[6])
    defparam i8146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8147_3_lut (.I0(\data_out_frame2[13] [7]), .I1(rand_data[31]), 
            .I2(n9606), .I3(GND_net), .O(n10563));   // coms.v(428[12] 532[6])
    defparam i8147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8007_3_lut (.I0(\data_in[12] [3]), .I1(\data_in[13] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10423));   // coms.v(402[9] 410[5])
    defparam i8007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8148_3_lut (.I0(\data_out_frame2[14] [0]), .I1(rand_data[16]), 
            .I2(n9606), .I3(GND_net), .O(n10564));   // coms.v(428[12] 532[6])
    defparam i8148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8149_3_lut (.I0(\data_out_frame2[14] [1]), .I1(rand_data[17]), 
            .I2(n9606), .I3(GND_net), .O(n10565));   // coms.v(428[12] 532[6])
    defparam i8149_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_15 (.CI(n16392), .I0(GND_net), .I1(n13), 
            .CO(n16393));
    SB_CARRY rand_data_2269_add_4_7 (.CI(n16323), .I0(GND_net), .I1(rand_data[5]), 
            .CO(n16324));
    SB_LUT4 rand_data_2269_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[4]), 
            .I3(n16322), .O(n161_adj_2592)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2271_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n16391), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8150_3_lut (.I0(\data_out_frame2[14] [2]), .I1(rand_data[18]), 
            .I2(n9606), .I3(GND_net), .O(n10566));   // coms.v(428[12] 532[6])
    defparam i8150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[19]), 
            .I3(n16337), .O(n146_adj_2593)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_14 (.CI(n16391), .I0(GND_net), .I1(n14), 
            .CO(n16392));
    SB_LUT4 i8151_3_lut (.I0(\data_out_frame2[14] [3]), .I1(rand_data[19]), 
            .I2(n9606), .I3(GND_net), .O(n10567));   // coms.v(428[12] 532[6])
    defparam i8151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2604));   // coms.v(383[12:25])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8152_3_lut (.I0(\data_out_frame2[14] [4]), .I1(rand_data[20]), 
            .I2(n9606), .I3(GND_net), .O(n10568));   // coms.v(428[12] 532[6])
    defparam i8152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[7] [0]), .I1(n9054), .I2(n9380), 
            .I3(n6_adj_2604), .O(n17547));   // coms.v(383[12:25])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n17547), .I1(n9051), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n17548));   // coms.v(383[12:25])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 blink_counter_2271_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n16390), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8153_3_lut (.I0(\data_out_frame2[14] [5]), .I1(rand_data[21]), 
            .I2(n9606), .I3(GND_net), .O(n10569));   // coms.v(428[12] 532[6])
    defparam i8153_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_13 (.CI(n16390), .I0(GND_net), .I1(n15), 
            .CO(n16391));
    SB_LUT4 i8154_3_lut (.I0(\data_out_frame2[14] [6]), .I1(rand_data[22]), 
            .I2(n9606), .I3(GND_net), .O(n10570));   // coms.v(428[12] 532[6])
    defparam i8154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8008_3_lut (.I0(\data_in[12] [4]), .I1(\data_in[13] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10424));   // coms.v(402[9] 410[5])
    defparam i8008_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_21 (.CI(n16337), .I0(GND_net), .I1(rand_data[19]), 
            .CO(n16338));
    SB_LUT4 i8009_3_lut (.I0(\data_in[12] [5]), .I1(\data_in[13] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10425));   // coms.v(402[9] 410[5])
    defparam i8009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17479));   // coms.v(383[12:25])
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(n17479), .I1(n6_adj_2583), .I2(\data_in_frame[9] [6]), 
            .I3(n9051), .O(n17480));   // coms.v(383[12:25])
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i8010_3_lut (.I0(\data_in[12] [6]), .I1(\data_in[13] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10426));   // coms.v(402[9] 410[5])
    defparam i8010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2271_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n16389), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_12 (.CI(n16389), .I0(GND_net), .I1(n16), 
            .CO(n16390));
    SB_LUT4 i8011_3_lut (.I0(\data_in[12] [7]), .I1(\data_in[13] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10427));   // coms.v(402[9] 410[5])
    defparam i8011_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_6 (.CI(n16322), .I0(GND_net), .I1(rand_data[4]), 
            .CO(n16323));
    SB_LUT4 i8012_3_lut (.I0(\data_in[13] [0]), .I1(\data_in[14] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10428));   // coms.v(402[9] 410[5])
    defparam i8012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8013_3_lut (.I0(\data_in[13] [1]), .I1(\data_in[14] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10429));   // coms.v(402[9] 410[5])
    defparam i8013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[18]), 
            .I3(n16336), .O(n147_adj_2646)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_2651));   // coms.v(383[12:25])
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i7973_3_lut (.I0(\data_in[8] [1]), .I1(\data_in[9] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10389));   // coms.v(402[9] 410[5])
    defparam i7973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8155_3_lut (.I0(\data_out_frame2[14] [7]), .I1(rand_data[23]), 
            .I2(n9606), .I3(GND_net), .O(n10571));   // coms.v(428[12] 532[6])
    defparam i8155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut_15992 (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[3]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n18438));
    defparam r_Bit_Index_2__bdd_4_lut_15992.LUT_INIT = 16'he4aa;
    SB_LUT4 blink_counter_2271_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n16388), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n18438_bdd_4_lut (.I0(n18438), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[1]), 
            .I3(r_Bit_Index[1]), .O(n18441));
    defparam n18438_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8156_3_lut (.I0(\data_out_frame2[15] [0]), .I1(rand_data[8]), 
            .I2(n9606), .I3(GND_net), .O(n10572));   // coms.v(428[12] 532[6])
    defparam i8156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[3]), 
            .I3(n16321), .O(n162_adj_2600)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_5 (.CI(n16321), .I0(GND_net), .I1(rand_data[3]), 
            .CO(n16322));
    SB_CARRY blink_counter_2271_add_4_11 (.CI(n16388), .I0(GND_net), .I1(n17), 
            .CO(n16389));
    SB_LUT4 blink_counter_2271_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n16387), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8157_3_lut (.I0(\data_out_frame2[15] [1]), .I1(rand_data[9]), 
            .I2(n9606), .I3(GND_net), .O(n10573));   // coms.v(428[12] 532[6])
    defparam i8157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8014_3_lut (.I0(\data_in[13] [2]), .I1(\data_in[14] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10430));   // coms.v(402[9] 410[5])
    defparam i8014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8015_3_lut (.I0(\data_in[13] [3]), .I1(\data_in[14] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10431));   // coms.v(402[9] 410[5])
    defparam i8015_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_10 (.CI(n16387), .I0(GND_net), .I1(n18), 
            .CO(n16388));
    SB_LUT4 i8016_3_lut (.I0(\data_in[13] [4]), .I1(\data_in[14] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10432));   // coms.v(402[9] 410[5])
    defparam i8016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2271_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n16386), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_20 (.CI(n16336), .I0(GND_net), .I1(rand_data[18]), 
            .CO(n16337));
    SB_LUT4 rand_data_2269_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[2]), 
            .I3(n16320), .O(n163_adj_2589)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7974_3_lut (.I0(\data_in[8] [2]), .I1(\data_in[9] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10390));   // coms.v(402[9] 410[5])
    defparam i7974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8158_3_lut (.I0(\data_out_frame2[15] [2]), .I1(rand_data[10]), 
            .I2(n9606), .I3(GND_net), .O(n10574));   // coms.v(428[12] 532[6])
    defparam i8158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8159_3_lut (.I0(\data_out_frame2[15] [3]), .I1(rand_data[11]), 
            .I2(n9606), .I3(GND_net), .O(n10575));   // coms.v(428[12] 532[6])
    defparam i8159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8160_3_lut (.I0(\data_out_frame2[15] [4]), .I1(rand_data[12]), 
            .I2(n9606), .I3(GND_net), .O(n10576));   // coms.v(428[12] 532[6])
    defparam i8160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8161_3_lut (.I0(\data_out_frame2[15] [5]), .I1(rand_data[13]), 
            .I2(n9606), .I3(GND_net), .O(n10577));   // coms.v(428[12] 532[6])
    defparam i8161_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_9 (.CI(n16386), .I0(GND_net), .I1(n19), 
            .CO(n16387));
    SB_LUT4 rand_data_2269_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[17]), 
            .I3(n16335), .O(n148_adj_2639)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2271_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n16385), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8162_3_lut (.I0(\data_out_frame2[15] [6]), .I1(rand_data[14]), 
            .I2(n9606), .I3(GND_net), .O(n10578));   // coms.v(428[12] 532[6])
    defparam i8162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8163_3_lut (.I0(\data_out_frame2[15] [7]), .I1(rand_data[15]), 
            .I2(n9606), .I3(GND_net), .O(n10579));   // coms.v(428[12] 532[6])
    defparam i8163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8164_3_lut (.I0(\data_out_frame2[16] [0]), .I1(rand_data[0]), 
            .I2(n9606), .I3(GND_net), .O(n10580));   // coms.v(428[12] 532[6])
    defparam i8164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8165_3_lut (.I0(\data_out_frame2[16] [1]), .I1(rand_data[1]), 
            .I2(n9606), .I3(GND_net), .O(n10581));   // coms.v(428[12] 532[6])
    defparam i8165_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_4 (.CI(n16320), .I0(GND_net), .I1(rand_data[2]), 
            .CO(n16321));
    SB_CARRY blink_counter_2271_add_4_8 (.CI(n16385), .I0(GND_net), .I1(n20), 
            .CO(n16386));
    SB_LUT4 i8166_3_lut (.I0(\data_out_frame2[16] [2]), .I1(rand_data[2]), 
            .I2(n9606), .I3(GND_net), .O(n10582));   // coms.v(428[12] 532[6])
    defparam i8166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8167_3_lut (.I0(\data_out_frame2[16] [3]), .I1(rand_data[3]), 
            .I2(n9606), .I3(GND_net), .O(n10583));   // coms.v(428[12] 532[6])
    defparam i8167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8168_3_lut (.I0(\data_out_frame2[16] [4]), .I1(rand_data[4]), 
            .I2(n9606), .I3(GND_net), .O(n10584));   // coms.v(428[12] 532[6])
    defparam i8168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2271_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n16384), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_19 (.CI(n16335), .I0(GND_net), .I1(rand_data[17]), 
            .CO(n16336));
    SB_LUT4 i8169_3_lut (.I0(\data_out_frame2[16] [5]), .I1(rand_data[5]), 
            .I2(n9606), .I3(GND_net), .O(n10585));   // coms.v(428[12] 532[6])
    defparam i8169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8170_3_lut (.I0(\data_out_frame2[16] [6]), .I1(rand_data[6]), 
            .I2(n9606), .I3(GND_net), .O(n10586));   // coms.v(428[12] 532[6])
    defparam i8170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8171_3_lut (.I0(\data_out_frame2[16] [7]), .I1(rand_data[7]), 
            .I2(n9606), .I3(GND_net), .O(n10587));   // coms.v(428[12] 532[6])
    defparam i8171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8218_3_lut (.I0(r_Tx_Data[3]), .I1(i_Tx_Byte[3]), .I2(n7734), 
            .I3(GND_net), .O(n10634));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8219_3_lut (.I0(r_Tx_Data[4]), .I1(i_Tx_Byte[4]), .I2(n7734), 
            .I3(GND_net), .O(n10635));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8172_3_lut (.I0(\data_out_frame2[17] [0]), .I1(rand_data[8]), 
            .I2(n9606), .I3(GND_net), .O(n10588));   // coms.v(428[12] 532[6])
    defparam i8172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8173_3_lut (.I0(\data_out_frame2[17] [1]), .I1(rand_data[9]), 
            .I2(n9606), .I3(GND_net), .O(n10589));   // coms.v(428[12] 532[6])
    defparam i8173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8174_3_lut (.I0(\data_out_frame2[17] [2]), .I1(rand_data[10]), 
            .I2(n9606), .I3(GND_net), .O(n10590));   // coms.v(428[12] 532[6])
    defparam i8174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8055_3_lut (.I0(\data_in[18] [3]), .I1(\data_in[19] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10471));   // coms.v(402[9] 410[5])
    defparam i8055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8175_3_lut (.I0(\data_out_frame2[17] [3]), .I1(rand_data[11]), 
            .I2(n9606), .I3(GND_net), .O(n10591));   // coms.v(428[12] 532[6])
    defparam i8175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8176_3_lut (.I0(\data_out_frame2[17] [4]), .I1(rand_data[12]), 
            .I2(n9606), .I3(GND_net), .O(n10592));   // coms.v(428[12] 532[6])
    defparam i8176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8177_3_lut (.I0(\data_out_frame2[17] [5]), .I1(rand_data[13]), 
            .I2(n9606), .I3(GND_net), .O(n10593));   // coms.v(428[12] 532[6])
    defparam i8177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8017_3_lut (.I0(\data_in[13] [5]), .I1(\data_in[14] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10433));   // coms.v(402[9] 410[5])
    defparam i8017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8018_3_lut (.I0(\data_in[13] [6]), .I1(\data_in[14] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10434));   // coms.v(402[9] 410[5])
    defparam i8018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8019_3_lut (.I0(\data_in[13] [7]), .I1(\data_in[14] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10435));   // coms.v(402[9] 410[5])
    defparam i8019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8020_3_lut (.I0(\data_in[14] [0]), .I1(\data_in[15] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10436));   // coms.v(402[9] 410[5])
    defparam i8020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8220_3_lut (.I0(r_Tx_Data[5]), .I1(i_Tx_Byte[5]), .I2(n7734), 
            .I3(GND_net), .O(n10636));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8056_3_lut (.I0(\data_in[18] [4]), .I1(\data_in[19] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10472));   // coms.v(402[9] 410[5])
    defparam i8056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8021_3_lut (.I0(\data_in[14] [1]), .I1(\data_in[15] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10437));   // coms.v(402[9] 410[5])
    defparam i8021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8022_3_lut (.I0(\data_in[14] [2]), .I1(\data_in[15] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10438));   // coms.v(402[9] 410[5])
    defparam i8022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8057_3_lut (.I0(\data_in[18] [5]), .I1(\data_in[19] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10473));   // coms.v(402[9] 410[5])
    defparam i8057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7975_3_lut (.I0(\data_in[8] [3]), .I1(\data_in[9] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10391));   // coms.v(402[9] 410[5])
    defparam i7975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7951_3_lut (.I0(\data_in[5] [3]), .I1(\data_in[6] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10367));   // coms.v(402[9] 410[5])
    defparam i7951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8178_3_lut (.I0(\data_out_frame2[17] [6]), .I1(rand_data[14]), 
            .I2(n9606), .I3(GND_net), .O(n10594));   // coms.v(428[12] 532[6])
    defparam i8178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut_adj_1132 (.I0(n18101), .I1(r_Clock_Count[1]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17084));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_1132.LUT_INIT = 16'hcaca;
    SB_LUT4 i8221_3_lut (.I0(r_Tx_Data[6]), .I1(i_Tx_Byte[6]), .I2(n7734), 
            .I3(GND_net), .O(n10637));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8179_3_lut (.I0(\data_out_frame2[17] [7]), .I1(rand_data[15]), 
            .I2(n9606), .I3(GND_net), .O(n10595));   // coms.v(428[12] 532[6])
    defparam i8179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8180_3_lut (.I0(\data_out_frame2[18] [0]), .I1(rand_data[0]), 
            .I2(n9606), .I3(GND_net), .O(n10596));   // coms.v(428[12] 532[6])
    defparam i8180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[1]), 
            .I3(n16319), .O(n164_adj_2588)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_7 (.CI(n16384), .I0(GND_net), .I1(n21), 
            .CO(n16385));
    SB_LUT4 i7972_3_lut (.I0(\data_in[8] [0]), .I1(\data_in[9] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10388));   // coms.v(402[9] 410[5])
    defparam i7972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[16]), 
            .I3(n16334), .O(n149_adj_2594)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8230_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_2582), 
            .I3(n8567), .O(n10646));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8230_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7953_3_lut (.I0(\data_in[5] [5]), .I1(\data_in[6] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10369));   // coms.v(402[9] 410[5])
    defparam i7953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2271_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_2655), .I3(n16383), .O(n131)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_6 (.CI(n16383), .I0(GND_net), .I1(n22_adj_2655), 
            .CO(n16384));
    SB_LUT4 i8058_3_lut (.I0(\data_in[18] [6]), .I1(\data_in[19] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10474));   // coms.v(402[9] 410[5])
    defparam i8058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8059_3_lut (.I0(\data_in[18] [7]), .I1(\data_in[19] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10475));   // coms.v(402[9] 410[5])
    defparam i8059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8229_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n13597), 
            .I3(n8562), .O(n10645));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8229_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i8060_3_lut (.I0(\data_in[19] [0]), .I1(\data_in[20] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10476));   // coms.v(402[9] 410[5])
    defparam i8060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8061_3_lut (.I0(\data_in[19] [1]), .I1(\data_in[20] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10477));   // coms.v(402[9] 410[5])
    defparam i8061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7954_3_lut (.I0(\data_in[5] [6]), .I1(\data_in[6] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10370));   // coms.v(402[9] 410[5])
    defparam i7954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2271_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23), .I3(n16382), .O(n132)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8228_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n13597), 
            .I3(n8567), .O(n10644));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8228_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i8062_3_lut (.I0(\data_in[19] [2]), .I1(\data_in[20] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10478));   // coms.v(402[9] 410[5])
    defparam i8062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8063_3_lut (.I0(\data_in[19] [3]), .I1(\data_in[20] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10479));   // coms.v(402[9] 410[5])
    defparam i8063_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_5 (.CI(n16382), .I0(GND_net), .I1(n23), 
            .CO(n16383));
    SB_LUT4 i7955_3_lut (.I0(\data_in[5] [7]), .I1(\data_in[6] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10371));   // coms.v(402[9] 410[5])
    defparam i7955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10787_3_lut (.I0(\data_in[6] [0]), .I1(\data_in[7] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10372));   // coms.v(377[7:20])
    defparam i10787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8227_4_lut (.I0(n9920), .I1(r_Bit_Index_adj_2661[1]), .I2(r_Bit_Index_adj_2661[0]), 
            .I3(n9646), .O(n10643));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8227_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i8064_3_lut (.I0(\data_in[19] [4]), .I1(\data_in[20] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10480));   // coms.v(402[9] 410[5])
    defparam i8064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7958_3_lut (.I0(\data_in[6] [2]), .I1(\data_in[7] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10374));   // coms.v(402[9] 410[5])
    defparam i7958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8065_3_lut (.I0(\data_in[19] [5]), .I1(\data_in[20] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10481));   // coms.v(402[9] 410[5])
    defparam i8065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8066_3_lut (.I0(\data_in[19] [6]), .I1(\data_in[20] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10482));   // coms.v(402[9] 410[5])
    defparam i8066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8067_3_lut (.I0(\data_in[19] [7]), .I1(\data_in[20] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10483));   // coms.v(402[9] 410[5])
    defparam i8067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8068_3_lut (.I0(\data_in[20] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10484));   // coms.v(402[9] 410[5])
    defparam i8068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8069_3_lut (.I0(\data_in[20] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10485));   // coms.v(402[9] 410[5])
    defparam i8069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_4_lut (.I0(byte_transmit_counter[5]), .I1(tx_transmit_N_2239[5]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8_adj_2611));   // coms.v(274[12] 374[6])
    defparam i25_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8070_3_lut (.I0(\data_in[20] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10486));   // coms.v(402[9] 410[5])
    defparam i8070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8071_3_lut (.I0(\data_in[20] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10487));   // coms.v(402[9] 410[5])
    defparam i8071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_4_lut_adj_1133 (.I0(byte_transmit_counter[4]), .I1(tx_transmit_N_2239[4]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8_adj_2654));   // coms.v(274[12] 374[6])
    defparam i25_4_lut_adj_1133.LUT_INIT = 16'h0aca;
    SB_CARRY rand_data_2269_add_4_3 (.CI(n16319), .I0(GND_net), .I1(rand_data[1]), 
            .CO(n16320));
    SB_LUT4 i8072_3_lut (.I0(\data_in[20] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10488));   // coms.v(402[9] 410[5])
    defparam i8072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7959_3_lut (.I0(\data_in[6] [3]), .I1(\data_in[7] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10375));   // coms.v(402[9] 410[5])
    defparam i7959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_4_lut_adj_1134 (.I0(byte_transmit_counter[3]), .I1(tx_transmit_N_2239[3]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8_adj_2605));   // coms.v(274[12] 374[6])
    defparam i25_4_lut_adj_1134.LUT_INIT = 16'h0aca;
    SB_LUT4 i8073_3_lut (.I0(\data_in[20] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10489));   // coms.v(402[9] 410[5])
    defparam i8073_3_lut.LUT_INIT = 16'hcaca;
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rand_data_2269_add_4_18 (.CI(n16334), .I0(GND_net), .I1(rand_data[16]), 
            .CO(n16335));
    SB_LUT4 rand_setpoint_2270_add_4_33_lut (.I0(GND_net), .I1(rand_data[31]), 
            .I2(rand_setpoint[31]), .I3(n16442), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25_4_lut_adj_1135 (.I0(byte_transmit_counter[2]), .I1(tx_transmit_N_2239[2]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8_adj_2647));   // coms.v(274[12] 374[6])
    defparam i25_4_lut_adj_1135.LUT_INIT = 16'h0aca;
    SB_LUT4 i8074_3_lut (.I0(\data_in[20] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10490));   // coms.v(402[9] 410[5])
    defparam i8074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9716_4_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(n17757), 
            .I3(n9796), .O(n12123));
    defparam i9716_4_lut.LUT_INIT = 16'ha6a0;
    SB_LUT4 i8075_3_lut (.I0(\data_in[20] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10491));   // coms.v(402[9] 410[5])
    defparam i8075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[15]), 
            .I3(n16333), .O(n150_adj_2644)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9717_4_lut (.I0(n17767), .I1(n12123), .I2(r_Bit_Index[0]), 
            .I3(r_Bit_Index[2]), .O(n10702));   // verilog/uart_tx.v(33[16:27])
    defparam i9717_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i8076_3_lut (.I0(\data_out_frame2[5] [0]), .I1(rand_data[24]), 
            .I2(n9606), .I3(GND_net), .O(n10492));   // coms.v(428[12] 532[6])
    defparam i8076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8077_3_lut (.I0(\data_out_frame2[5] [1]), .I1(rand_data[25]), 
            .I2(n9606), .I3(GND_net), .O(n10493));   // coms.v(428[12] 532[6])
    defparam i8077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8078_3_lut (.I0(\data_out_frame2[5] [2]), .I1(rand_data[26]), 
            .I2(n9606), .I3(GND_net), .O(n10494));   // coms.v(428[12] 532[6])
    defparam i8078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8079_3_lut (.I0(\data_out_frame2[5] [3]), .I1(rand_data[27]), 
            .I2(n9606), .I3(GND_net), .O(n10495));   // coms.v(428[12] 532[6])
    defparam i8079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_32_lut (.I0(GND_net), .I1(rand_data[30]), 
            .I2(rand_setpoint[30]), .I3(n16441), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8080_3_lut (.I0(\data_out_frame2[5] [4]), .I1(rand_data[28]), 
            .I2(n9606), .I3(GND_net), .O(n10496));   // coms.v(428[12] 532[6])
    defparam i8080_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_32 (.CI(n16441), .I0(rand_data[30]), 
            .I1(rand_setpoint[30]), .CO(n16442));
    SB_CARRY rand_data_2269_add_4_17 (.CI(n16333), .I0(GND_net), .I1(rand_data[15]), 
            .CO(n16334));
    SB_LUT4 i15317_2_lut (.I0(n17757), .I1(n9796), .I2(GND_net), .I3(GND_net), 
            .O(n17767));
    defparam i15317_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8081_3_lut (.I0(\data_out_frame2[5] [5]), .I1(rand_data[29]), 
            .I2(n9606), .I3(GND_net), .O(n10497));   // coms.v(428[12] 532[6])
    defparam i8081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8082_3_lut (.I0(\data_out_frame2[5] [6]), .I1(rand_data[30]), 
            .I2(n9606), .I3(GND_net), .O(n10498));   // coms.v(428[12] 532[6])
    defparam i8082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8083_3_lut (.I0(\data_out_frame2[5] [7]), .I1(rand_data[31]), 
            .I2(n9606), .I3(GND_net), .O(n10499));   // coms.v(428[12] 532[6])
    defparam i8083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8084_3_lut (.I0(\data_out_frame2[6] [0]), .I1(rand_data[16]), 
            .I2(n9606), .I3(GND_net), .O(n10500));   // coms.v(428[12] 532[6])
    defparam i8084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_31_lut (.I0(GND_net), .I1(rand_data[29]), 
            .I2(rand_setpoint[29]), .I3(n16440), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8085_3_lut (.I0(\data_out_frame2[6] [1]), .I1(rand_data[17]), 
            .I2(n9606), .I3(GND_net), .O(n10501));   // coms.v(428[12] 532[6])
    defparam i8085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8086_3_lut (.I0(\data_out_frame2[6] [2]), .I1(rand_data[18]), 
            .I2(n9606), .I3(GND_net), .O(n10502));   // coms.v(428[12] 532[6])
    defparam i8086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7683_3_lut (.I0(\data_in[4] [2]), .I1(\data_in[5] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10099));   // coms.v(402[9] 410[5])
    defparam i7683_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_31 (.CI(n16440), .I0(rand_data[29]), 
            .I1(rand_setpoint[29]), .CO(n16441));
    SB_LUT4 rand_setpoint_2270_add_4_30_lut (.I0(GND_net), .I1(rand_data[28]), 
            .I2(rand_setpoint[28]), .I3(n16439), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_30 (.CI(n16439), .I0(rand_data[28]), 
            .I1(rand_setpoint[28]), .CO(n16440));
    SB_LUT4 blink_counter_2271_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n16381), .O(n133)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2269_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[14]), 
            .I3(n16332), .O(n151_adj_2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7945_3_lut (.I0(\data_out[8] [0]), .I1(rand_setpoint[0]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10361));   // coms.v(274[12] 374[6])
    defparam i7945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_29_lut (.I0(GND_net), .I1(rand_data[27]), 
            .I2(rand_setpoint[27]), .I3(n16438), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_29 (.CI(n16438), .I0(rand_data[27]), 
            .I1(rand_setpoint[27]), .CO(n16439));
    SB_LUT4 rand_setpoint_2270_add_4_28_lut (.I0(GND_net), .I1(rand_data[26]), 
            .I2(rand_setpoint[26]), .I3(n16437), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_28 (.CI(n16437), .I0(rand_data[26]), 
            .I1(rand_setpoint[26]), .CO(n16438));
    SB_LUT4 i7576_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[1]), .I2(n320), 
            .I3(r_SM_Main_adj_2665[2]), .O(n9992));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7576_4_lut.LUT_INIT = 16'h88a0;
    SB_CARRY blink_counter_2271_add_4_4 (.CI(n16381), .I0(GND_net), .I1(n24), 
            .CO(n16382));
    SB_LUT4 i7580_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[2]), .I2(n319), 
            .I3(r_SM_Main_adj_2665[2]), .O(n9996));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7580_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 blink_counter_2271_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(n16380), .O(n134_adj_2614)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7684_3_lut (.I0(\data_in[4] [5]), .I1(\data_in[5] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10100));   // coms.v(402[9] 410[5])
    defparam i7684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10793_3_lut (.I0(\data_in[4] [0]), .I1(\data_in[5] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10101));   // coms.v(377[7:20])
    defparam i10793_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_3 (.CI(n16380), .I0(GND_net), .I1(n25), 
            .CO(n16381));
    SB_LUT4 i7686_3_lut (.I0(\data_in[3] [5]), .I1(\data_in[4] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10102));   // coms.v(402[9] 410[5])
    defparam i7686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7688_3_lut (.I0(\data_in[3] [3]), .I1(\data_in[4] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10104));   // coms.v(402[9] 410[5])
    defparam i7688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7689_3_lut (.I0(\data_in[3] [2]), .I1(\data_in[4] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10105));   // coms.v(402[9] 410[5])
    defparam i7689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7690_3_lut (.I0(\data_in[3] [1]), .I1(\data_in[4] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10106));   // coms.v(402[9] 410[5])
    defparam i7690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7692_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10108));   // coms.v(402[9] 410[5])
    defparam i7692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7693_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10109));   // coms.v(402[9] 410[5])
    defparam i7693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8087_3_lut (.I0(\data_out_frame2[6] [3]), .I1(rand_data[19]), 
            .I2(n9606), .I3(GND_net), .O(n10503));   // coms.v(428[12] 532[6])
    defparam i8087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8088_3_lut (.I0(\data_out_frame2[6] [4]), .I1(rand_data[20]), 
            .I2(n9606), .I3(GND_net), .O(n10504));   // coms.v(428[12] 532[6])
    defparam i8088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7694_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10110));   // coms.v(402[9] 410[5])
    defparam i7694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8089_3_lut (.I0(\data_out_frame2[6] [5]), .I1(rand_data[21]), 
            .I2(n9606), .I3(GND_net), .O(n10505));   // coms.v(428[12] 532[6])
    defparam i8089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8090_3_lut (.I0(\data_out_frame2[6] [6]), .I1(rand_data[22]), 
            .I2(n9606), .I3(GND_net), .O(n10506));   // coms.v(428[12] 532[6])
    defparam i8090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7583_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[3]), .I2(n318), 
            .I3(r_SM_Main_adj_2665[2]), .O(n9999));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7583_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i8091_3_lut (.I0(\data_out_frame2[6] [7]), .I1(rand_data[23]), 
            .I2(n9606), .I3(GND_net), .O(n10507));   // coms.v(428[12] 532[6])
    defparam i8091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7586_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[4]), .I2(n317), 
            .I3(r_SM_Main_adj_2665[2]), .O(n10002));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7586_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i7592_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[5]), .I2(n316), 
            .I3(r_SM_Main_adj_2665[2]), .O(n10008));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7592_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i7981_3_lut (.I0(\data_in[9] [1]), .I1(\data_in[10] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10397));   // coms.v(402[9] 410[5])
    defparam i7981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8092_3_lut (.I0(\data_out_frame2[7] [0]), .I1(rand_data[8]), 
            .I2(n9606), .I3(GND_net), .O(n10508));   // coms.v(428[12] 532[6])
    defparam i8092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut_adj_1136 (.I0(n18097), .I1(r_Clock_Count[4]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17030));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_1136.LUT_INIT = 16'hcaca;
    SB_LUT4 i7524_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4), .I3(n8567), 
            .O(n9940));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7696_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10112));   // coms.v(402[9] 410[5])
    defparam i7696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7525_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4), .I3(n8562), 
            .O(n9941));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7525_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7982_3_lut (.I0(\data_in[9] [2]), .I1(\data_in[10] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10398));   // coms.v(402[9] 410[5])
    defparam i7982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7526_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_2649), 
            .I3(n8567), .O(n9942));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7526_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8093_3_lut (.I0(\data_out_frame2[7] [1]), .I1(rand_data[9]), 
            .I2(n9606), .I3(GND_net), .O(n10509));   // coms.v(428[12] 532[6])
    defparam i8093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_27_lut (.I0(GND_net), .I1(rand_data[25]), 
            .I2(rand_setpoint[25]), .I3(n16436), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8275_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10691));   // coms.v(402[9] 410[5])
    defparam i8275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7531_2_lut (.I0(n1396), .I1(n2560), .I2(GND_net), .I3(GND_net), 
            .O(n9947));   // coms.v(428[12] 532[6])
    defparam i7531_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8094_3_lut (.I0(\data_out_frame2[7] [2]), .I1(rand_data[10]), 
            .I2(n9606), .I3(GND_net), .O(n10510));   // coms.v(428[12] 532[6])
    defparam i8094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7560_2_lut (.I0(n1396), .I1(n2561), .I2(GND_net), .I3(GND_net), 
            .O(n9976));   // coms.v(428[12] 532[6])
    defparam i7560_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8095_3_lut (.I0(\data_out_frame2[7] [3]), .I1(rand_data[11]), 
            .I2(n9606), .I3(GND_net), .O(n10511));   // coms.v(428[12] 532[6])
    defparam i8095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7698_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10114));   // coms.v(402[9] 410[5])
    defparam i7698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7522_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9938));   // coms.v(402[9] 410[5])
    defparam i7522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7561_2_lut (.I0(n1396), .I1(n2562), .I2(GND_net), .I3(GND_net), 
            .O(n9977));   // coms.v(428[12] 532[6])
    defparam i7561_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7562_2_lut (.I0(n1396), .I1(n2563), .I2(GND_net), .I3(GND_net), 
            .O(n9978));   // coms.v(428[12] 532[6])
    defparam i7562_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7983_3_lut (.I0(\data_in[9] [3]), .I1(\data_in[10] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10399));   // coms.v(402[9] 410[5])
    defparam i7983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8096_3_lut (.I0(\data_out_frame2[7] [4]), .I1(rand_data[12]), 
            .I2(n9606), .I3(GND_net), .O(n10512));   // coms.v(428[12] 532[6])
    defparam i8096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8267_4_lut (.I0(n1396), .I1(\data_in_frame[8] [7]), .I2(\data_in[8] [7]), 
            .I3(n9419), .O(n10683));   // coms.v(428[12] 532[6])
    defparam i8267_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i7563_2_lut (.I0(n1396), .I1(n2564), .I2(GND_net), .I3(GND_net), 
            .O(n9979));   // coms.v(428[12] 532[6])
    defparam i7563_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7984_3_lut (.I0(\data_in[9] [4]), .I1(\data_in[10] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10400));   // coms.v(402[9] 410[5])
    defparam i7984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7564_2_lut (.I0(n1396), .I1(n2565), .I2(GND_net), .I3(GND_net), 
            .O(n9980));   // coms.v(428[12] 532[6])
    defparam i7564_2_lut.LUT_INIT = 16'h4444;
    SB_DFF rand_data_2269__i31 (.Q(rand_data[31]), .C(CLK_c), .D(n134_adj_2602));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i15288_2_lut (.I0(delay_counter[13]), .I1(delay_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17737));
    defparam i15288_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8097_3_lut (.I0(\data_out_frame2[7] [5]), .I1(rand_data[13]), 
            .I2(n9606), .I3(GND_net), .O(n10513));   // coms.v(428[12] 532[6])
    defparam i8097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n8529), .I1(n4_adj_2612), .I2(\UART_TRANSMITTER.state [2]), 
            .I3(n121_adj_2606), .O(n13_adj_2652));   // coms.v(274[12] 374[6])
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1137 (.I0(delay_counter[14]), .I1(n13_adj_2652), 
            .I2(n13415), .I3(n17737), .O(n17312));   // coms.v(274[12] 374[6])
    defparam i4_4_lut_adj_1137.LUT_INIT = 16'h0004;
    SB_LUT4 i7700_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10116));   // coms.v(402[9] 410[5])
    defparam i7700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7985_3_lut (.I0(\data_in[9] [5]), .I1(\data_in[10] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10401));   // coms.v(402[9] 410[5])
    defparam i7985_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2269__i30 (.Q(rand_data[30]), .C(CLK_c), .D(n135_adj_2601));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i7565_2_lut (.I0(n1396), .I1(n2566), .I2(GND_net), .I3(GND_net), 
            .O(n9981));   // coms.v(428[12] 532[6])
    defparam i7565_2_lut.LUT_INIT = 16'h4444;
    SB_DFF rand_data_2269__i29 (.Q(rand_data[29]), .C(CLK_c), .D(n136_adj_2598));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i28 (.Q(rand_data[28]), .C(CLK_c), .D(n137_adj_2641));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i27 (.Q(rand_data[27]), .C(CLK_c), .D(n138_adj_2638));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i26 (.Q(rand_data[26]), .C(CLK_c), .D(n139_adj_2603));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i25 (.Q(rand_data[25]), .C(CLK_c), .D(n140_adj_2597));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i24 (.Q(rand_data[24]), .C(CLK_c), .D(n141_adj_2640));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i23 (.Q(rand_data[23]), .C(CLK_c), .D(n142_adj_2610));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i22 (.Q(rand_data[22]), .C(CLK_c), .D(n143_adj_2599));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i21 (.Q(rand_data[21]), .C(CLK_c), .D(n144_adj_2643));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i20 (.Q(rand_data[20]), .C(CLK_c), .D(n145_adj_2645));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i19 (.Q(rand_data[19]), .C(CLK_c), .D(n146_adj_2593));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8098_3_lut (.I0(\data_out_frame2[7] [6]), .I1(rand_data[14]), 
            .I2(n9606), .I3(GND_net), .O(n10514));   // coms.v(428[12] 532[6])
    defparam i8098_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2269__i18 (.Q(rand_data[18]), .C(CLK_c), .D(n147_adj_2646));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i17 (.Q(rand_data[17]), .C(CLK_c), .D(n148_adj_2639));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i16 (.Q(rand_data[16]), .C(CLK_c), .D(n149_adj_2594));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i15 (.Q(rand_data[15]), .C(CLK_c), .D(n150_adj_2644));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF blink_counter_2271__i0 (.Q(n26), .C(CLK_c), .D(n135_adj_2585));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF rand_data_2269__i14 (.Q(rand_data[14]), .C(CLK_c), .D(n151_adj_2609));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i13 (.Q(rand_data[13]), .C(CLK_c), .D(n152_adj_2590));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i12 (.Q(rand_data[12]), .C(CLK_c), .D(n153_adj_2595));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i11 (.Q(rand_data[11]), .C(CLK_c), .D(n154_adj_2591));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i10 (.Q(rand_data[10]), .C(CLK_c), .D(n155_adj_2586));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i9 (.Q(rand_data[9]), .C(CLK_c), .D(n156_adj_2596));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i8 (.Q(rand_data[8]), .C(CLK_c), .D(n157));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i7 (.Q(rand_data[7]), .C(CLK_c), .D(n158_adj_2608));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i6 (.Q(rand_data[6]), .C(CLK_c), .D(n159));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i5 (.Q(rand_data[5]), .C(CLK_c), .D(n160_adj_2607));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i4 (.Q(rand_data[4]), .C(CLK_c), .D(n161_adj_2592));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i3 (.Q(rand_data[3]), .C(CLK_c), .D(n162_adj_2600));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i2 (.Q(rand_data[2]), .C(CLK_c), .D(n163_adj_2589));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2269__i1 (.Q(rand_data[1]), .C(CLK_c), .D(n164_adj_2588));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_setpoint_2270__i0 (.Q(rand_setpoint[0]), .C(CLK_c), .D(n165));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i7566_2_lut (.I0(n1396), .I1(n2567), .I2(GND_net), .I3(GND_net), 
            .O(n9982));   // coms.v(428[12] 532[6])
    defparam i7566_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7567_2_lut (.I0(n1396), .I1(n2568), .I2(GND_net), .I3(GND_net), 
            .O(n9983));   // coms.v(428[12] 532[6])
    defparam i7567_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7569_2_lut (.I0(n1396), .I1(n2570), .I2(GND_net), .I3(GND_net), 
            .O(n9985));   // coms.v(428[12] 532[6])
    defparam i7569_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7570_2_lut (.I0(n1396), .I1(n2571), .I2(GND_net), .I3(GND_net), 
            .O(n9986));   // coms.v(428[12] 532[6])
    defparam i7570_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i10278_3_lut (.I0(\data_in[9] [6]), .I1(\data_in[10] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10402));   // coms.v(377[7:20])
    defparam i10278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7571_2_lut (.I0(n1396), .I1(n2572), .I2(GND_net), .I3(GND_net), 
            .O(n9987));   // coms.v(428[12] 532[6])
    defparam i7571_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(n12_adj_2618), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n22));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_4_lut_adj_1138 (.I0(n16466), .I1(n9390), .I2(n22), .I3(n8517), 
            .O(n17366));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_1138.LUT_INIT = 16'h5150;
    SB_CARRY rand_setpoint_2270_add_4_27 (.CI(n16436), .I0(rand_data[25]), 
            .I1(rand_setpoint[25]), .CO(n16437));
    SB_LUT4 i1_2_lut_adj_1139 (.I0(n2573), .I1(n1396), .I2(GND_net), .I3(GND_net), 
            .O(n9988));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h2222;
    SB_LUT4 i7702_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10118));   // coms.v(402[9] 410[5])
    defparam i7702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7573_2_lut (.I0(n1396), .I1(n2574), .I2(GND_net), .I3(GND_net), 
            .O(n9989));   // coms.v(428[12] 532[6])
    defparam i7573_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7703_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10119));   // coms.v(402[9] 410[5])
    defparam i7703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8099_3_lut (.I0(\data_out_frame2[7] [7]), .I1(rand_data[15]), 
            .I2(n9606), .I3(GND_net), .O(n10515));   // coms.v(428[12] 532[6])
    defparam i8099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_26_lut (.I0(GND_net), .I1(rand_data[24]), 
            .I2(rand_setpoint[24]), .I3(n16435), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8100_3_lut (.I0(\data_out_frame2[8] [0]), .I1(rand_data[0]), 
            .I2(n9606), .I3(GND_net), .O(n10516));   // coms.v(428[12] 532[6])
    defparam i8100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7667_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[1]), .I2(n225), 
            .I3(n3), .O(n10083));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7667_4_lut.LUT_INIT = 16'h4450;
    SB_CARRY rand_setpoint_2270_add_4_26 (.CI(n16435), .I0(rand_data[24]), 
            .I1(rand_setpoint[24]), .CO(n16436));
    SB_LUT4 i7577_2_lut (.I0(n1396), .I1(n2575), .I2(GND_net), .I3(GND_net), 
            .O(n9993));   // coms.v(428[12] 532[6])
    defparam i7577_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8101_3_lut (.I0(\data_out_frame2[8] [1]), .I1(rand_data[1]), 
            .I2(n9606), .I3(GND_net), .O(n10517));   // coms.v(428[12] 532[6])
    defparam i8101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_25_lut (.I0(GND_net), .I1(rand_data[23]), 
            .I2(rand_setpoint[23]), .I3(n16434), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_25 (.CI(n16434), .I0(rand_data[23]), 
            .I1(rand_setpoint[23]), .CO(n16435));
    SB_LUT4 i7987_3_lut (.I0(\data_in[9] [7]), .I1(\data_in[10] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10403));   // coms.v(402[9] 410[5])
    defparam i7987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_24_lut (.I0(GND_net), .I1(rand_data[22]), 
            .I2(rand_setpoint[22]), .I3(n16433), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2271_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26), .I3(VCC_net), .O(n135_adj_2585)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8102_3_lut (.I0(\data_out_frame2[8] [2]), .I1(rand_data[2]), 
            .I2(n9606), .I3(GND_net), .O(n10518));   // coms.v(428[12] 532[6])
    defparam i8102_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_24 (.CI(n16433), .I0(rand_data[22]), 
            .I1(rand_setpoint[22]), .CO(n16434));
    SB_CARRY rand_data_2269_add_4_16 (.CI(n16332), .I0(GND_net), .I1(rand_data[14]), 
            .CO(n16333));
    SB_LUT4 i7670_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[2]), .I2(n224), 
            .I3(n3), .O(n10086));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7670_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7587_2_lut (.I0(n1396), .I1(n2584), .I2(GND_net), .I3(GND_net), 
            .O(n10003));   // coms.v(428[12] 532[6])
    defparam i7587_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rand_setpoint_2270_add_4_23_lut (.I0(GND_net), .I1(rand_data[21]), 
            .I2(rand_setpoint[21]), .I3(n16432), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8103_3_lut (.I0(\data_out_frame2[8] [3]), .I1(rand_data[3]), 
            .I2(n9606), .I3(GND_net), .O(n10519));   // coms.v(428[12] 532[6])
    defparam i8103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7588_2_lut (.I0(n1396), .I1(n2585), .I2(GND_net), .I3(GND_net), 
            .O(n10004));   // coms.v(428[12] 532[6])
    defparam i7588_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8255_4_lut (.I0(n1396), .I1(\data_in_frame[8] [6]), .I2(\data_in[8] [6]), 
            .I3(n9419), .O(n10671));   // coms.v(428[12] 532[6])
    defparam i8255_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i7988_3_lut (.I0(\data_in[10] [0]), .I1(\data_in[11] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10404));   // coms.v(402[9] 410[5])
    defparam i7988_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_23 (.CI(n16432), .I0(rand_data[21]), 
            .I1(rand_setpoint[21]), .CO(n16433));
    SB_LUT4 rand_setpoint_2270_add_4_22_lut (.I0(GND_net), .I1(rand_data[20]), 
            .I2(rand_setpoint[20]), .I3(n16431), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33_3_lut_adj_1140 (.I0(n18054), .I1(r_Clock_Count[5]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16998));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_1140.LUT_INIT = 16'hcaca;
    SB_LUT4 i7589_2_lut (.I0(n1396), .I1(n2586), .I2(GND_net), .I3(GND_net), 
            .O(n10005));   // coms.v(428[12] 532[6])
    defparam i7589_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8104_3_lut (.I0(\data_out_frame2[8] [4]), .I1(rand_data[4]), 
            .I2(n9606), .I3(GND_net), .O(n10520));   // coms.v(428[12] 532[6])
    defparam i8104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8105_3_lut (.I0(\data_out_frame2[8] [5]), .I1(rand_data[5]), 
            .I2(n9606), .I3(GND_net), .O(n10521));   // coms.v(428[12] 532[6])
    defparam i8105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8106_3_lut (.I0(\data_out_frame2[8] [6]), .I1(rand_data[6]), 
            .I2(n9606), .I3(GND_net), .O(n10522));   // coms.v(428[12] 532[6])
    defparam i8106_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n26), 
            .CO(n16380));
    SB_LUT4 i7705_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10121));   // coms.v(402[9] 410[5])
    defparam i7705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7593_2_lut (.I0(n1396), .I1(n2587), .I2(GND_net), .I3(GND_net), 
            .O(n10009));   // coms.v(428[12] 532[6])
    defparam i7593_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7673_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[3]), .I2(n223), 
            .I3(n3), .O(n10089));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7673_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7600_2_lut (.I0(n1396), .I1(n2588), .I2(GND_net), .I3(GND_net), 
            .O(n10016));   // coms.v(428[12] 532[6])
    defparam i7600_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8107_3_lut (.I0(\data_out_frame2[8] [7]), .I1(rand_data[7]), 
            .I2(n9606), .I3(GND_net), .O(n10523));   // coms.v(428[12] 532[6])
    defparam i8107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8108_3_lut (.I0(\data_out_frame2[9] [0]), .I1(rand_data[24]), 
            .I2(n9606), .I3(GND_net), .O(n10524));   // coms.v(428[12] 532[6])
    defparam i8108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7601_2_lut (.I0(n1396), .I1(n2589), .I2(GND_net), .I3(GND_net), 
            .O(n10017));   // coms.v(428[12] 532[6])
    defparam i7601_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY rand_setpoint_2270_add_4_22 (.CI(n16431), .I0(rand_data[20]), 
            .I1(rand_setpoint[20]), .CO(n16432));
    SB_LUT4 i7676_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[4]), .I2(n222), 
            .I3(n3), .O(n10092));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7676_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7602_2_lut (.I0(n1396), .I1(n2590), .I2(GND_net), .I3(GND_net), 
            .O(n10018));   // coms.v(428[12] 532[6])
    defparam i7602_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rand_setpoint_2270_add_4_21_lut (.I0(GND_net), .I1(rand_data[19]), 
            .I2(rand_setpoint[19]), .I3(n16430), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2269_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[31]), 
            .I3(n16349), .O(n134_adj_2602)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_21 (.CI(n16430), .I0(rand_data[19]), 
            .I1(rand_setpoint[19]), .CO(n16431));
    SB_LUT4 rand_data_2269_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[13]), 
            .I3(n16331), .O(n152_adj_2590)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_15 (.CI(n16331), .I0(GND_net), .I1(rand_data[13]), 
            .CO(n16332));
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n2591), .I1(n1396), .I2(GND_net), .I3(GND_net), 
            .O(n10019));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h2222;
    SB_LUT4 i7679_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[5]), .I2(n221), 
            .I3(n3), .O(n10095));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7679_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 rand_data_2269_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[12]), 
            .I3(n16330), .O(n153_adj_2595)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2269_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[30]), 
            .I3(n16348), .O(n135_adj_2601)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2270_add_4_20_lut (.I0(GND_net), .I1(rand_data[18]), 
            .I2(rand_setpoint[18]), .I3(n16429), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_20 (.CI(n16429), .I0(rand_data[18]), 
            .I1(rand_setpoint[18]), .CO(n16430));
    SB_LUT4 rand_setpoint_2270_add_4_19_lut (.I0(GND_net), .I1(rand_data[17]), 
            .I2(rand_setpoint[17]), .I3(n16428), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_19 (.CI(n16428), .I0(rand_data[17]), 
            .I1(rand_setpoint[17]), .CO(n16429));
    SB_LUT4 i7605_2_lut (.I0(n1396), .I1(n2593), .I2(GND_net), .I3(GND_net), 
            .O(n10021));   // coms.v(428[12] 532[6])
    defparam i7605_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rand_setpoint_2270_add_4_18_lut (.I0(GND_net), .I1(rand_data[16]), 
            .I2(rand_setpoint[16]), .I3(n16427), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8109_3_lut (.I0(\data_out_frame2[9] [1]), .I1(rand_data[25]), 
            .I2(n9606), .I3(GND_net), .O(n10525));   // coms.v(428[12] 532[6])
    defparam i8109_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_32 (.CI(n16348), .I0(GND_net), .I1(rand_data[30]), 
            .CO(n16349));
    SB_CARRY rand_setpoint_2270_add_4_18 (.CI(n16427), .I0(rand_data[16]), 
            .I1(rand_setpoint[16]), .CO(n16428));
    SB_LUT4 rand_setpoint_2270_add_4_17_lut (.I0(GND_net), .I1(rand_data[15]), 
            .I2(rand_setpoint[15]), .I3(n16426), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8110_3_lut (.I0(\data_out_frame2[9] [2]), .I1(rand_data[26]), 
            .I2(n9606), .I3(GND_net), .O(n10526));   // coms.v(428[12] 532[6])
    defparam i8110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7829_4_lut (.I0(n10244), .I1(r_Clock_Count_adj_2666[0]), .I2(n321), 
            .I3(r_SM_Main_adj_2665[2]), .O(n10245));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7829_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i8111_3_lut (.I0(\data_out_frame2[9] [3]), .I1(rand_data[27]), 
            .I2(n9606), .I3(GND_net), .O(n10527));   // coms.v(428[12] 532[6])
    defparam i8111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8246_4_lut (.I0(n1396), .I1(\data_in_frame[8] [5]), .I2(\data_in[8] [5]), 
            .I3(n9419), .O(n10662));   // coms.v(428[12] 532[6])
    defparam i8246_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY rand_setpoint_2270_add_4_17 (.CI(n16426), .I0(rand_data[15]), 
            .I1(rand_setpoint[15]), .CO(n16427));
    SB_LUT4 i8112_3_lut (.I0(\data_out_frame2[9] [4]), .I1(rand_data[28]), 
            .I2(n9606), .I3(GND_net), .O(n10528));   // coms.v(428[12] 532[6])
    defparam i8112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8243_4_lut (.I0(n1396), .I1(\data_in_frame[8] [4]), .I2(\data_in[8] [4]), 
            .I3(n9419), .O(n10659));   // coms.v(428[12] 532[6])
    defparam i8243_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 rand_setpoint_2270_add_4_16_lut (.I0(GND_net), .I1(rand_data[14]), 
            .I2(rand_setpoint[14]), .I3(n16425), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_16 (.CI(n16425), .I0(rand_data[14]), 
            .I1(rand_setpoint[14]), .CO(n16426));
    SB_LUT4 rand_data_2269_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[29]), 
            .I3(n16347), .O(n136_adj_2598)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1142 (.I0(n1396), .I1(\data_in_frame[8] [3]), .I2(\data_in[8] [3]), 
            .I3(n9419), .O(n10655));
    defparam i1_4_lut_adj_1142.LUT_INIT = 16'h5044;
    SB_LUT4 i8113_3_lut (.I0(\data_out_frame2[9] [5]), .I1(rand_data[29]), 
            .I2(n9606), .I3(GND_net), .O(n10529));   // coms.v(428[12] 532[6])
    defparam i8113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7989_3_lut (.I0(\data_in[10] [1]), .I1(\data_in[11] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10405));   // coms.v(402[9] 410[5])
    defparam i7989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7606_2_lut (.I0(n1396), .I1(n2594), .I2(GND_net), .I3(GND_net), 
            .O(n10022));   // coms.v(428[12] 532[6])
    defparam i7606_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8114_3_lut (.I0(\data_out_frame2[9] [6]), .I1(rand_data[30]), 
            .I2(n9606), .I3(GND_net), .O(n10530));   // coms.v(428[12] 532[6])
    defparam i8114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8236_4_lut (.I0(n1396), .I1(\data_in_frame[8] [2]), .I2(\data_in[8] [2]), 
            .I3(n9419), .O(n10652));   // coms.v(428[12] 532[6])
    defparam i8236_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i7607_2_lut (.I0(n1396), .I1(n2595), .I2(GND_net), .I3(GND_net), 
            .O(n10023));   // coms.v(428[12] 532[6])
    defparam i7607_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8115_3_lut (.I0(\data_out_frame2[9] [7]), .I1(rand_data[31]), 
            .I2(n9606), .I3(GND_net), .O(n10531));   // coms.v(428[12] 532[6])
    defparam i8115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7990_3_lut (.I0(\data_in[10] [2]), .I1(\data_in[11] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10406));   // coms.v(402[9] 410[5])
    defparam i7990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8116_3_lut (.I0(\data_out_frame2[10] [0]), .I1(rand_data[16]), 
            .I2(n9606), .I3(GND_net), .O(n10532));   // coms.v(428[12] 532[6])
    defparam i8116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7608_2_lut (.I0(n1396), .I1(n2596), .I2(GND_net), .I3(GND_net), 
            .O(n10024));   // coms.v(428[12] 532[6])
    defparam i7608_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rand_setpoint_2270_add_4_15_lut (.I0(GND_net), .I1(rand_data[13]), 
            .I2(rand_setpoint[13]), .I3(n16424), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8233_4_lut (.I0(n1396), .I1(\data_in_frame[8] [1]), .I2(\data_in[8] [1]), 
            .I3(n9419), .O(n10649));   // coms.v(428[12] 532[6])
    defparam i8233_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i7609_2_lut (.I0(n1396), .I1(n2597), .I2(GND_net), .I3(GND_net), 
            .O(n10025));   // coms.v(428[12] 532[6])
    defparam i7609_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7991_3_lut (.I0(\data_in[10] [3]), .I1(\data_in[11] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10407));   // coms.v(402[9] 410[5])
    defparam i7991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8117_3_lut (.I0(\data_out_frame2[10] [1]), .I1(rand_data[17]), 
            .I2(n9606), .I3(GND_net), .O(n10533));   // coms.v(428[12] 532[6])
    defparam i8117_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_14 (.CI(n16330), .I0(GND_net), .I1(rand_data[12]), 
            .CO(n16331));
    SB_LUT4 i7610_2_lut (.I0(n1396), .I1(n2598), .I2(GND_net), .I3(GND_net), 
            .O(n10026));   // coms.v(428[12] 532[6])
    defparam i7610_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8181_3_lut (.I0(\data_out_frame2[18] [1]), .I1(rand_data[1]), 
            .I2(n9606), .I3(GND_net), .O(n10597));   // coms.v(428[12] 532[6])
    defparam i8181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7611_2_lut (.I0(n1396), .I1(n2599), .I2(GND_net), .I3(GND_net), 
            .O(n10027));   // coms.v(428[12] 532[6])
    defparam i7611_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25_4_lut_adj_1143 (.I0(byte_transmit_counter[7]), .I1(tx_transmit_N_2239[7]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8));   // coms.v(274[12] 374[6])
    defparam i25_4_lut_adj_1143.LUT_INIT = 16'h0aca;
    SB_CARRY rand_setpoint_2270_add_4_15 (.CI(n16424), .I0(rand_data[13]), 
            .I1(rand_setpoint[13]), .CO(n16425));
    SB_LUT4 i1_2_lut_adj_1144 (.I0(n17306), .I1(n17312), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_2615));   // coms.v(274[12] 374[6])
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h4444;
    SB_LUT4 i8118_3_lut (.I0(\data_out_frame2[10] [2]), .I1(rand_data[18]), 
            .I2(n9606), .I3(GND_net), .O(n10534));   // coms.v(428[12] 532[6])
    defparam i8118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_4_lut_adj_1145 (.I0(byte_transmit_counter[6]), .I1(tx_transmit_N_2239[6]), 
            .I2(n9631), .I3(n14_adj_2615), .O(n8_adj_2613));   // coms.v(274[12] 374[6])
    defparam i25_4_lut_adj_1145.LUT_INIT = 16'h0aca;
    SB_LUT4 i7744_3_lut (.I0(n9922), .I1(r_Bit_Index_adj_2667[0]), .I2(n9652), 
            .I3(GND_net), .O(n10160));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7744_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i7961_3_lut (.I0(\data_in[6] [5]), .I1(\data_in[7] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10377));   // coms.v(402[9] 410[5])
    defparam i7961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8182_3_lut (.I0(\data_out_frame2[18] [2]), .I1(rand_data[2]), 
            .I2(n9606), .I3(GND_net), .O(n10598));   // coms.v(428[12] 532[6])
    defparam i8182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8183_3_lut (.I0(\data_out_frame2[18] [3]), .I1(rand_data[3]), 
            .I2(n9606), .I3(GND_net), .O(n10599));   // coms.v(428[12] 532[6])
    defparam i8183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8184_3_lut (.I0(\data_out_frame2[18] [4]), .I1(rand_data[4]), 
            .I2(n9606), .I3(GND_net), .O(n10600));   // coms.v(428[12] 532[6])
    defparam i8184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[11]), 
            .I3(n16329), .O(n154_adj_2591)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_31 (.CI(n16347), .I0(GND_net), .I1(rand_data[29]), 
            .CO(n16348));
    SB_CARRY rand_data_2269_add_4_13 (.CI(n16329), .I0(GND_net), .I1(rand_data[11]), 
            .CO(n16330));
    SB_LUT4 i7992_3_lut (.I0(\data_in[10] [4]), .I1(\data_in[11] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10408));   // coms.v(402[9] 410[5])
    defparam i7992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8185_3_lut (.I0(\data_out_frame2[18] [5]), .I1(rand_data[5]), 
            .I2(n9606), .I3(GND_net), .O(n10601));   // coms.v(428[12] 532[6])
    defparam i8185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[0]), 
            .I3(VCC_net), .O(n165_adj_2587)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2270_add_4_14_lut (.I0(GND_net), .I1(rand_data[12]), 
            .I2(rand_setpoint[12]), .I3(n16423), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_14 (.CI(n16423), .I0(rand_data[12]), 
            .I1(rand_setpoint[12]), .CO(n16424));
    SB_LUT4 rand_setpoint_2270_add_4_13_lut (.I0(GND_net), .I1(rand_data[11]), 
            .I2(rand_setpoint[11]), .I3(n16422), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2269_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[28]), 
            .I3(n16346), .O(n137_adj_2641)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_13 (.CI(n16422), .I0(rand_data[11]), 
            .I1(rand_setpoint[11]), .CO(n16423));
    SB_LUT4 i8186_3_lut (.I0(\data_out_frame2[18] [6]), .I1(rand_data[6]), 
            .I2(n9606), .I3(GND_net), .O(n10602));   // coms.v(428[12] 532[6])
    defparam i8186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8119_3_lut (.I0(\data_out_frame2[10] [3]), .I1(rand_data[19]), 
            .I2(n9606), .I3(GND_net), .O(n10535));   // coms.v(428[12] 532[6])
    defparam i8119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_12_lut (.I0(GND_net), .I1(rand_data[10]), 
            .I2(rand_setpoint[10]), .I3(n16421), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8187_3_lut (.I0(\data_out_frame2[18] [7]), .I1(rand_data[7]), 
            .I2(n9606), .I3(GND_net), .O(n10603));   // coms.v(428[12] 532[6])
    defparam i8187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15277_4_lut (.I0(n16466), .I1(n13601), .I2(n17681), .I3(n12_adj_2618), 
            .O(n17356));
    defparam i15277_4_lut.LUT_INIT = 16'h1505;
    SB_LUT4 i7993_3_lut (.I0(\data_in[10] [5]), .I1(\data_in[11] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10409));   // coms.v(402[9] 410[5])
    defparam i7993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8120_3_lut (.I0(\data_out_frame2[10] [4]), .I1(rand_data[20]), 
            .I2(n9606), .I3(GND_net), .O(n10536));   // coms.v(428[12] 532[6])
    defparam i8120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7994_3_lut (.I0(\data_in[10] [6]), .I1(\data_in[11] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10410));   // coms.v(402[9] 410[5])
    defparam i7994_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_30 (.CI(n16346), .I0(GND_net), .I1(rand_data[28]), 
            .CO(n16347));
    SB_LUT4 i8121_3_lut (.I0(\data_out_frame2[10] [5]), .I1(rand_data[21]), 
            .I2(n9606), .I3(GND_net), .O(n10537));   // coms.v(428[12] 532[6])
    defparam i8121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8122_3_lut (.I0(\data_out_frame2[10] [6]), .I1(rand_data[22]), 
            .I2(n9606), .I3(GND_net), .O(n10538));   // coms.v(428[12] 532[6])
    defparam i8122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8188_3_lut (.I0(\data_out_frame2[19] [0]), .I1(n9135), .I2(n9606), 
            .I3(GND_net), .O(n10604));   // coms.v(428[12] 532[6])
    defparam i8188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8023_3_lut (.I0(\data_in[14] [3]), .I1(\data_in[15] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10439));   // coms.v(402[9] 410[5])
    defparam i8023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8024_3_lut (.I0(\data_in[14] [4]), .I1(\data_in[15] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10440));   // coms.v(402[9] 410[5])
    defparam i8024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8025_3_lut (.I0(\data_in[14] [5]), .I1(\data_in[15] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10441));   // coms.v(402[9] 410[5])
    defparam i8025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8026_3_lut (.I0(\data_in[14] [6]), .I1(\data_in[15] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10442));   // coms.v(402[9] 410[5])
    defparam i8026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8027_3_lut (.I0(\data_in[14] [7]), .I1(\data_in[15] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10443));   // coms.v(402[9] 410[5])
    defparam i8027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7995_3_lut (.I0(\data_in[10] [7]), .I1(\data_in[11] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10411));   // coms.v(402[9] 410[5])
    defparam i7995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8123_3_lut (.I0(\data_out_frame2[10] [7]), .I1(rand_data[23]), 
            .I2(n9606), .I3(GND_net), .O(n10539));   // coms.v(428[12] 532[6])
    defparam i8123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7996_3_lut (.I0(\data_in[11] [0]), .I1(\data_in[12] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10412));   // coms.v(402[9] 410[5])
    defparam i7996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8028_3_lut (.I0(\data_in[15] [0]), .I1(\data_in[16] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10444));   // coms.v(402[9] 410[5])
    defparam i8028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8029_3_lut (.I0(\data_in[15] [1]), .I1(\data_in[16] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10445));   // coms.v(402[9] 410[5])
    defparam i8029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8124_3_lut (.I0(\data_out_frame2[11] [0]), .I1(rand_data[8]), 
            .I2(n9606), .I3(GND_net), .O(n10540));   // coms.v(428[12] 532[6])
    defparam i8124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7997_3_lut (.I0(\data_in[11] [1]), .I1(\data_in[12] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10413));   // coms.v(402[9] 410[5])
    defparam i7997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8125_3_lut (.I0(\data_out_frame2[11] [1]), .I1(rand_data[9]), 
            .I2(n9606), .I3(GND_net), .O(n10541));   // coms.v(428[12] 532[6])
    defparam i8125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[27]), 
            .I3(n16345), .O(n138_adj_2638)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_29 (.CI(n16345), .I0(GND_net), .I1(rand_data[27]), 
            .CO(n16346));
    SB_LUT4 i8030_3_lut (.I0(\data_in[15] [2]), .I1(\data_in[16] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10446));   // coms.v(402[9] 410[5])
    defparam i8030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8031_3_lut (.I0(\data_in[15] [3]), .I1(\data_in[16] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10447));   // coms.v(402[9] 410[5])
    defparam i8031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7998_3_lut (.I0(\data_in[11] [2]), .I1(\data_in[12] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10414));   // coms.v(402[9] 410[5])
    defparam i7998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7930_4_lut (.I0(n9922), .I1(r_Bit_Index_adj_2667[2]), .I2(n4980), 
            .I3(n9652), .O(n10346));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7930_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i8126_3_lut (.I0(\data_out_frame2[11] [2]), .I1(rand_data[10]), 
            .I2(n9606), .I3(GND_net), .O(n10542));   // coms.v(428[12] 532[6])
    defparam i8126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut_adj_1146 (.I0(n18103), .I1(r_Clock_Count[3]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17080));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_1146.LUT_INIT = 16'hcaca;
    SB_DFF blink_counter_2271__i1 (.Q(n25), .C(CLK_c), .D(n134_adj_2614));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i7750_3_lut (.I0(n9920), .I1(r_Bit_Index_adj_2661[0]), .I2(n9646), 
            .I3(GND_net), .O(n10166));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7750_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i7999_3_lut (.I0(\data_in[11] [3]), .I1(\data_in[12] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10415));   // coms.v(402[9] 410[5])
    defparam i7999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8127_3_lut (.I0(\data_out_frame2[11] [3]), .I1(rand_data[11]), 
            .I2(n9606), .I3(GND_net), .O(n10543));   // coms.v(428[12] 532[6])
    defparam i8127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15704_4_lut (.I0(n119), .I1(\UART_TRANSMITTER.state [0]), .I2(n29), 
            .I3(n13415), .O(n17958));   // coms.v(274[12] 374[6])
    defparam i15704_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i1_3_lut_adj_1147 (.I0(\UART_TRANSMITTER.state [1]), .I1(n17364), 
            .I2(n17709), .I3(GND_net), .O(n47));   // coms.v(274[12] 374[6])
    defparam i1_3_lut_adj_1147.LUT_INIT = 16'h8a8a;
    SB_LUT4 i8000_3_lut (.I0(\data_in[11] [4]), .I1(\data_in[12] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10416));   // coms.v(402[9] 410[5])
    defparam i8000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8128_3_lut (.I0(\data_out_frame2[11] [4]), .I1(rand_data[12]), 
            .I2(n9606), .I3(GND_net), .O(n10544));   // coms.v(428[12] 532[6])
    defparam i8128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8001_3_lut (.I0(\data_in[11] [5]), .I1(\data_in[12] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10417));   // coms.v(402[9] 410[5])
    defparam i8001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8129_3_lut (.I0(\data_out_frame2[11] [5]), .I1(rand_data[13]), 
            .I2(n9606), .I3(GND_net), .O(n10545));   // coms.v(428[12] 532[6])
    defparam i8129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8002_3_lut (.I0(\data_in[11] [6]), .I1(\data_in[12] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10418));   // coms.v(402[9] 410[5])
    defparam i8002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8130_3_lut (.I0(\data_out_frame2[11] [6]), .I1(rand_data[14]), 
            .I2(n9606), .I3(GND_net), .O(n10546));   // coms.v(428[12] 532[6])
    defparam i8130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8003_3_lut (.I0(\data_in[11] [7]), .I1(\data_in[12] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10419));   // coms.v(402[9] 410[5])
    defparam i8003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8032_3_lut (.I0(\data_in[15] [4]), .I1(\data_in[16] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10448));   // coms.v(402[9] 410[5])
    defparam i8032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7979_3_lut (.I0(\data_in[8] [7]), .I1(\data_in[9] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10395));   // coms.v(402[9] 410[5])
    defparam i7979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8131_3_lut (.I0(\data_out_frame2[11] [7]), .I1(rand_data[15]), 
            .I2(n9606), .I3(GND_net), .O(n10547));   // coms.v(428[12] 532[6])
    defparam i8131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i64_4_lut (.I0(n17958), .I1(n17709), .I2(\UART_TRANSMITTER.state [1]), 
            .I3(n6878), .O(n43));   // coms.v(274[12] 374[6])
    defparam i64_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1148 (.I0(\UART_TRANSMITTER.state [2]), .I1(n47), 
            .I2(n2615), .I3(n8488), .O(n41));   // coms.v(274[12] 374[6])
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h5545;
    SB_LUT4 i8033_3_lut (.I0(\data_in[15] [5]), .I1(\data_in[16] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10449));   // coms.v(402[9] 410[5])
    defparam i8033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15884_4_lut (.I0(n41), .I1(n2615), .I2(n8488), .I3(n43), 
            .O(n38));   // coms.v(274[12] 374[6])
    defparam i15884_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i8034_3_lut (.I0(\data_in[15] [6]), .I1(\data_in[16] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10450));   // coms.v(402[9] 410[5])
    defparam i8034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15893_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026 [1]), 
            .I2(\FRAME_MATCHER.next_state [1]), .I3(n63_adj_2642), .O(n6_adj_2616));   // coms.v(428[12] 532[6])
    defparam i15893_4_lut.LUT_INIT = 16'hc4cc;
    SB_LUT4 rand_data_2269_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[10]), 
            .I3(n16328), .O(n155_adj_2586)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(rand_data[0]), 
            .CO(n16319));
    SB_LUT4 i7516_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9932));   // coms.v(402[9] 410[5])
    defparam i7516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7517_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_2582), 
            .I3(n8562), .O(n9933));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7517_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7518_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9934));   // coms.v(402[9] 410[5])
    defparam i7518_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_12 (.CI(n16421), .I0(rand_data[10]), 
            .I1(rand_setpoint[10]), .CO(n16422));
    SB_LUT4 i7519_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9935));   // coms.v(402[9] 410[5])
    defparam i7519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_11_lut (.I0(GND_net), .I1(rand_data[9]), 
            .I2(rand_setpoint[9]), .I3(n16420), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_11 (.CI(n16420), .I0(rand_data[9]), 
            .I1(rand_setpoint[9]), .CO(n16421));
    SB_LUT4 i8209_4_lut (.I0(n9922), .I1(r_Bit_Index_adj_2667[1]), .I2(r_Bit_Index_adj_2667[0]), 
            .I3(n9652), .O(n10625));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8209_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 rand_setpoint_2270_add_4_10_lut (.I0(GND_net), .I1(rand_data[8]), 
            .I2(rand_setpoint[8]), .I3(n16419), .O(n157_adj_2581)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_10 (.CI(n16419), .I0(rand_data[8]), 
            .I1(rand_setpoint[8]), .CO(n16420));
    SB_LUT4 i7969_3_lut (.I0(\data_in[7] [5]), .I1(\data_in[8] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10385));   // coms.v(402[9] 410[5])
    defparam i7969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7521_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9937));   // coms.v(402[9] 410[5])
    defparam i7521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7980_3_lut (.I0(\data_in[9] [0]), .I1(\data_in[10] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10396));   // coms.v(402[9] 410[5])
    defparam i7980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8212_4_lut (.I0(n9920), .I1(r_Bit_Index_adj_2661[2]), .I2(n4958), 
            .I3(n9646), .O(n10628));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8212_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i8035_3_lut (.I0(\data_in[15] [7]), .I1(\data_in[16] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10451));   // coms.v(402[9] 410[5])
    defparam i8035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7947_3_lut (.I0(\data_in[4] [7]), .I1(\data_in[5] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10363));   // coms.v(402[9] 410[5])
    defparam i7947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7728_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10144));   // coms.v(402[9] 410[5])
    defparam i7728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8036_3_lut (.I0(\data_in[16] [0]), .I1(\data_in[17] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10452));   // coms.v(402[9] 410[5])
    defparam i8036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2270_add_4_9_lut (.I0(GND_net), .I1(rand_data[7]), 
            .I2(rand_setpoint[7]), .I3(n16418), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8037_3_lut (.I0(\data_in[16] [1]), .I1(\data_in[17] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10453));   // coms.v(402[9] 410[5])
    defparam i8037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7977_3_lut (.I0(\data_in[8] [5]), .I1(\data_in[9] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10393));   // coms.v(402[9] 410[5])
    defparam i7977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7978_3_lut (.I0(\data_in[8] [6]), .I1(\data_in[9] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10394));   // coms.v(402[9] 410[5])
    defparam i7978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7950_3_lut (.I0(\data_in[5] [2]), .I1(\data_in[6] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10366));   // coms.v(402[9] 410[5])
    defparam i7950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8038_3_lut (.I0(\data_in[16] [2]), .I1(\data_in[17] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10454));   // coms.v(402[9] 410[5])
    defparam i8038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7754_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_2649), 
            .I3(n8562), .O(n10170));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7754_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY rand_setpoint_2270_add_4_9 (.CI(n16418), .I0(rand_data[7]), 
            .I1(rand_setpoint[7]), .CO(n16419));
    SB_DFF blink_counter_2271__i2 (.Q(n24), .C(CLK_c), .D(n133));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i3 (.Q(n23), .C(CLK_c), .D(n132));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i4 (.Q(n22_adj_2655), .C(CLK_c), .D(n131));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i5 (.Q(n21), .C(CLK_c), .D(n130));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i6 (.Q(n20), .C(CLK_c), .D(n129));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i7 (.Q(n19), .C(CLK_c), .D(n128));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i8 (.Q(n18), .C(CLK_c), .D(n127));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i9 (.Q(n17), .C(CLK_c), .D(n126));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i10 (.Q(n16), .C(CLK_c), .D(n125));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i11 (.Q(n15), .C(CLK_c), .D(n124));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i12 (.Q(n14), .C(CLK_c), .D(n123));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i13 (.Q(n13), .C(CLK_c), .D(n122));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i14 (.Q(n12), .C(CLK_c), .D(n121));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i15 (.Q(n11), .C(CLK_c), .D(n120));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i16 (.Q(n10), .C(CLK_c), .D(n119_adj_2648));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i17 (.Q(n9), .C(CLK_c), .D(n118));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i18 (.Q(n8_adj_2617), .C(CLK_c), .D(n117));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i19 (.Q(n7), .C(CLK_c), .D(n116));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i20 (.Q(n6), .C(CLK_c), .D(n115));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i21 (.Q(blink_counter[21]), .C(CLK_c), .D(n114));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i22 (.Q(blink_counter[22]), .C(CLK_c), .D(n113));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i23 (.Q(blink_counter[23]), .C(CLK_c), .D(n112));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i24 (.Q(blink_counter[24]), .C(CLK_c), .D(n111));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2271__i25 (.Q(blink_counter[25]), .C(CLK_c), .D(n110));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF rand_setpoint_2270__i1 (.Q(rand_setpoint[1]), .C(CLK_c), .D(n164));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n7364), .I1(n18098), .I2(n7086), .I3(r_SM_Main[2]), 
            .O(n17028));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'hafec;
    SB_DFF rand_setpoint_2270__i2 (.Q(rand_setpoint[2]), .C(CLK_c), .D(n163));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i8039_3_lut (.I0(\data_in[16] [3]), .I1(\data_in[17] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10455));   // coms.v(402[9] 410[5])
    defparam i8039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8040_3_lut (.I0(\data_in[16] [4]), .I1(\data_in[17] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10456));   // coms.v(402[9] 410[5])
    defparam i8040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8041_3_lut (.I0(\data_in[16] [5]), .I1(\data_in[17] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10457));   // coms.v(402[9] 410[5])
    defparam i8041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8] [4]), 
            .I2(\data_in_frame[6] [5]), .I3(n9283), .O(n16_adj_2656));   // coms.v(383[12:25])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8042_3_lut (.I0(\data_in[16] [6]), .I1(\data_in[17] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10458));   // coms.v(402[9] 410[5])
    defparam i8042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8004_3_lut (.I0(\data_in[12] [0]), .I1(\data_in[13] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10420));   // coms.v(402[9] 410[5])
    defparam i8004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8132_3_lut (.I0(\data_out_frame2[12] [0]), .I1(rand_data[0]), 
            .I2(n9606), .I3(GND_net), .O(n10548));   // coms.v(428[12] 532[6])
    defparam i8132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8043_3_lut (.I0(\data_in[16] [7]), .I1(\data_in[17] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10459));   // coms.v(402[9] 410[5])
    defparam i8043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut_adj_1150 (.I0(n18104), .I1(r_Clock_Count[0]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17078));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_1150.LUT_INIT = 16'hcaca;
    SB_LUT4 i8044_3_lut (.I0(\data_in[17] [0]), .I1(\data_in[18] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10460));   // coms.v(402[9] 410[5])
    defparam i8044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8133_3_lut (.I0(\data_out_frame2[12] [1]), .I1(rand_data[1]), 
            .I2(n9606), .I3(GND_net), .O(n10549));   // coms.v(428[12] 532[6])
    defparam i8133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8134_3_lut (.I0(\data_out_frame2[12] [2]), .I1(rand_data[2]), 
            .I2(n9606), .I3(GND_net), .O(n10550));   // coms.v(428[12] 532[6])
    defparam i8134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8045_3_lut (.I0(\data_in[17] [1]), .I1(\data_in[18] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10461));   // coms.v(402[9] 410[5])
    defparam i8045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8046_3_lut (.I0(\data_in[17] [2]), .I1(\data_in[18] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10462));   // coms.v(402[9] 410[5])
    defparam i8046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15406_4_lut (.I0(blink_counter[22]), .I1(blink_counter[23]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17856));
    defparam i15406_4_lut.LUT_INIT = 16'hfec4;
    SB_LUT4 i15405_4_lut (.I0(blink_counter[23]), .I1(blink_counter[22]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17855));
    defparam i15405_4_lut.LUT_INIT = 16'hcf08;
    SB_LUT4 i15407_3_lut (.I0(n17855), .I1(n17856), .I2(blink_counter[25]), 
            .I3(GND_net), .O(LED_c));
    defparam i15407_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i8135_3_lut (.I0(\data_out_frame2[12] [3]), .I1(rand_data[3]), 
            .I2(n9606), .I3(GND_net), .O(n10551));   // coms.v(428[12] 532[6])
    defparam i8135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8047_3_lut (.I0(\data_in[17] [3]), .I1(\data_in[18] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10463));   // coms.v(402[9] 410[5])
    defparam i8047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8048_3_lut (.I0(\data_in[17] [4]), .I1(\data_in[18] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10464));   // coms.v(402[9] 410[5])
    defparam i8048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7721_3_lut_4_lut (.I0(\data_out[1] [2]), .I1(\UART_TRANSMITTER.state [2]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n9519), .O(n10137));   // coms.v(274[12] 374[6])
    defparam i7721_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i8136_3_lut (.I0(\data_out_frame2[12] [4]), .I1(rand_data[4]), 
            .I2(n9606), .I3(GND_net), .O(n10552));   // coms.v(428[12] 532[6])
    defparam i8136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8137_3_lut (.I0(\data_out_frame2[12] [5]), .I1(rand_data[5]), 
            .I2(n9606), .I3(GND_net), .O(n10553));   // coms.v(428[12] 532[6])
    defparam i8137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8138_3_lut (.I0(\data_out_frame2[12] [6]), .I1(rand_data[6]), 
            .I2(n9606), .I3(GND_net), .O(n10554));   // coms.v(428[12] 532[6])
    defparam i8138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7778_4_lut (.I0(n13880), .I1(r_Clock_Count_adj_2660[0]), .I2(n226), 
            .I3(n3), .O(n10194));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7778_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[8] [3]), .I1(n19_adj_2651), 
            .I2(n9100), .I3(n9148), .O(n17585));   // coms.v(383[12:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8049_3_lut (.I0(\data_in[17] [5]), .I1(\data_in[18] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10465));   // coms.v(402[9] 410[5])
    defparam i8049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1151 (.I0(\FRAME_MATCHER.next_state [0]), .I1(n63_adj_2642), 
            .I2(n63), .I3(\FRAME_MATCHER.next_state_31__N_2026 [1]), .O(n17092));   // coms.v(428[12] 532[6])
    defparam i1_4_lut_adj_1151.LUT_INIT = 16'hb3ff;
    SB_LUT4 i11594214_i1_3_lut (.I0(n18465), .I1(n18441), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n1));
    defparam i11594214_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8222_3_lut (.I0(r_Tx_Data[7]), .I1(i_Tx_Byte[7]), .I2(n7734), 
            .I3(GND_net), .O(n10638));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[26]), 
            .I3(n16344), .O(n139_adj_2603)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2270_add_4_8_lut (.I0(GND_net), .I1(rand_data[6]), 
            .I2(rand_setpoint[6]), .I3(n16417), .O(n159_adj_2580)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_28 (.CI(n16344), .I0(GND_net), .I1(rand_data[26]), 
            .CO(n16345));
    SB_LUT4 i7907_3_lut (.I0(tx_o_adj_2584), .I1(n3_adj_2650), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n10323));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7962_3_lut (.I0(\data_in[6] [6]), .I1(\data_in[7] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10378));   // coms.v(402[9] 410[5])
    defparam i7962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7963_3_lut (.I0(\data_in[6] [7]), .I1(\data_in[7] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10379));   // coms.v(402[9] 410[5])
    defparam i7963_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2270_add_4_8 (.CI(n16417), .I0(rand_data[6]), 
            .I1(rand_setpoint[6]), .CO(n16418));
    SB_LUT4 rand_setpoint_2270_add_4_7_lut (.I0(GND_net), .I1(rand_data[5]), 
            .I2(rand_setpoint[5]), .I3(n16416), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2270__i3 (.Q(rand_setpoint[3]), .C(CLK_c), .D(n162));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i4 (.Q(rand_setpoint[4]), .C(CLK_c), .D(n161));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i5 (.Q(rand_setpoint[5]), .C(CLK_c), .D(n160));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i6 (.Q(rand_setpoint[6]), .C(CLK_c), .D(n159_adj_2580));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i7 (.Q(rand_setpoint[7]), .C(CLK_c), .D(n158));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i8 (.Q(rand_setpoint[8]), .C(CLK_c), .D(n157_adj_2581));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i9 (.Q(rand_setpoint[9]), .C(CLK_c), .D(n156));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i10 (.Q(rand_setpoint[10]), .C(CLK_c), .D(n155));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i11 (.Q(rand_setpoint[11]), .C(CLK_c), .D(n154));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i12 (.Q(rand_setpoint[12]), .C(CLK_c), .D(n153));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i13 (.Q(rand_setpoint[13]), .C(CLK_c), .D(n152));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i14 (.Q(rand_setpoint[14]), .C(CLK_c), .D(n151));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i15 (.Q(rand_setpoint[15]), .C(CLK_c), .D(n150));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i16 (.Q(rand_setpoint[16]), .C(CLK_c), .D(n149));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i17 (.Q(rand_setpoint[17]), .C(CLK_c), .D(n148));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i18 (.Q(rand_setpoint[18]), .C(CLK_c), .D(n147));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i19 (.Q(rand_setpoint[19]), .C(CLK_c), .D(n146));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i20 (.Q(rand_setpoint[20]), .C(CLK_c), .D(n145));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i21 (.Q(rand_setpoint[21]), .C(CLK_c), .D(n144));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i22 (.Q(rand_setpoint[22]), .C(CLK_c), .D(n143));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i23 (.Q(rand_setpoint[23]), .C(CLK_c), .D(n142));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i24 (.Q(rand_setpoint[24]), .C(CLK_c), .D(n141));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i25 (.Q(rand_setpoint[25]), .C(CLK_c), .D(n140));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i26 (.Q(rand_setpoint[26]), .C(CLK_c), .D(n139));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i27 (.Q(rand_setpoint[27]), .C(CLK_c), .D(n138));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i28 (.Q(rand_setpoint[28]), .C(CLK_c), .D(n137));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i29 (.Q(rand_setpoint[29]), .C(CLK_c), .D(n136));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i30 (.Q(rand_setpoint[30]), .C(CLK_c), .D(n135));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2270__i31 (.Q(rand_setpoint[31]), .C(CLK_c), .D(n134));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_CARRY rand_setpoint_2270_add_4_7 (.CI(n16416), .I0(rand_data[5]), 
            .I1(rand_setpoint[5]), .CO(n16417));
    SB_LUT4 rand_setpoint_2270_add_4_6_lut (.I0(GND_net), .I1(rand_data[4]), 
            .I2(rand_setpoint[4]), .I3(n16415), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_6 (.CI(n16415), .I0(rand_data[4]), 
            .I1(rand_setpoint[4]), .CO(n16416));
    SB_LUT4 i2_3_lut_adj_1152 (.I0(\UART_TRANSMITTER.state [0]), .I1(n96), 
            .I2(n29), .I3(GND_net), .O(n17364));   // coms.v(274[12] 374[6])
    defparam i2_3_lut_adj_1152.LUT_INIT = 16'h4040;
    SB_LUT4 rand_data_2269_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[25]), 
            .I3(n16343), .O(n140_adj_2597)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15721_4_lut (.I0(\UART_TRANSMITTER.state_7__N_1749 [2]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(\UART_TRANSMITTER.state [2]), 
            .O(n18032));   // coms.v(274[12] 374[6])
    defparam i15721_4_lut.LUT_INIT = 16'h0203;
    SB_LUT4 i12_4_lut (.I0(\UART_TRANSMITTER.state [0]), .I1(n18032), .I2(n16485), 
            .I3(n17672), .O(n16864));   // coms.v(274[12] 374[6])
    defparam i12_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 rand_setpoint_2270_add_4_5_lut (.I0(GND_net), .I1(rand_data[3]), 
            .I2(rand_setpoint[3]), .I3(n16414), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_27 (.CI(n16343), .I0(GND_net), .I1(rand_data[25]), 
            .CO(n16344));
    SB_CARRY rand_setpoint_2270_add_4_5 (.CI(n16414), .I0(rand_data[3]), 
            .I1(rand_setpoint[3]), .CO(n16415));
    SB_LUT4 i25_3_lut (.I0(r_Clock_Count[6]), .I1(n18010), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16968));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rand_setpoint_2270_add_4_4_lut (.I0(GND_net), .I1(rand_data[2]), 
            .I2(rand_setpoint[2]), .I3(n16413), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_4 (.CI(n16413), .I0(rand_data[2]), 
            .I1(rand_setpoint[2]), .CO(n16414));
    SB_CARRY rand_data_2269_add_4_12 (.CI(n16328), .I0(GND_net), .I1(rand_data[10]), 
            .CO(n16329));
    SB_LUT4 rand_data_2269_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[24]), 
            .I3(n16342), .O(n141_adj_2640)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25_3_lut_adj_1153 (.I0(r_Clock_Count[7]), .I1(n17952), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16954));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_1153.LUT_INIT = 16'hacac;
    SB_LUT4 i25_3_lut_adj_1154 (.I0(r_Clock_Count[8]), .I1(n17950), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16932));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_1154.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut (.I0(n17757), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17054));   // verilog/uart_tx.v(33[16:27])
    defparam i12_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 i7711_3_lut_4_lut (.I0(data_out_5__4__N_959), .I1(n2720), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n4430), .O(n10127));   // coms.v(274[12] 374[6])
    defparam i7711_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7908_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n4_adj_2653), .O(n10324));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7908_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i7628_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [0]), .I2(\data_in[5] [0]), 
            .I3(n16468), .O(n10044));   // coms.v(428[12] 532[6])
    defparam i7628_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7970_3_lut (.I0(\data_in[7] [6]), .I1(\data_in[8] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10386));   // coms.v(402[9] 410[5])
    defparam i7970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15234_3_lut_4_lut (.I0(n12_adj_2618), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n9390), .O(n17681));
    defparam i15234_3_lut_4_lut.LUT_INIT = 16'hf7f3;
    SB_LUT4 i7627_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [1]), .I2(\data_in[5] [1]), 
            .I3(n16468), .O(n10043));   // coms.v(428[12] 532[6])
    defparam i7627_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7909_3_lut (.I0(r_Tx_Data[0]), .I1(i_Tx_Byte[0]), .I2(n7734), 
            .I3(GND_net), .O(n10325));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7971_3_lut (.I0(\data_in[7] [7]), .I1(\data_in[8] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10387));   // coms.v(402[9] 410[5])
    defparam i7971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1155 (.I0(n1396), .I1(\data_in_frame[8] [0]), .I2(\data_in[8] [0]), 
            .I3(n9419), .O(n10631));
    defparam i1_4_lut_adj_1155.LUT_INIT = 16'h5044;
    SB_LUT4 i7910_4_lut (.I0(r_SM_Main[2]), .I1(n7080), .I2(r_SM_Main_2__N_2323[1]), 
            .I3(r_SM_Main[0]), .O(n10326));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7910_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i7623_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [2]), .I2(\data_in[5] [2]), 
            .I3(n16468), .O(n10039));   // coms.v(428[12] 532[6])
    defparam i7623_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7622_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [3]), .I2(\data_in[5] [3]), 
            .I3(n16468), .O(n10038));   // coms.v(428[12] 532[6])
    defparam i7622_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7710_3_lut_4_lut (.I0(\data_out[3] [4]), .I1(n2720), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n4430), .O(n10126));   // coms.v(274[12] 374[6])
    defparam i7710_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7618_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [4]), .I2(\data_in[5] [4]), 
            .I3(n16468), .O(n10034));   // coms.v(428[12] 532[6])
    defparam i7618_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i9728_3_lut (.I0(r_Tx_Data[1]), .I1(i_Tx_Byte[1]), .I2(n7734), 
            .I3(GND_net), .O(n10632));
    defparam i9728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7617_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [5]), .I2(\data_in[5] [5]), 
            .I3(n16468), .O(n10033));   // coms.v(428[12] 532[6])
    defparam i7617_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i8050_3_lut (.I0(\data_in[17] [6]), .I1(\data_in[18] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10466));   // coms.v(402[9] 410[5])
    defparam i8050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7616_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [6]), .I2(\data_in[5] [6]), 
            .I3(n16468), .O(n10032));   // coms.v(428[12] 532[6])
    defparam i7616_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i8051_3_lut (.I0(\data_in[17] [7]), .I1(\data_in[18] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10467));   // coms.v(402[9] 410[5])
    defparam i8051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7615_2_lut_4_lut (.I0(n1396), .I1(\data_in_frame[5] [7]), .I2(\data_in[5] [7]), 
            .I3(n16468), .O(n10031));   // coms.v(428[12] 532[6])
    defparam i7615_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i7964_3_lut (.I0(\data_in[7] [0]), .I1(\data_in[8] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10380));   // coms.v(402[9] 410[5])
    defparam i7964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7966_3_lut (.I0(\data_in[7] [2]), .I1(\data_in[8] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10382));   // coms.v(402[9] 410[5])
    defparam i7966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7967_3_lut (.I0(\data_in[7] [3]), .I1(\data_in[8] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10383));   // coms.v(402[9] 410[5])
    defparam i7967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8052_3_lut (.I0(\data_in[18] [0]), .I1(\data_in[19] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10468));   // coms.v(402[9] 410[5])
    defparam i8052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7708_3_lut_4_lut (.I0(\data_out[3] [6]), .I1(\UART_TRANSMITTER.state [2]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n9519), .O(n10124));   // coms.v(274[12] 374[6])
    defparam i7708_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i8053_3_lut (.I0(\data_in[18] [1]), .I1(\data_in[19] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10469));   // coms.v(402[9] 410[5])
    defparam i8053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8054_3_lut (.I0(\data_in[18] [2]), .I1(\data_in[19] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10470));   // coms.v(402[9] 410[5])
    defparam i8054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9727_3_lut (.I0(r_Tx_Data[2]), .I1(i_Tx_Byte[2]), .I2(n7734), 
            .I3(GND_net), .O(n10633));
    defparam i9727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7724_3_lut_4_lut (.I0(\data_out[0] [3]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10140));   // coms.v(274[12] 374[6])
    defparam i7724_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 rand_setpoint_2270_add_4_3_lut (.I0(GND_net), .I1(rand_data[1]), 
            .I2(rand_setpoint[1]), .I3(n16412), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_3 (.CI(n16412), .I0(rand_data[1]), 
            .I1(rand_setpoint[1]), .CO(n16413));
    SB_LUT4 rand_setpoint_2270_add_4_2_lut (.I0(GND_net), .I1(rand_data[0]), 
            .I2(rand_setpoint[0]), .I3(GND_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2270_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2270_add_4_2 (.CI(GND_net), .I0(rand_data[0]), 
            .I1(rand_setpoint[0]), .CO(n16412));
    SB_CARRY rand_data_2269_add_4_26 (.CI(n16342), .I0(GND_net), .I1(rand_data[24]), 
            .CO(n16343));
    SB_LUT4 rand_data_2269_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[23]), 
            .I3(n16341), .O(n142_adj_2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7556_4_lut_4_lut (.I0(n17757), .I1(n9796), .I2(r_Bit_Index[1]), 
            .I3(r_Bit_Index[0]), .O(n9972));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7556_4_lut_4_lut.LUT_INIT = 16'ha4e0;
    SB_LUT4 i7726_3_lut_4_lut_4_lut (.I0(\data_out[0] [0]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10142));   // coms.v(274[12] 374[6])
    defparam i7726_3_lut_4_lut_4_lut.LUT_INIT = 16'haaca;
    SB_CARRY rand_data_2269_add_4_25 (.CI(n16341), .I0(GND_net), .I1(rand_data[23]), 
            .CO(n16342));
    SB_LUT4 rand_data_2269_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[9]), 
            .I3(n16327), .O(n156_adj_2596)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7931_3_lut (.I0(\data_in[4] [3]), .I1(\data_in[5] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10347));   // coms.v(402[9] 410[5])
    defparam i7931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2269_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[22]), 
            .I3(n16340), .O(n143_adj_2599)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7935_3_lut (.I0(\data_out[8] [7]), .I1(rand_setpoint[7]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10351));   // coms.v(274[12] 374[6])
    defparam i7935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7936_3_lut (.I0(\data_out[8] [6]), .I1(rand_setpoint[6]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10352));   // coms.v(274[12] 374[6])
    defparam i7936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7937_3_lut (.I0(\data_out[8] [5]), .I1(rand_setpoint[5]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10353));   // coms.v(274[12] 374[6])
    defparam i7937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7941_3_lut (.I0(\data_out[8] [4]), .I1(rand_setpoint[4]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10357));   // coms.v(274[12] 374[6])
    defparam i7941_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_24 (.CI(n16340), .I0(GND_net), .I1(rand_data[22]), 
            .CO(n16341));
    SB_LUT4 i7942_3_lut (.I0(\data_out[8] [3]), .I1(rand_setpoint[3]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10358));   // coms.v(274[12] 374[6])
    defparam i7942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7943_3_lut (.I0(\data_out[8] [2]), .I1(rand_setpoint[2]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10359));   // coms.v(274[12] 374[6])
    defparam i7943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2269_add_4_11 (.CI(n16327), .I0(GND_net), .I1(rand_data[9]), 
            .CO(n16328));
    SB_LUT4 i7944_3_lut (.I0(\data_out[8] [1]), .I1(rand_setpoint[1]), .I2(data_out_10__7__N_114), 
            .I3(GND_net), .O(n10360));   // coms.v(274[12] 374[6])
    defparam i7944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7723_3_lut_4_lut (.I0(\data_out[0] [5]), .I1(n2720), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n4430), .O(n10139));   // coms.v(274[12] 374[6])
    defparam i7723_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rand_data_2269_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[21]), 
            .I3(n16339), .O(n144_adj_2643)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7707_3_lut_4_lut_4_lut (.I0(data_out_5__7__N_931), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10123));   // coms.v(274[12] 374[6])
    defparam i7707_3_lut_4_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 blink_counter_2271_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[25]), .I3(n16404), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7725_3_lut_4_lut (.I0(\data_out[0] [1]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10141));   // coms.v(274[12] 374[6])
    defparam i7725_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 blink_counter_2271_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[24]), .I3(n16403), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7709_3_lut_4_lut_4_lut (.I0(\data_out[3] [5]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10125));   // coms.v(274[12] 374[6])
    defparam i7709_3_lut_4_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rand_data_2269_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[8]), 
            .I3(n16326), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_26 (.CI(n16403), .I0(GND_net), .I1(blink_counter[24]), 
            .CO(n16404));
    SB_LUT4 blink_counter_2271_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[23]), .I3(n16402), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7719_3_lut_4_lut_4_lut (.I0(\data_out[1] [6]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10135));   // coms.v(274[12] 374[6])
    defparam i7719_3_lut_4_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7718_3_lut_4_lut (.I0(\data_out[1] [7]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10134));   // coms.v(274[12] 374[6])
    defparam i7718_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 i2_3_lut_4_lut_adj_1156 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[8] [0]), 
            .I2(n6_adj_2583), .I3(n2573), .O(n17481));   // coms.v(383[12:25])
    defparam i2_3_lut_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_CARRY blink_counter_2271_add_4_25 (.CI(n16402), .I0(GND_net), .I1(blink_counter[23]), 
            .CO(n16403));
    SB_LUT4 blink_counter_2271_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[22]), .I3(n16401), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_10 (.CI(n16326), .I0(GND_net), .I1(rand_data[8]), 
            .CO(n16327));
    SB_CARRY blink_counter_2271_add_4_24 (.CI(n16401), .I0(GND_net), .I1(blink_counter[22]), 
            .CO(n16402));
    GND i1 (.Y(GND_net));
    SB_LUT4 blink_counter_2271_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[21]), .I3(n16400), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_23 (.CI(n16400), .I0(GND_net), .I1(blink_counter[21]), 
            .CO(n16401));
    SB_LUT4 blink_counter_2271_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n16399), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7717_3_lut_4_lut (.I0(\data_out[2] [0]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10133));   // coms.v(274[12] 374[6])
    defparam i7717_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_CARRY blink_counter_2271_add_4_22 (.CI(n16399), .I0(GND_net), .I1(n6), 
            .CO(n16400));
    SB_LUT4 blink_counter_2271_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n16398), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_21 (.CI(n16398), .I0(GND_net), .I1(n7), 
            .CO(n16399));
    SB_LUT4 rand_data_2269_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[7]), 
            .I3(n16325), .O(n158_adj_2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2271_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_2617), .I3(n16397), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_20 (.CI(n16397), .I0(GND_net), .I1(n8_adj_2617), 
            .CO(n16398));
    SB_LUT4 blink_counter_2271_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n16396), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_23 (.CI(n16339), .I0(GND_net), .I1(rand_data[21]), 
            .CO(n16340));
    SB_CARRY blink_counter_2271_add_4_19 (.CI(n16396), .I0(GND_net), .I1(n9), 
            .CO(n16397));
    SB_LUT4 blink_counter_2271_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10), .I3(n16395), .O(n119_adj_2648)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2269_add_4_9 (.CI(n16325), .I0(GND_net), .I1(rand_data[7]), 
            .CO(n16326));
    SB_LUT4 i7716_3_lut_4_lut (.I0(data_out_6__6__N_729), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10132));   // coms.v(274[12] 374[6])
    defparam i7716_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 i7714_3_lut_4_lut (.I0(data_out_6__7__N_678), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10130));   // coms.v(274[12] 374[6])
    defparam i7714_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 i7713_3_lut_4_lut (.I0(data_out_6__1__N_850), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(n4430), .O(n10129));   // coms.v(274[12] 374[6])
    defparam i7713_3_lut_4_lut.LUT_INIT = 16'haa3a;
    SB_LUT4 i8139_3_lut (.I0(\data_out_frame2[12] [7]), .I1(rand_data[7]), 
            .I2(n9606), .I3(GND_net), .O(n10555));   // coms.v(428[12] 532[6])
    defparam i8139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8140_3_lut (.I0(\data_out_frame2[13] [0]), .I1(rand_data[24]), 
            .I2(n9606), .I3(GND_net), .O(n10556));   // coms.v(428[12] 532[6])
    defparam i8140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8141_3_lut (.I0(\data_out_frame2[13] [1]), .I1(rand_data[25]), 
            .I2(n9606), .I3(GND_net), .O(n10557));   // coms.v(428[12] 532[6])
    defparam i8141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8142_3_lut (.I0(\data_out_frame2[13] [2]), .I1(rand_data[26]), 
            .I2(n9606), .I3(GND_net), .O(n10558));   // coms.v(428[12] 532[6])
    defparam i8142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10788_3_lut (.I0(\data_in[5] [0]), .I1(\data_in[6] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10364));   // coms.v(377[7:20])
    defparam i10788_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2271_add_4_18 (.CI(n16395), .I0(GND_net), .I1(n10), 
            .CO(n16396));
    SB_LUT4 i7712_3_lut_4_lut (.I0(data_out_6__2__N_804), .I1(n2720), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n4430), .O(n10128));   // coms.v(274[12] 374[6])
    defparam i7712_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 blink_counter_2271_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n16394), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2269_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[6]), 
            .I3(n16324), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2269_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_17 (.CI(n16394), .I0(GND_net), .I1(n11), 
            .CO(n16395));
    SB_LUT4 blink_counter_2271_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n16393), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2271_add_4_16 (.CI(n16393), .I0(GND_net), .I1(n12), 
            .CO(n16394));
    coms c0 (.n16485(n16485), .\UART_TRANSMITTER.state[1] (\UART_TRANSMITTER.state [1]), 
         .\UART_TRANSMITTER.state[0] (\UART_TRANSMITTER.state [0]), .i_Tx_Byte({i_Tx_Byte}), 
         .n10383(n10383), .\data_in[7] ({Open_0, Open_1, Open_2, Open_3, 
         \data_in[7] [3:2], Open_4, Open_5}), .CLK_c(CLK_c), .\data_out[3][6] (\data_out[3] [6]), 
         .n10382(n10382), .n10380(n10380), .\data_in[7][0] (\data_in[7] [0]), 
         .n10379(n10379), .\data_in[6] ({\data_in[6] [7:5], Open_6, Open_7, 
         Open_8, Open_9, Open_10}), .n10378(n10378), .GND_net(GND_net), 
         .VCC_net(VCC_net), .\data_in_frame[8] ({\data_in_frame[8] }), .n10377(n10377), 
         .\UART_TRANSMITTER.state[2] (\UART_TRANSMITTER.state [2]), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n9380(n9380), .n16(n16_adj_2656), .\rand_setpoint[8] (rand_setpoint[8]), 
         .n2565(n2565), .n2574(n2574), .\data_out[8] ({\data_out[8] }), 
         .\data_out_frame2[13] ({\data_out_frame2[13] }), .\data_out_frame2[12] ({\data_out_frame2[12] }), 
         .n9519(n9519), .\data_out_frame2[18] ({\data_out_frame2[18] }), 
         .\data_in_frame[1][1] (\data_in_frame[1] [1]), .data_out_6__7__N_678(data_out_6__7__N_678), 
         .data_out_6__1__N_850(data_out_6__1__N_850), .\data_out_frame2[17] ({\data_out_frame2[17] }), 
         .\data_out_frame2[16] ({\data_out_frame2[16] }), .\data_in[5] ({\data_in[5] }), 
         .rx_data_ready(rx_data_ready), .\data_in_frame[10][6] (\data_in_frame[10] [6]), 
         .n10375(n10375), .\data_in[6][3] (\data_in[6] [3]), .data_out_10__7__N_114(data_out_10__7__N_114), 
         .n10374(n10374), .\data_in[6][2] (\data_in[6] [2]), .\data_out[0][1] (\data_out[0] [1]), 
         .\data_out[0][3] (\data_out[0] [3]), .n2561(n2561), .n2566(n2566), 
         .n9148(n9148), .n10372(n10372), .\data_in[6][0] (\data_in[6] [0]), 
         .n10371(n10371), .n10370(n10370), .n10369(n10369), .n10367(n10367), 
         .n4430(n4430), .n17585(n17585), .n10631(n10631), .n9631(n9631), 
         .n2568(n2568), .n2564(n2564), .n29(n29), .data_out_5__7__N_931(data_out_5__7__N_931), 
         .data_out_6__6__N_729(data_out_6__6__N_729), .\data_out[2][0] (\data_out[2] [0]), 
         .n16864(n16864), .\delay_counter[0] (delay_counter[0]), .\rand_setpoint[9] (rand_setpoint[9]), 
         .n2567(n2567), .\data_out[3][4] (\data_out[3] [4]), .\data_out[1][6] (\data_out[1] [6]), 
         .\data_out[0][0] (\data_out[0] [0]), .n10366(n10366), .\rand_setpoint[10] (rand_setpoint[10]), 
         .\data_out[1][7] (\data_out[1] [7]), .n2560(n2560), .n2572(n2572), 
         .n10394(n10394), .\data_in[8] ({\data_in[8] }), .n10393(n10393), 
         .n2571(n2571), .n17547(n17547), .tx_transmit_N_2239({tx_transmit_N_2239[7:2], 
         Open_11, Open_12}), .\byte_transmit_counter[7] (byte_transmit_counter[7]), 
         .\byte_transmit_counter[6] (byte_transmit_counter[6]), .n19(n19_adj_2651), 
         .\data_in[4] ({Open_13, Open_14, Open_15, Open_16, Open_17, 
         Open_18, \data_in[4] [1], Open_19}), .\rand_setpoint[11] (rand_setpoint[11]), 
         .\rand_setpoint[12] (rand_setpoint[12]), .n2575(n2575), .\rand_setpoint[13] (rand_setpoint[13]), 
         .n10144(n10144), .\data_in[1] ({Open_20, Open_21, Open_22, 
         Open_23, Open_24, \data_in[1] [2:1], Open_25}), .n6(n6_adj_2616), 
         .\FRAME_MATCHER.next_state[1] (\FRAME_MATCHER.next_state [1]), .n2562(n2562), 
         .n17481(n17481), .n38(n38), .\byte_transmit_counter[5] (byte_transmit_counter[5]), 
         .n10604(n10604), .\data_out_frame2[19][0] (\data_out_frame2[19] [0]), 
         .n10603(n10603), .n10602(n10602), .n10601(n10601), .n10600(n10600), 
         .n10599(n10599), .n10598(n10598), .n2570(n2570), .n8(n8_adj_2613), 
         .n8_adj_3(n8), .n10597(n10597), .\data_out[0][5] (\data_out[0] [5]), 
         .\rand_setpoint[14] (rand_setpoint[14]), .n10649(n10649), .n10652(n10652), 
         .n10655(n10655), .n10659(n10659), .n10662(n10662), .n10671(n10671), 
         .\delay_counter[14] (delay_counter[14]), .\delay_counter[13] (delay_counter[13]), 
         .n10683(n10683), .n10691(n10691), .\data_in[0] ({\data_in[0] [7], 
         Open_26, Open_27, Open_28, Open_29, Open_30, Open_31, Open_32}), 
         .n8_adj_4(n8_adj_2647), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n8_adj_5(n8_adj_2605), .\byte_transmit_counter[3] (byte_transmit_counter[3]), 
         .n8_adj_6(n8_adj_2654), .\byte_transmit_counter[4] (byte_transmit_counter[4]), 
         .n8_adj_7(n8_adj_2611), .\rand_setpoint[15] (rand_setpoint[15]), 
         .\data_out[3][5] (\data_out[3] [5]), .n10596(n10596), .n10595(n10595), 
         .n13415(n13415), .n10594(n10594), .n10391(n10391), .n10438(n10438), 
         .\data_in[14] ({\data_in[14] }), .n10437(n10437), .n10436(n10436), 
         .n10435(n10435), .\data_in[13] ({\data_in[13] }), .n10434(n10434), 
         .n10433(n10433), .n10593(n10593), .n10592(n10592), .n10591(n10591), 
         .data_out_6__2__N_804(data_out_6__2__N_804), .\data_in[9] ({\data_in[9] }), 
         .n10590(n10590), .n10589(n10589), .n10588(n10588), .n10587(n10587), 
         .n10586(n10586), .n10585(n10585), .n10584(n10584), .n10583(n10583), 
         .n10582(n10582), .n10581(n10581), .n10580(n10580), .n10579(n10579), 
         .\data_out_frame2[15] ({\data_out_frame2[15] }), .n10578(n10578), 
         .n10577(n10577), .n10576(n10576), .n10575(n10575), .n10574(n10574), 
         .n10390(n10390), .n10432(n10432), .n10431(n10431), .n10430(n10430), 
         .n10573(n10573), .n10572(n10572), .n10571(n10571), .\data_out_frame2[14] ({\data_out_frame2[14] }), 
         .n10389(n10389), .n10429(n10429), .n10428(n10428), .n10427(n10427), 
         .\data_in[12] ({\data_in[12] }), .n10426(n10426), .n10425(n10425), 
         .n10424(n10424), .n10570(n10570), .n10569(n10569), .n10568(n10568), 
         .n10567(n10567), .n10566(n10566), .n10565(n10565), .n10564(n10564), 
         .n10423(n10423), .n10563(n10563), .n10562(n10562), .n10561(n10561), 
         .n10560(n10560), .n10142(n10142), .n10141(n10141), .n2590(n2590), 
         .n10422(n10422), .n10421(n10421), .n10559(n10559), .\data_out_frame2[6] ({\data_out_frame2[6] }), 
         .\data_out_frame2[7] ({\data_out_frame2[7] }), .\data_out_frame2[5] ({\data_out_frame2[5] }), 
         .n2614({n2615}), .n10140(n10140), .n10364(n10364), .\data_out[1][2] (\data_out[1] [2]), 
         .n2599(n2599), .n2587(n2587), .n2598(n2598), .n10558(n10558), 
         .n10557(n10557), .n10556(n10556), .n10555(n10555), .n10139(n10139), 
         .tx_active(tx_active), .tx_o(tx_o), .tx_o_adj_8(tx_o_adj_2584), 
         .tx_enable(tx_enable), .n7364(n7364), .n10554(n10554), .n10553(n10553), 
         .n10552(n10552), .n10551(n10551), .n10550(n10550), .n10549(n10549), 
         .n10548(n10548), .n10420(n10420), .n10137(n10137), .n10363(n10363), 
         .\data_in[4][7] (\data_in[4] [7]), .n10385(n10385), .\data_in[7][5] (\data_in[7] [5]), 
         .n2593(n2593), .n2597(n2597), .n10135(n10135), .n10134(n10134), 
         .n10133(n10133), .n10132(n10132), .n2595(n2595), .n2589(n2589), 
         .n9054(n9054), .n10130(n10130), .n10129(n10129), .n10547(n10547), 
         .\data_out_frame2[11] ({\data_out_frame2[11] }), .n10419(n10419), 
         .\data_in[11] ({\data_in[11] }), .n10128(n10128), .n10546(n10546), 
         .n2596(n2596), .n2584(n2584), .n10418(n10418), .n10545(n10545), 
         .n10417(n10417), .n10544(n10544), .n10416(n10416), .n10543(n10543), 
         .n10415(n10415), .n10127(n10127), .data_out_5__4__N_959(data_out_5__4__N_959), 
         .n10542(n10542), .n10414(n10414), .n10541(n10541), .n10413(n10413), 
         .n10540(n10540), .n10412(n10412), .n10539(n10539), .\data_out_frame2[10] ({\data_out_frame2[10] }), 
         .n10411(n10411), .\data_in[10] ({\data_in[10] }), .n10126(n10126), 
         .n10538(n10538), .n10537(n10537), .n10410(n10410), .n10536(n10536), 
         .n10409(n10409), .n10535(n10535), .n10408(n10408), .n10125(n10125), 
         .n10534(n10534), .n10533(n10533), .n10407(n10407), .n10532(n10532), 
         .n10406(n10406), .n10531(n10531), .\data_out_frame2[9] ({\data_out_frame2[9] }), 
         .n10530(n10530), .n10405(n10405), .n10529(n10529), .n2591(n2591), 
         .n10528(n10528), .n10527(n10527), .n10124(n10124), .n10526(n10526), 
         .n10525(n10525), .n10123(n10123), .\data_in[4][0] (\data_in[4] [0]), 
         .n10524(n10524), .\data_in[2] ({Open_33, Open_34, Open_35, 
         \data_in[2] [4], Open_36, \data_in[2] [2], Open_37, Open_38}), 
         .n10523(n10523), .\data_out_frame2[8] ({\data_out_frame2[8] }), 
         .n10121(n10121), .n10522(n10522), .n121(n121_adj_2606), .n10521(n10521), 
         .n10520(n10520), .\data_in[3][7] (\data_in[3] [7]), .n2594(n2594), 
         .n9100(n9100), .n2588(n2588), .n2586(n2586), .n10404(n10404), 
         .n10519(n10519), .n10518(n10518), .n10403(n10403), .n10517(n10517), 
         .n10516(n10516), .n10515(n10515), .n10119(n10119), .\data_in[1][4] (\data_in[1] [4]), 
         .n10118(n10118), .\data_in[1][5] (\data_in[1] [5]), .n10402(n10402), 
         .\data_in[3][2] (\data_in[3] [2]), .n119(n119), .\data_in[1][6] (\data_in[1] [6]), 
         .n8529(n8529), .n4(n4_adj_2612), .n10514(n10514), .n10401(n10401), 
         .n10116(n10116), .\data_in[1][7] (\data_in[1] [7]), .n10513(n10513), 
         .n10400(n10400), .n10512(n10512), .n10399(n10399), .n17312(n17312), 
         .n9938(n9938), .\data_in[0][1] (\data_in[0] [1]), .n10114(n10114), 
         .\data_in[2][1] (\data_in[2] [1]), .n10511(n10511), .n10510(n10510), 
         .n10509(n10509), .n10398(n10398), .n10112(n10112), .\data_in[2][3] (\data_in[2] [3]), 
         .n10508(n10508), .n10397(n10397), .n10507(n10507), .n10506(n10506), 
         .n10505(n10505), .n10110(n10110), .\data_in[2][5] (\data_in[2] [5]), 
         .\data_in[2][6] (\data_in[2] [6]), .n1396(n1396), .n10504(n10504), 
         .n10503(n10503), .n10109(n10109), .n10108(n10108), .\data_in[2][7] (\data_in[2] [7]), 
         .\data_in[3][6] (\data_in[3] [6]), .\data_in[3][3] (\data_in[3] [3]), 
         .\data_in[0][4] (\data_in[0] [4]), .n10106(n10106), .\data_in[3][1] (\data_in[3] [1]), 
         .n10105(n10105), .\data_in[0][2] (\data_in[0] [2]), .n10104(n10104), 
         .n63(n63_adj_2642), .\FRAME_MATCHER.next_state_31__N_2026[1] (\FRAME_MATCHER.next_state_31__N_2026 [1]), 
         .n10102(n10102), .\data_in[3][5] (\data_in[3] [5]), .n10101(n10101), 
         .n10100(n10100), .\data_in[4][5] (\data_in[4] [5]), .n10361(n10361), 
         .n2563(n2563), .n10099(n10099), .\data_in[4][2] (\data_in[4] [2]), 
         .n10502(n10502), .n10501(n10501), .n10500(n10500), .n10499(n10499), 
         .n10498(n10498), .n10497(n10497), .n10496(n10496), .n10495(n10495), 
         .n10494(n10494), .n10493(n10493), .n10492(n10492), .n10491(n10491), 
         .\data_in[20] ({\data_in[20] }), .n10490(n10490), .n10489(n10489), 
         .n10488(n10488), .n10487(n10487), .n10486(n10486), .n10485(n10485), 
         .n10484(n10484), .n10483(n10483), .\data_in[19] ({\data_in[19] }), 
         .n10482(n10482), .n10481(n10481), .n10480(n10480), .n10479(n10479), 
         .n10478(n10478), .n10477(n10477), .n10476(n10476), .n10475(n10475), 
         .\data_in[18] ({\data_in[18] }), .n10474(n10474), .n10388(n10388), 
         .\data_in_frame[9][6] (\data_in_frame[9] [6]), .n9419(n9419), .n2573(n2573), 
         .n10473(n10473), .n10472(n10472), .n10471(n10471), .\data_in[0][6] (\data_in[0] [6]), 
         .\data_in[0][5] (\data_in[0] [5]), .n63_adj_9(n63), .n9606(n9606), 
         .n17480(n17480), .n17548(n17548), .n10360(n10360), .n10359(n10359), 
         .n10358(n10358), .n10357(n10357), .n10353(n10353), .n10352(n10352), 
         .n10351(n10351), .n10347(n10347), .\data_in[4][3] (\data_in[4] [3]), 
         .n10470(n10470), .n10469(n10469), .n10468(n10468), .n10467(n10467), 
         .\data_in[17] ({\data_in[17] }), .n10466(n10466), .n10387(n10387), 
         .\data_in[7][7] (\data_in[7] [7]), .n9135(n9135), .\FRAME_MATCHER.next_state[0] (\FRAME_MATCHER.next_state [0]), 
         .n10386(n10386), .\data_in[7][6] (\data_in[7] [6]), .n17092(n17092), 
         .n10465(n10465), .\data_in_frame[7][0] (\data_in_frame[7] [0]), 
         .n9283(n9283), .n6_adj_10(n6_adj_2583), .n16468(n16468), .n10464(n10464), 
         .n10463(n10463), .n10462(n10462), .n10461(n10461), .n10460(n10460), 
         .n10459(n10459), .\data_in[16] ({\data_in[16] }), .n10458(n10458), 
         .n10457(n10457), .n10456(n10456), .n10455(n10455), .n10454(n10454), 
         .n10453(n10453), .n10452(n10452), .n10451(n10451), .\data_in[15] ({\data_in[15] }), 
         .n10396(n10396), .n9937(n9937), .\UART_TRANSMITTER.state_7__N_1749[2] (\UART_TRANSMITTER.state_7__N_1749 [2]), 
         .n9935(n9935), .n9934(n9934), .n9932(n9932), .n8488(n8488), 
         .n96(n96), .n17709(n17709), .n10450(n10450), .n10449(n10449), 
         .n10395(n10395), .n6878(n6878), .n17364(n17364), .n17672(n17672), 
         .n10448(n10448), .n17306(n17306), .\rand_setpoint[24] (rand_setpoint[24]), 
         .\rand_setpoint[25] (rand_setpoint[25]), .n2585(n2585), .\rand_setpoint[26] (rand_setpoint[26]), 
         .\rand_setpoint[27] (rand_setpoint[27]), .n10447(n10447), .n10446(n10446), 
         .\rand_setpoint[28] (rand_setpoint[28]), .\rand_setpoint[29] (rand_setpoint[29]), 
         .n2719({n2720}), .\rand_setpoint[30] (rand_setpoint[30]), .n10445(n10445), 
         .n10444(n10444), .n10443(n10443), .n10442(n10442), .\rand_setpoint[31] (rand_setpoint[31]), 
         .n10441(n10441), .n10440(n10440), .n10439(n10439), .\rand_setpoint[16] (rand_setpoint[16]), 
         .n10044(n10044), .\rand_setpoint[17] (rand_setpoint[17]), .\rand_setpoint[18] (rand_setpoint[18]), 
         .\rand_setpoint[19] (rand_setpoint[19]), .n9051(n9051), .n10043(n10043), 
         .n10039(n10039), .n10038(n10038), .n10034(n10034), .n10033(n10033), 
         .n10032(n10032), .n10031(n10031), .n10027(n10027), .n10026(n10026), 
         .n10025(n10025), .n10024(n10024), .n10023(n10023), .\rand_setpoint[20] (rand_setpoint[20]), 
         .n10022(n10022), .\data_in_frame[6][5] (\data_in_frame[6] [5]), 
         .n10021(n10021), .n10019(n10019), .n10018(n10018), .n10017(n10017), 
         .n10016(n10016), .n10009(n10009), .n10005(n10005), .n10004(n10004), 
         .n10003(n10003), .n9993(n9993), .n9989(n9989), .n9988(n9988), 
         .n9987(n9987), .n9986(n9986), .n9985(n9985), .\rand_setpoint[21] (rand_setpoint[21]), 
         .n9983(n9983), .n9982(n9982), .n9981(n9981), .n9980(n9980), 
         .n9979(n9979), .n9978(n9978), .n9977(n9977), .n9976(n9976), 
         .\rand_setpoint[22] (rand_setpoint[22]), .n9947(n9947), .\rand_setpoint[23] (rand_setpoint[23]), 
         .r_SM_Main({r_SM_Main}), .n10638(n10638), .r_Tx_Data({r_Tx_Data}), 
         .r_Clock_Count({r_Clock_Count}), .n16998(n16998), .n18103(n18103), 
         .n17366(n17366), .n10637(n10637), .n10636(n10636), .n10635(n10635), 
         .n10634(n10634), .n10633(n10633), .n10632(n10632), .n18102(n18102), 
         .n17054(n17054), .r_Bit_Index({r_Bit_Index}), .n16932(n16932), 
         .n16954(n16954), .n16968(n16968), .n17078(n17078), .n18101(n18101), 
         .n17028(n17028), .n18104(n18104), .n9972(n9972), .n10702(n10702), 
         .n17084(n17084), .n17082(n17082), .n17080(n17080), .n17030(n17030), 
         .\r_SM_Main_2__N_2323[1] (r_SM_Main_2__N_2323[1]), .n18098(n18098), 
         .n4_adj_11(n4_adj_2653), .n8517(n8517), .n12(n12_adj_2618), .n9390(n9390), 
         .n16466(n16466), .n10326(n10326), .n10325(n10325), .n10324(n10324), 
         .n10323(n10323), .n7086(n7086), .n7734(n7734), .n13601(n13601), 
         .n1(n1), .n3(n3_adj_2650), .n17757(n17757), .n7080(n7080), 
         .n9796(n9796), .n17950(n17950), .n17356(n17356), .n17952(n17952), 
         .n18010(n18010), .n18054(n18054), .n18097(n18097), .n10245(n10245), 
         .\r_Clock_Count[0]_adj_12 (r_Clock_Count_adj_2666[0]), .r_Bit_Index_adj_35({r_Bit_Index_adj_2667}), 
         .n10625(n10625), .n10346(n10346), .n10008(n10008), .\r_Clock_Count[5]_adj_16 (r_Clock_Count_adj_2666[5]), 
         .n10002(n10002), .\r_Clock_Count[4]_adj_17 (r_Clock_Count_adj_2666[4]), 
         .n9999(n9999), .\r_Clock_Count[3]_adj_18 (r_Clock_Count_adj_2666[3]), 
         .n9996(n9996), .\r_Clock_Count[2]_adj_19 (r_Clock_Count_adj_2666[2]), 
         .n9992(n9992), .\r_Clock_Count[1]_adj_20 (r_Clock_Count_adj_2666[1]), 
         .n10160(n10160), .\r_SM_Main[2]_adj_21 (r_SM_Main_adj_2665[2]), 
         .n10244(n10244), .n316(n316), .n317(n317), .tx2_o(tx2_o), .n318(n318), 
         .n4980(n4980), .n9652(n9652), .n319(n319), .n9922(n9922), .n320(n320), 
         .n321(n321), .tx2_enable(tx2_enable), .n10166(n10166), .r_Bit_Index_adj_36({r_Bit_Index_adj_2661}), 
         .n10194(n10194), .\r_Clock_Count[0]_adj_25 (r_Clock_Count_adj_2660[0]), 
         .n10170(n10170), .rx_data({rx_data}), .n10628(n10628), .n10095(n10095), 
         .\r_Clock_Count[5]_adj_26 (r_Clock_Count_adj_2660[5]), .n10092(n10092), 
         .\r_Clock_Count[4]_adj_27 (r_Clock_Count_adj_2660[4]), .n10089(n10089), 
         .\r_Clock_Count[3]_adj_28 (r_Clock_Count_adj_2660[3]), .n10086(n10086), 
         .\r_Clock_Count[2]_adj_29 (r_Clock_Count_adj_2660[2]), .n10083(n10083), 
         .\r_Clock_Count[1]_adj_30 (r_Clock_Count_adj_2660[1]), .n10643(n10643), 
         .n10644(n10644), .n10645(n10645), .n10646(n10646), .n3_adj_31(n3), 
         .n4_adj_32(n4_adj_2582), .n13597(n13597), .r_Rx_Data(r_Rx_Data), 
         .rx_i(rx_i), .n4_adj_33(n4), .n4958(n4958), .n13880(n13880), 
         .n4_adj_34(n4_adj_2649), .n9933(n9933), .n8567(n8567), .n8562(n8562), 
         .n9646(n9646), .n221(n221), .n222(n222), .n223(n223), .n224(n224), 
         .n225(n225), .n9920(n9920), .n226(n226), .n9942(n9942), .n9941(n9941), 
         .n9940(n9940)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(84[8] 97[4])
    SB_LUT4 blink_counter_2271_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n16392), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2271_add_4_15_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n16485, \UART_TRANSMITTER.state[1] , \UART_TRANSMITTER.state[0] , 
            i_Tx_Byte, n10383, \data_in[7] , CLK_c, \data_out[3][6] , 
            n10382, n10380, \data_in[7][0] , n10379, \data_in[6] , 
            n10378, GND_net, VCC_net, \data_in_frame[8] , n10377, 
            \UART_TRANSMITTER.state[2] , \data_in_frame[5] , n9380, n16, 
            \rand_setpoint[8] , n2565, n2574, \data_out[8] , \data_out_frame2[13] , 
            \data_out_frame2[12] , n9519, \data_out_frame2[18] , \data_in_frame[1][1] , 
            data_out_6__7__N_678, data_out_6__1__N_850, \data_out_frame2[17] , 
            \data_out_frame2[16] , \data_in[5] , rx_data_ready, \data_in_frame[10][6] , 
            n10375, \data_in[6][3] , data_out_10__7__N_114, n10374, 
            \data_in[6][2] , \data_out[0][1] , \data_out[0][3] , n2561, 
            n2566, n9148, n10372, \data_in[6][0] , n10371, n10370, 
            n10369, n10367, n4430, n17585, n10631, n9631, n2568, 
            n2564, n29, data_out_5__7__N_931, data_out_6__6__N_729, 
            \data_out[2][0] , n16864, \delay_counter[0] , \rand_setpoint[9] , 
            n2567, \data_out[3][4] , \data_out[1][6] , \data_out[0][0] , 
            n10366, \rand_setpoint[10] , \data_out[1][7] , n2560, n2572, 
            n10394, \data_in[8] , n10393, n2571, n17547, tx_transmit_N_2239, 
            \byte_transmit_counter[7] , \byte_transmit_counter[6] , n19, 
            \data_in[4] , \rand_setpoint[11] , \rand_setpoint[12] , n2575, 
            \rand_setpoint[13] , n10144, \data_in[1] , n6, \FRAME_MATCHER.next_state[1] , 
            n2562, n17481, n38, \byte_transmit_counter[5] , n10604, 
            \data_out_frame2[19][0] , n10603, n10602, n10601, n10600, 
            n10599, n10598, n2570, n8, n8_adj_3, n10597, \data_out[0][5] , 
            \rand_setpoint[14] , n10649, n10652, n10655, n10659, n10662, 
            n10671, \delay_counter[14] , \delay_counter[13] , n10683, 
            n10691, \data_in[0] , n8_adj_4, \byte_transmit_counter[2] , 
            n8_adj_5, \byte_transmit_counter[3] , n8_adj_6, \byte_transmit_counter[4] , 
            n8_adj_7, \rand_setpoint[15] , \data_out[3][5] , n10596, 
            n10595, n13415, n10594, n10391, n10438, \data_in[14] , 
            n10437, n10436, n10435, \data_in[13] , n10434, n10433, 
            n10593, n10592, n10591, data_out_6__2__N_804, \data_in[9] , 
            n10590, n10589, n10588, n10587, n10586, n10585, n10584, 
            n10583, n10582, n10581, n10580, n10579, \data_out_frame2[15] , 
            n10578, n10577, n10576, n10575, n10574, n10390, n10432, 
            n10431, n10430, n10573, n10572, n10571, \data_out_frame2[14] , 
            n10389, n10429, n10428, n10427, \data_in[12] , n10426, 
            n10425, n10424, n10570, n10569, n10568, n10567, n10566, 
            n10565, n10564, n10423, n10563, n10562, n10561, n10560, 
            n10142, n10141, n2590, n10422, n10421, n10559, \data_out_frame2[6] , 
            \data_out_frame2[7] , \data_out_frame2[5] , n2614, n10140, 
            n10364, \data_out[1][2] , n2599, n2587, n2598, n10558, 
            n10557, n10556, n10555, n10139, tx_active, tx_o, tx_o_adj_8, 
            tx_enable, n7364, n10554, n10553, n10552, n10551, n10550, 
            n10549, n10548, n10420, n10137, n10363, \data_in[4][7] , 
            n10385, \data_in[7][5] , n2593, n2597, n10135, n10134, 
            n10133, n10132, n2595, n2589, n9054, n10130, n10129, 
            n10547, \data_out_frame2[11] , n10419, \data_in[11] , n10128, 
            n10546, n2596, n2584, n10418, n10545, n10417, n10544, 
            n10416, n10543, n10415, n10127, data_out_5__4__N_959, 
            n10542, n10414, n10541, n10413, n10540, n10412, n10539, 
            \data_out_frame2[10] , n10411, \data_in[10] , n10126, n10538, 
            n10537, n10410, n10536, n10409, n10535, n10408, n10125, 
            n10534, n10533, n10407, n10532, n10406, n10531, \data_out_frame2[9] , 
            n10530, n10405, n10529, n2591, n10528, n10527, n10124, 
            n10526, n10525, n10123, \data_in[4][0] , n10524, \data_in[2] , 
            n10523, \data_out_frame2[8] , n10121, n10522, n121, n10521, 
            n10520, \data_in[3][7] , n2594, n9100, n2588, n2586, 
            n10404, n10519, n10518, n10403, n10517, n10516, n10515, 
            n10119, \data_in[1][4] , n10118, \data_in[1][5] , n10402, 
            \data_in[3][2] , n119, \data_in[1][6] , n8529, n4, n10514, 
            n10401, n10116, \data_in[1][7] , n10513, n10400, n10512, 
            n10399, n17312, n9938, \data_in[0][1] , n10114, \data_in[2][1] , 
            n10511, n10510, n10509, n10398, n10112, \data_in[2][3] , 
            n10508, n10397, n10507, n10506, n10505, n10110, \data_in[2][5] , 
            \data_in[2][6] , n1396, n10504, n10503, n10109, n10108, 
            \data_in[2][7] , \data_in[3][6] , \data_in[3][3] , \data_in[0][4] , 
            n10106, \data_in[3][1] , n10105, \data_in[0][2] , n10104, 
            n63, \FRAME_MATCHER.next_state_31__N_2026[1] , n10102, \data_in[3][5] , 
            n10101, n10100, \data_in[4][5] , n10361, n2563, n10099, 
            \data_in[4][2] , n10502, n10501, n10500, n10499, n10498, 
            n10497, n10496, n10495, n10494, n10493, n10492, n10491, 
            \data_in[20] , n10490, n10489, n10488, n10487, n10486, 
            n10485, n10484, n10483, \data_in[19] , n10482, n10481, 
            n10480, n10479, n10478, n10477, n10476, n10475, \data_in[18] , 
            n10474, n10388, \data_in_frame[9][6] , n9419, n2573, n10473, 
            n10472, n10471, \data_in[0][6] , \data_in[0][5] , n63_adj_9, 
            n9606, n17480, n17548, n10360, n10359, n10358, n10357, 
            n10353, n10352, n10351, n10347, \data_in[4][3] , n10470, 
            n10469, n10468, n10467, \data_in[17] , n10466, n10387, 
            \data_in[7][7] , n9135, \FRAME_MATCHER.next_state[0] , n10386, 
            \data_in[7][6] , n17092, n10465, \data_in_frame[7][0] , 
            n9283, n6_adj_10, n16468, n10464, n10463, n10462, n10461, 
            n10460, n10459, \data_in[16] , n10458, n10457, n10456, 
            n10455, n10454, n10453, n10452, n10451, \data_in[15] , 
            n10396, n9937, \UART_TRANSMITTER.state_7__N_1749[2] , n9935, 
            n9934, n9932, n8488, n96, n17709, n10450, n10449, 
            n10395, n6878, n17364, n17672, n10448, n17306, \rand_setpoint[24] , 
            \rand_setpoint[25] , n2585, \rand_setpoint[26] , \rand_setpoint[27] , 
            n10447, n10446, \rand_setpoint[28] , \rand_setpoint[29] , 
            n2719, \rand_setpoint[30] , n10445, n10444, n10443, n10442, 
            \rand_setpoint[31] , n10441, n10440, n10439, \rand_setpoint[16] , 
            n10044, \rand_setpoint[17] , \rand_setpoint[18] , \rand_setpoint[19] , 
            n9051, n10043, n10039, n10038, n10034, n10033, n10032, 
            n10031, n10027, n10026, n10025, n10024, n10023, \rand_setpoint[20] , 
            n10022, \data_in_frame[6][5] , n10021, n10019, n10018, 
            n10017, n10016, n10009, n10005, n10004, n10003, n9993, 
            n9989, n9988, n9987, n9986, n9985, \rand_setpoint[21] , 
            n9983, n9982, n9981, n9980, n9979, n9978, n9977, n9976, 
            \rand_setpoint[22] , n9947, \rand_setpoint[23] , r_SM_Main, 
            n10638, r_Tx_Data, r_Clock_Count, n16998, n18103, n17366, 
            n10637, n10636, n10635, n10634, n10633, n10632, n18102, 
            n17054, r_Bit_Index, n16932, n16954, n16968, n17078, 
            n18101, n17028, n18104, n9972, n10702, n17084, n17082, 
            n17080, n17030, \r_SM_Main_2__N_2323[1] , n18098, n4_adj_11, 
            n8517, n12, n9390, n16466, n10326, n10325, n10324, 
            n10323, n7086, n7734, n13601, n1, n3, n17757, n7080, 
            n9796, n17950, n17356, n17952, n18010, n18054, n18097, 
            n10245, \r_Clock_Count[0]_adj_12 , r_Bit_Index_adj_35, n10625, 
            n10346, n10008, \r_Clock_Count[5]_adj_16 , n10002, \r_Clock_Count[4]_adj_17 , 
            n9999, \r_Clock_Count[3]_adj_18 , n9996, \r_Clock_Count[2]_adj_19 , 
            n9992, \r_Clock_Count[1]_adj_20 , n10160, \r_SM_Main[2]_adj_21 , 
            n10244, n316, n317, tx2_o, n318, n4980, n9652, n319, 
            n9922, n320, n321, tx2_enable, n10166, r_Bit_Index_adj_36, 
            n10194, \r_Clock_Count[0]_adj_25 , n10170, rx_data, n10628, 
            n10095, \r_Clock_Count[5]_adj_26 , n10092, \r_Clock_Count[4]_adj_27 , 
            n10089, \r_Clock_Count[3]_adj_28 , n10086, \r_Clock_Count[2]_adj_29 , 
            n10083, \r_Clock_Count[1]_adj_30 , n10643, n10644, n10645, 
            n10646, n3_adj_31, n4_adj_32, n13597, r_Rx_Data, rx_i, 
            n4_adj_33, n4958, n13880, n4_adj_34, n9933, n8567, n8562, 
            n9646, n221, n222, n223, n224, n225, n9920, n226, 
            n9942, n9941, n9940) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n16485;
    output \UART_TRANSMITTER.state[1] ;
    output \UART_TRANSMITTER.state[0] ;
    output [7:0]i_Tx_Byte;
    input n10383;
    output [7:0]\data_in[7] ;
    input CLK_c;
    output \data_out[3][6] ;
    input n10382;
    input n10380;
    output \data_in[7][0] ;
    input n10379;
    output [7:0]\data_in[6] ;
    input n10378;
    input GND_net;
    input VCC_net;
    output [7:0]\data_in_frame[8] ;
    input n10377;
    output \UART_TRANSMITTER.state[2] ;
    output [7:0]\data_in_frame[5] ;
    output n9380;
    input n16;
    input \rand_setpoint[8] ;
    output n2565;
    output n2574;
    output [7:0]\data_out[8] ;
    output [7:0]\data_out_frame2[13] ;
    output [7:0]\data_out_frame2[12] ;
    output n9519;
    output [7:0]\data_out_frame2[18] ;
    output \data_in_frame[1][1] ;
    output data_out_6__7__N_678;
    output data_out_6__1__N_850;
    output [7:0]\data_out_frame2[17] ;
    output [7:0]\data_out_frame2[16] ;
    output [7:0]\data_in[5] ;
    output rx_data_ready;
    output \data_in_frame[10][6] ;
    input n10375;
    output \data_in[6][3] ;
    output data_out_10__7__N_114;
    input n10374;
    output \data_in[6][2] ;
    output \data_out[0][1] ;
    output \data_out[0][3] ;
    output n2561;
    output n2566;
    output n9148;
    input n10372;
    output \data_in[6][0] ;
    input n10371;
    input n10370;
    input n10369;
    input n10367;
    output n4430;
    input n17585;
    input n10631;
    output n9631;
    output n2568;
    output n2564;
    output n29;
    output data_out_5__7__N_931;
    output data_out_6__6__N_729;
    output \data_out[2][0] ;
    input n16864;
    output \delay_counter[0] ;
    input \rand_setpoint[9] ;
    output n2567;
    output \data_out[3][4] ;
    output \data_out[1][6] ;
    output \data_out[0][0] ;
    input n10366;
    input \rand_setpoint[10] ;
    output \data_out[1][7] ;
    output n2560;
    output n2572;
    input n10394;
    output [7:0]\data_in[8] ;
    input n10393;
    output n2571;
    input n17547;
    output [7:0]tx_transmit_N_2239;
    output \byte_transmit_counter[7] ;
    output \byte_transmit_counter[6] ;
    input n19;
    output [7:0]\data_in[4] ;
    input \rand_setpoint[11] ;
    input \rand_setpoint[12] ;
    output n2575;
    input \rand_setpoint[13] ;
    input n10144;
    output [7:0]\data_in[1] ;
    input n6;
    output \FRAME_MATCHER.next_state[1] ;
    output n2562;
    input n17481;
    input n38;
    output \byte_transmit_counter[5] ;
    input n10604;
    output \data_out_frame2[19][0] ;
    input n10603;
    input n10602;
    input n10601;
    input n10600;
    input n10599;
    input n10598;
    output n2570;
    input n8;
    input n8_adj_3;
    input n10597;
    output \data_out[0][5] ;
    input \rand_setpoint[14] ;
    input n10649;
    input n10652;
    input n10655;
    input n10659;
    input n10662;
    input n10671;
    output \delay_counter[14] ;
    output \delay_counter[13] ;
    input n10683;
    input n10691;
    output [7:0]\data_in[0] ;
    input n8_adj_4;
    output \byte_transmit_counter[2] ;
    input n8_adj_5;
    output \byte_transmit_counter[3] ;
    input n8_adj_6;
    output \byte_transmit_counter[4] ;
    input n8_adj_7;
    input \rand_setpoint[15] ;
    output \data_out[3][5] ;
    input n10596;
    input n10595;
    output n13415;
    input n10594;
    input n10391;
    input n10438;
    output [7:0]\data_in[14] ;
    input n10437;
    input n10436;
    input n10435;
    output [7:0]\data_in[13] ;
    input n10434;
    input n10433;
    input n10593;
    input n10592;
    input n10591;
    output data_out_6__2__N_804;
    output [7:0]\data_in[9] ;
    input n10590;
    input n10589;
    input n10588;
    input n10587;
    input n10586;
    input n10585;
    input n10584;
    input n10583;
    input n10582;
    input n10581;
    input n10580;
    input n10579;
    output [7:0]\data_out_frame2[15] ;
    input n10578;
    input n10577;
    input n10576;
    input n10575;
    input n10574;
    input n10390;
    input n10432;
    input n10431;
    input n10430;
    input n10573;
    input n10572;
    input n10571;
    output [7:0]\data_out_frame2[14] ;
    input n10389;
    input n10429;
    input n10428;
    input n10427;
    output [7:0]\data_in[12] ;
    input n10426;
    input n10425;
    input n10424;
    input n10570;
    input n10569;
    input n10568;
    input n10567;
    input n10566;
    input n10565;
    input n10564;
    input n10423;
    input n10563;
    input n10562;
    input n10561;
    input n10560;
    input n10142;
    input n10141;
    output n2590;
    input n10422;
    input n10421;
    input n10559;
    output [7:0]\data_out_frame2[6] ;
    output [7:0]\data_out_frame2[7] ;
    output [7:0]\data_out_frame2[5] ;
    output [0:0]n2614;
    input n10140;
    input n10364;
    output \data_out[1][2] ;
    output n2599;
    output n2587;
    output n2598;
    input n10558;
    input n10557;
    input n10556;
    input n10555;
    input n10139;
    output tx_active;
    output tx_o;
    output tx_o_adj_8;
    output tx_enable;
    output n7364;
    input n10554;
    input n10553;
    input n10552;
    input n10551;
    input n10550;
    input n10549;
    input n10548;
    input n10420;
    input n10137;
    input n10363;
    output \data_in[4][7] ;
    input n10385;
    output \data_in[7][5] ;
    output n2593;
    output n2597;
    input n10135;
    input n10134;
    input n10133;
    input n10132;
    output n2595;
    output n2589;
    output n9054;
    input n10130;
    input n10129;
    input n10547;
    output [7:0]\data_out_frame2[11] ;
    input n10419;
    output [7:0]\data_in[11] ;
    input n10128;
    input n10546;
    output n2596;
    output n2584;
    input n10418;
    input n10545;
    input n10417;
    input n10544;
    input n10416;
    input n10543;
    input n10415;
    input n10127;
    output data_out_5__4__N_959;
    input n10542;
    input n10414;
    input n10541;
    input n10413;
    input n10540;
    input n10412;
    input n10539;
    output [7:0]\data_out_frame2[10] ;
    input n10411;
    output [7:0]\data_in[10] ;
    input n10126;
    input n10538;
    input n10537;
    input n10410;
    input n10536;
    input n10409;
    input n10535;
    input n10408;
    input n10125;
    input n10534;
    input n10533;
    input n10407;
    input n10532;
    input n10406;
    input n10531;
    output [7:0]\data_out_frame2[9] ;
    input n10530;
    input n10405;
    input n10529;
    output n2591;
    input n10528;
    input n10527;
    input n10124;
    input n10526;
    input n10525;
    input n10123;
    output \data_in[4][0] ;
    input n10524;
    output [7:0]\data_in[2] ;
    input n10523;
    output [7:0]\data_out_frame2[8] ;
    input n10121;
    input n10522;
    output n121;
    input n10521;
    input n10520;
    output \data_in[3][7] ;
    output n2594;
    output n9100;
    output n2588;
    output n2586;
    input n10404;
    input n10519;
    input n10518;
    input n10403;
    input n10517;
    input n10516;
    input n10515;
    input n10119;
    output \data_in[1][4] ;
    input n10118;
    output \data_in[1][5] ;
    input n10402;
    output \data_in[3][2] ;
    output n119;
    output \data_in[1][6] ;
    output n8529;
    output n4;
    input n10514;
    input n10401;
    input n10116;
    output \data_in[1][7] ;
    input n10513;
    input n10400;
    input n10512;
    input n10399;
    input n17312;
    input n9938;
    output \data_in[0][1] ;
    input n10114;
    output \data_in[2][1] ;
    input n10511;
    input n10510;
    input n10509;
    input n10398;
    input n10112;
    output \data_in[2][3] ;
    input n10508;
    input n10397;
    input n10507;
    input n10506;
    input n10505;
    input n10110;
    output \data_in[2][5] ;
    output \data_in[2][6] ;
    output n1396;
    input n10504;
    input n10503;
    input n10109;
    input n10108;
    output \data_in[2][7] ;
    output \data_in[3][6] ;
    output \data_in[3][3] ;
    output \data_in[0][4] ;
    input n10106;
    output \data_in[3][1] ;
    input n10105;
    output \data_in[0][2] ;
    input n10104;
    output n63;
    output \FRAME_MATCHER.next_state_31__N_2026[1] ;
    input n10102;
    output \data_in[3][5] ;
    input n10101;
    input n10100;
    output \data_in[4][5] ;
    input n10361;
    output n2563;
    input n10099;
    output \data_in[4][2] ;
    input n10502;
    input n10501;
    input n10500;
    input n10499;
    input n10498;
    input n10497;
    input n10496;
    input n10495;
    input n10494;
    input n10493;
    input n10492;
    input n10491;
    output [7:0]\data_in[20] ;
    input n10490;
    input n10489;
    input n10488;
    input n10487;
    input n10486;
    input n10485;
    input n10484;
    input n10483;
    output [7:0]\data_in[19] ;
    input n10482;
    input n10481;
    input n10480;
    input n10479;
    input n10478;
    input n10477;
    input n10476;
    input n10475;
    output [7:0]\data_in[18] ;
    input n10474;
    input n10388;
    output \data_in_frame[9][6] ;
    output n9419;
    output n2573;
    input n10473;
    input n10472;
    input n10471;
    output \data_in[0][6] ;
    output \data_in[0][5] ;
    output n63_adj_9;
    output n9606;
    input n17480;
    input n17548;
    input n10360;
    input n10359;
    input n10358;
    input n10357;
    input n10353;
    input n10352;
    input n10351;
    input n10347;
    output \data_in[4][3] ;
    input n10470;
    input n10469;
    input n10468;
    input n10467;
    output [7:0]\data_in[17] ;
    input n10466;
    input n10387;
    output \data_in[7][7] ;
    output n9135;
    output \FRAME_MATCHER.next_state[0] ;
    input n10386;
    output \data_in[7][6] ;
    input n17092;
    input n10465;
    output \data_in_frame[7][0] ;
    output n9283;
    output n6_adj_10;
    output n16468;
    input n10464;
    input n10463;
    input n10462;
    input n10461;
    input n10460;
    input n10459;
    output [7:0]\data_in[16] ;
    input n10458;
    input n10457;
    input n10456;
    input n10455;
    input n10454;
    input n10453;
    input n10452;
    input n10451;
    output [7:0]\data_in[15] ;
    input n10396;
    input n9937;
    output \UART_TRANSMITTER.state_7__N_1749[2] ;
    input n9935;
    input n9934;
    input n9932;
    output n8488;
    output n96;
    output n17709;
    input n10450;
    input n10449;
    input n10395;
    output n6878;
    input n17364;
    output n17672;
    input n10448;
    output n17306;
    input \rand_setpoint[24] ;
    input \rand_setpoint[25] ;
    output n2585;
    input \rand_setpoint[26] ;
    input \rand_setpoint[27] ;
    input n10447;
    input n10446;
    input \rand_setpoint[28] ;
    input \rand_setpoint[29] ;
    output [0:0]n2719;
    input \rand_setpoint[30] ;
    input n10445;
    input n10444;
    input n10443;
    input n10442;
    input \rand_setpoint[31] ;
    input n10441;
    input n10440;
    input n10439;
    input \rand_setpoint[16] ;
    input n10044;
    input \rand_setpoint[17] ;
    input \rand_setpoint[18] ;
    input \rand_setpoint[19] ;
    output n9051;
    input n10043;
    input n10039;
    input n10038;
    input n10034;
    input n10033;
    input n10032;
    input n10031;
    input n10027;
    input n10026;
    input n10025;
    input n10024;
    input n10023;
    input \rand_setpoint[20] ;
    input n10022;
    output \data_in_frame[6][5] ;
    input n10021;
    input n10019;
    input n10018;
    input n10017;
    input n10016;
    input n10009;
    input n10005;
    input n10004;
    input n10003;
    input n9993;
    input n9989;
    input n9988;
    input n9987;
    input n9986;
    input n9985;
    input \rand_setpoint[21] ;
    input n9983;
    input n9982;
    input n9981;
    input n9980;
    input n9979;
    input n9978;
    input n9977;
    input n9976;
    input \rand_setpoint[22] ;
    input n9947;
    input \rand_setpoint[23] ;
    output [2:0]r_SM_Main;
    input n10638;
    output [7:0]r_Tx_Data;
    output [8:0]r_Clock_Count;
    input n16998;
    output n18103;
    input n17366;
    input n10637;
    input n10636;
    input n10635;
    input n10634;
    input n10633;
    input n10632;
    output n18102;
    input n17054;
    output [2:0]r_Bit_Index;
    input n16932;
    input n16954;
    input n16968;
    input n17078;
    output n18101;
    input n17028;
    output n18104;
    input n9972;
    input n10702;
    input n17084;
    input n17082;
    input n17080;
    input n17030;
    output \r_SM_Main_2__N_2323[1] ;
    output n18098;
    output n4_adj_11;
    output n8517;
    output n12;
    output n9390;
    output n16466;
    input n10326;
    input n10325;
    input n10324;
    input n10323;
    output n7086;
    output n7734;
    output n13601;
    input n1;
    output n3;
    output n17757;
    output n7080;
    output n9796;
    output n17950;
    input n17356;
    output n17952;
    output n18010;
    output n18054;
    output n18097;
    input n10245;
    output \r_Clock_Count[0]_adj_12 ;
    output [2:0]r_Bit_Index_adj_35;
    input n10625;
    input n10346;
    input n10008;
    output \r_Clock_Count[5]_adj_16 ;
    input n10002;
    output \r_Clock_Count[4]_adj_17 ;
    input n9999;
    output \r_Clock_Count[3]_adj_18 ;
    input n9996;
    output \r_Clock_Count[2]_adj_19 ;
    input n9992;
    output \r_Clock_Count[1]_adj_20 ;
    input n10160;
    output \r_SM_Main[2]_adj_21 ;
    output n10244;
    output n316;
    output n317;
    output tx2_o;
    output n318;
    output n4980;
    output n9652;
    output n319;
    output n9922;
    output n320;
    output n321;
    output tx2_enable;
    input n10166;
    output [2:0]r_Bit_Index_adj_36;
    input n10194;
    output \r_Clock_Count[0]_adj_25 ;
    input n10170;
    output [7:0]rx_data;
    input n10628;
    input n10095;
    output \r_Clock_Count[5]_adj_26 ;
    input n10092;
    output \r_Clock_Count[4]_adj_27 ;
    input n10089;
    output \r_Clock_Count[3]_adj_28 ;
    input n10086;
    output \r_Clock_Count[2]_adj_29 ;
    input n10083;
    output \r_Clock_Count[1]_adj_30 ;
    input n10643;
    input n10644;
    input n10645;
    input n10646;
    output n3_adj_31;
    output n4_adj_32;
    output n13597;
    output r_Rx_Data;
    input rx_i;
    output n4_adj_33;
    output n4958;
    output n13880;
    output n4_adj_34;
    input n9933;
    output n8567;
    output n8562;
    output n9646;
    output n221;
    output n222;
    output n223;
    output n224;
    output n225;
    output n9920;
    output n226;
    input n9942;
    input n9941;
    input n9940;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n7428, n16870, data_out_7__5__N_543, n17578, n17641, n9276, 
        n10381;
    wire [7:0]\data_in[7]_c ;   // coms.v(382[12:19])
    wire [7:0]\data_in_frame[9] ;   // coms.v(383[12:25])
    
    wire n17488, n10259;
    wire [7:0]\data_in_frame[1] ;   // coms.v(383[12:25])
    
    wire n10255, n10252;
    wire [7:0]\data_out[5] ;   // coms.v(21[11:19])
    
    wire n8634, n17457, n17623;
    wire [7:0]\data_in_frame[7] ;   // coms.v(383[12:25])
    
    wire n17473, data_out_7__1__N_626, n8926, n17916;
    wire [7:0]\data_out[6] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[7] ;   // coms.v(21[11:19])
    wire [7:0]byte_transmit_counter;   // coms.v(19[11:32])
    
    wire n5, n10311;
    wire [7:0]\data_in_frame[3] ;   // coms.v(383[12:25])
    
    wire n8666, n17519, n9204, n9365, n8695, n17430, n22, n17605;
    wire [7:0]\data_in_frame[6] ;   // coms.v(383[12:25])
    
    wire n20, n9208, n24, n9355, n8645, data_out_7__7__N_519, n18017;
    wire [0:0]n2019;
    
    wire n17412, n17594, n23, n9087;
    wire [7:0]\data_in_frame[4] ;   // coms.v(383[12:25])
    
    wire n17513, n10249, n18474;
    wire [7:0]byte_transmit_counter2;   // coms.v(413[12:34])
    
    wire n17836;
    wire [7:0]n37;
    
    wire n9605, n9900, n8812, n10242, data_out_7__2__N_574, data_out_10__2__N_179;
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    
    wire n10131;
    wire [7:0]\data_out_frame2[19] ;   // coms.v(384[12:27])
    
    wire n18468, n10239, n10236, n17445, n18471, n10232;
    wire [7:0]\data_in[6]_c ;   // coms.v(382[12:19])
    
    wire n10365, data_out_6__3__N_788;
    wire [7:0]\data_in_frame[10] ;   // coms.v(383[12:25])
    
    wire n8995, n10, n9131, n17418, n17420, data_out_5__5__N_950, 
        n8767, n10308, n10229;
    wire [7:0]\data_in_frame[0] ;   // coms.v(383[12:25])
    
    wire n10226, n8964, n17525, n17415, n9043, n8886, n17535, 
        n16856, n10376, n10222, data_out_10__5__N_132;
    wire [7:0]\data_out[10] ;   // coms.v(21[11:19])
    
    wire data_out_7__6__N_530, n17504, n9240, n17537, n8777, n8056, 
        n17544, n19_c, n10136, n17955, n5_adj_2425, n18456, n10373, 
        n10219, n10368;
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    
    wire n10138, n17482, data_out_10__4__N_147, n10216, tx_active_prev, 
        n17339, tx_transmit;
    wire [0:0]n1774;
    
    wire n9518;
    wire [0:0]n1809;
    wire [0:0]n1844;
    wire [0:0]n1879;
    wire [0:0]n1914;
    wire [0:0]n1949;
    wire [0:0]n1984;
    wire [0:0]n2054;
    wire [0:0]n2089;
    wire [0:0]n2124;
    wire [0:0]n2159;
    wire [0:0]n2194;
    wire [0:0]n2229;
    wire [0:0]n2264;
    wire [0:0]n2299;
    wire [0:0]n2334;
    wire [0:0]n2369;
    wire [0:0]n2404;
    wire [0:0]n2439;
    
    wire data_out_7__4__N_556;
    wire [0:0]n2474;
    wire [0:0]n2509;
    wire [0:0]n2544;
    wire [0:0]n2579;
    wire [0:0]n3203;
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    
    wire n9685;
    wire [7:0]\data_out_frame2[0] ;   // coms.v(384[12:27])
    
    wire n10213, n17214;
    wire [31:0]\FRAME_MATCHER.state ;   // coms.v(422[11:16])
    
    wire n1_c, n6_c, n17587, n23_adj_2426;
    wire [14:0]n7260;
    wire [14:0]delay_counter;   // coms.v(266[12:25])
    
    wire n16314, n10210, n17538, n21, n18012, n16309, n16306, 
        n16307, n20_adj_2427, n10_adj_2428, n17611, n17659, n17918, 
        n17499, n8674, n9324, n11, n12_c, n18444, n9144, n6_adj_2429, 
        n9151, n17588, n17433, n17590, n16315, n10196, n9, n8_c, 
        n18447, n10188, n10305, n17647, n8890, n17648, data_out_10__3__N_163, 
        n16310, n17644;
    wire [7:0]\data_in_frame[2] ;   // coms.v(383[12:25])
    
    wire n9317, data_out_6__3__N_781, n17921, n16313, n8600, n17582, 
        n18, n9176, n10_adj_2430, n17536, n28, n17635, n17922, 
        n16356, n16355, n9254, n8725, n16308, n10148, n17485, 
        n17931, n18011, n16312, n16305, data_out_7__4__N_550, n17592, 
        n26, n17925, n18372, n6_adj_2432, n18082, n18375, n17773, 
        n17779, n18432, n10622, n10619, n10143;
    wire [7:0]\data_in[4]_c ;   // coms.v(382[12:19])
    
    wire n17541, n27, n10614, n10611, n10608, n16354, n10350, 
        n10356, n25, n6_adj_2436, n18074, n18435, n14631, n142, 
        n9671, n17465, n17906, n9674, n1_adj_2437, n18459, n31, 
        n5_adj_2438, n136, n17400, n10663, n10314, n10262, n10674, 
        n10675, n10676, n10071, n10068, n10065, n10680, n10059, 
        n10056, n10686, n10050, n10047, n10042, n10037, n16858, 
        n10302, n1_adj_2443, n157, data_out_6__7__N_675, n17928, n9677, 
        n5_adj_2444, n97, n16_adj_2445, n17949, n149;
    wire [0:0]n2649;
    
    wire n19_adj_2446, n8550, n17556, n17492, data_out_10__7__N_101, 
        n10392, n17941, n5_adj_2447, n18396, n17620, n17510, n17638, 
        data_out_9__1__N_462, n8950, n8922, data_out_9__2__N_446, n18094, 
        n18095, n16353, n16352, n16311, n6_adj_2448, data_out_9__3__N_430, 
        n9306, n8867, n17406, n12_adj_2449, n8687, n10_adj_2450, 
        n8064, n17470, n17532, n17534, n18426, n6_adj_2451, n8062, 
        n8751, n20_adj_2452, n11_adj_2453, n17522, n24_adj_2454, n2, 
        n18089, n18429, n17424, n1_adj_2455;
    wire [2:0]r_SM_Main_2__N_2326;
    
    wire data_out_10__1__N_196, n9039, n16351;
    wire [7:0]tx_transmit_N_2239_c;
    
    wire n17349, data_out_10__0__N_259, n2839, n8874, n8_adj_2459, 
        n2604, n11_adj_2460, n17529, n22_adj_2461, n8658, n17575, 
        n9103, n23_adj_2462, n18084, n17785, n17788, n18420, n5_adj_2463, 
        n6_adj_2464, n18076, n18423, n21_adj_2465, n6_adj_2466;
    wire [7:0]\data_in[3] ;   // coms.v(382[12:19])
    
    wire n10103, n251, data_out_9__7__N_323;
    wire [7:0]\data_out[9] ;   // coms.v(21[11:19])
    
    wire n18093, n18092, n18399, n17533, n10122;
    wire [7:0]\data_in[0]_c ;   // coms.v(382[12:19])
    
    wire n10107, n6_adj_2467, n10111, n9345, data_out_9__6__N_386, 
        n9939, n8061, n18_adj_2468, n8857, n26_adj_2469, n10384, 
        n10120;
    wire [7:0]\data_in[1]_c ;   // coms.v(382[12:19])
    
    wire n8970, n17600, n17387, n17467, n30, n10113, n10_adj_2470, 
        n17409, n17618, n17442, n17507, n1314, n16350, n17;
    wire [7:0]\data_in[2]_c ;   // coms.v(382[12:19])
    
    wire n10115, n81, n9662, data_out_9__5__N_401, n10117, n16450, 
        n9665, n9668, n8486, n17619, n9680, data_out_9__4__N_414, 
        n17753, n17755, n9091, n17398, n15927, n9984, data_out_6__5__N_752, 
        n17454, n8572, n18009, n17815, n17818, n17824, n17827, 
        n18366, n17697, n12_adj_2472, n17765, n17218, n18008, n17656, 
        n18105, n8556, n17715, n17516, n8976, n6_adj_2473, n8_adj_2474, 
        n18369, n28_adj_2475, n17216, n17833, n18360, n18390, n18393, 
        data_out_9__0__N_475, n8559, n18091, n2_adj_2476, data_out_10__6__N_118, 
        n5_adj_2477, n6_adj_2478, n17743, n18414, n17550, n8460, 
        n7, n17745, n17649;
    wire [7:0]\data_out_frame2[20] ;   // coms.v(384[12:27])
    
    wire n17490, n17540, n17593, n17543, n17545, n17584, n4_adj_2480, 
        n10342, n10266, n10269, n10272, n10276, n10279, n10333, 
        n10330, n10286, n17553, n5_adj_2481, n17943, n17626, n17608, 
        n17662, n12_adj_2482, n17665, n17650, n18096, n17559, n17629, 
        n2_adj_2483, n18090, n1_adj_2484, n18417, n17794, n17797, 
        n18408, n16_adj_2485, n18088, n17_adj_2486, n9219, n8063, 
        n2_adj_2487, n5_adj_2488, n17911, n9349, n30_adj_2489, n9334, 
        n17476, n5_adj_2490, n17937, n9368, n25_adj_2491, n9163, 
        n17602, n12_adj_2492, n2600, n10_adj_2493, n9279, n2601, 
        n11_adj_2494, n18080, n5_adj_2495, n6_adj_2496, n2605, n10_adj_2498, 
        n5_adj_2499, n2607, n2602, n9_adj_2500, n9058, tx2_transmit_N_2287, 
        n17936, n5_adj_2501, n18086, n6_adj_2502, n8989, n5_adj_2503, 
        n17478, n6_adj_2504, n17591, n2603, n17569, n10_adj_2505, 
        n2606, n17428, n14, n6_adj_2506, n18078, n18411, n17325, 
        n17632, n9_adj_2507, n17403, n17614, n22_adj_2508, n9186, 
        n9936, n5_adj_2509, n10289, n10293, n10296, n10299, n134, 
        n18603, n22_adj_2510;
    wire [7:0]tx2_data;   // coms.v(416[13:21])
    
    wire n18606, n113, n17668, n9195, n8_adj_2511, n18600, n4_adj_2512, 
        n16_adj_2513, n17_adj_2514, n18588, n5_adj_2515, n18016, n17741, 
        n8_adj_2516, n93, n18582, n18015, n25_adj_2517, n18501, 
        n18576, n18363, n45_adj_2518, n18579, n18073, n8_adj_2519, 
        n22_adj_2520, n18555, n22_adj_2521, n46, n18570, n1_adj_2522, 
        n18378, n18014, n18384, n18387, n18564, n18537, n22_adj_2523, 
        n44_adj_2524, n18531, n22_adj_2525, n15, n18558, n18071, 
        n8_adj_2526, n18513, n22_adj_2527, n18552, n18546, n17803, 
        n18072, n18381, n8_adj_2528, n18540, n18489, n22_adj_2529, 
        n17806, n9328, n18534, n18528, n18069, n22_adj_2530, n18522, 
        n8_adj_2531, n18070, n10_adj_2532, n18516, n14_adj_2533, n6_adj_2534, 
        n18510, n18067, n8_adj_2535, n8953, n18068, n18504, n10_adj_2536, 
        n18064, n8_adj_2537, n18065, n18405, n18060, n8_adj_2538, 
        n18061, n18498, n18062, n17957, n8_adj_2539, n18063, n18492, 
        n17962, n18486, n17389, data_out_6__1__N_849, n17964, n18480, 
        data_out_6__2__N_803, n17966, data_out_5__3__N_964, n17967, 
        n16411, n16410, n16409, n17970, n10020, n16408, n17972, 
        n16407, n17974, n16406, n17438, n17653, n17976, n17566, 
        n16405, data_out_6__4__N_765, n17654, n17693;
    wire [0:0]n2250;
    wire [0:0]n2215;
    
    wire data_out_6__3__N_785;
    wire [0:0]n2180;
    
    wire n67, n13530, n19_adj_2540, n16318, n16317, n18402;
    wire [0:0]n2145;
    
    wire n6_adj_2541, n12_adj_2542, n9028, n4_adj_2543, n18_adj_2544, 
        n9656, n16316, n9658, n18_adj_2545, n17562, n16_adj_2546, 
        n20_adj_2547, n4_adj_2548;
    wire [0:0]n2040;
    
    wire n12_adj_2549, n6_adj_2550;
    
    assign tx_o = tx_o_adj_8;
    SB_LUT4 i12_3_lut_4_lut (.I0(n7428), .I1(n16485), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n16870));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'he3e0;
    SB_DFF data_in_0___i60 (.Q(\data_in[7] [3]), .C(CLK_c), .D(n10383));   // coms.v(402[9] 410[5])
    SB_LUT4 i3_4_lut (.I0(data_out_7__5__N_543), .I1(n17578), .I2(\data_out[3][6] ), 
            .I3(n17641), .O(n9276));   // coms.v(62[15:196])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i59 (.Q(\data_in[7] [2]), .C(CLK_c), .D(n10382));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i58 (.Q(\data_in[7]_c [1]), .C(CLK_c), .D(n10381));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i57 (.Q(\data_in[7][0] ), .C(CLK_c), .D(n10380));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i56 (.Q(\data_in[6] [7]), .C(CLK_c), .D(n10379));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i55 (.Q(\data_in[6] [6]), .C(CLK_c), .D(n10378));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17488));   // coms.v(228[15:344])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), 
            .E(VCC_net), .D(n10259));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), 
            .E(VCC_net), .D(n10255));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), 
            .E(VCC_net), .D(n10252));   // coms.v(428[12] 532[6])
    SB_LUT4 i3_4_lut_adj_827 (.I0(\data_out[5] [3]), .I1(n9276), .I2(n8634), 
            .I3(n17457), .O(n17623));   // coms.v(116[16:91])
    defparam i3_4_lut_adj_827.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_828 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17473));   // coms.v(224[15:379])
    defparam i1_2_lut_adj_828.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i54 (.Q(\data_in[6] [5]), .C(CLK_c), .D(n10377));   // coms.v(402[9] 410[5])
    SB_LUT4 i15771_4_lut (.I0(data_out_7__1__N_626), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n8926), .I3(n17623), .O(n17916));   // coms.v(277[4] 373[11])
    defparam i15771_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out[6] [7]), 
            .I1(\data_out[7] [7]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), 
            .E(VCC_net), .D(n10311));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_829 (.I0(\data_in_frame[5] [7]), .I1(n8666), .I2(GND_net), 
            .I3(GND_net), .O(n17519));   // coms.v(116[16:91])
    defparam i1_2_lut_adj_829.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(n9204), .I1(n9365), .I2(n8695), .I3(n17430), 
            .O(n22));   // coms.v(517[9:65])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n17605), .I1(n9380), .I2(\data_in_frame[6] [3]), 
            .I3(GND_net), .O(n20));   // coms.v(517[9:65])
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(n9208), .I1(n22), .I2(n16), .I3(\data_in_frame[6] [6]), 
            .O(n24));   // coms.v(517[9:65])
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n17473), .I1(n24), .I2(n20), .I3(n17519), 
            .O(n9355));   // coms.v(517[9:65])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_830 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[3] [3]), .O(n8645));   // coms.v(452[9:67])
    defparam i3_4_lut_adj_830.LUT_INIT = 16'h6996;
    SB_LUT4 i15753_2_lut (.I0(data_out_7__7__N_519), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18017));
    defparam i15753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_687_i1_4_lut (.I0(n17916), .I1(\rand_setpoint[8] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2019[0]));   // coms.v(277[4] 373[11])
    defparam mux_687_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7_4_lut (.I0(n2565), .I1(n2574), .I2(n17412), .I3(n17594), 
            .O(n23));
    defparam i7_4_lut.LUT_INIT = 16'hb7ed;
    SB_LUT4 i1_2_lut_adj_831 (.I0(\data_out[8] [6]), .I1(\data_out[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9087));   // coms.v(169[15:130])
    defparam i1_2_lut_adj_831.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_832 (.I0(\data_in_frame[4] [7]), .I1(n8645), .I2(GND_net), 
            .I3(GND_net), .O(n17513));   // coms.v(74[16:53])
    defparam i1_2_lut_adj_832.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), 
            .E(VCC_net), .D(n10249));   // coms.v(428[12] 532[6])
    SB_LUT4 n18474_bdd_4_lut (.I0(n18474), .I1(\data_out_frame2[13] [1]), 
            .I2(\data_out_frame2[12] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n17836));
    defparam n18474_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR byte_transmit_counter2_2272__i0 (.Q(byte_transmit_counter2[0]), 
            .C(CLK_c), .E(n9605), .D(n37[0]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_LUT4 i1_2_lut_adj_833 (.I0(\data_out[7] [5]), .I1(\data_out[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n8812));   // coms.v(173[15:115])
    defparam i1_2_lut_adj_833.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), 
            .E(VCC_net), .D(n10242));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_4_lut (.I0(n8812), .I1(n9087), .I2(data_out_7__2__N_574), 
            .I3(\data_out[7] [1]), .O(data_out_10__2__N_179));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i7715_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n9519), .I3(\data_out[2] [3]), .O(n10131));
    defparam i7715_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16001 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [1]), .I2(\data_out_frame2[19] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18468));
    defparam byte_transmit_counter2_0__bdd_4_lut_16001.LUT_INIT = 16'he4aa;
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), 
            .E(VCC_net), .D(n10239));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1][1] ), .C(CLK_c), 
            .E(VCC_net), .D(n10236));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_834 (.I0(data_out_6__7__N_678), .I1(data_out_6__1__N_850), 
            .I2(GND_net), .I3(GND_net), .O(n17445));   // coms.v(180[16:109])
    defparam i1_2_lut_adj_834.LUT_INIT = 16'h6666;
    SB_LUT4 n18468_bdd_4_lut (.I0(n18468), .I1(\data_out_frame2[17] [1]), 
            .I2(\data_out_frame2[16] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n18471));
    defparam n18468_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), 
            .E(VCC_net), .D(n10232));   // coms.v(428[12] 532[6])
    SB_LUT4 i9088_3_lut (.I0(\data_in[5] [1]), .I1(\data_in[6]_c [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10365));   // coms.v(377[7:20])
    defparam i9088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_835 (.I0(data_out_6__3__N_788), .I1(\data_out[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n8634));   // coms.v(180[16:109])
    defparam i1_2_lut_adj_835.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[10] [2]), .I1(n8995), .I2(n9355), 
            .I3(\data_in_frame[10] [5]), .O(n10));   // coms.v(229[15:344])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n9131), .I1(n10), .I2(n17418), .I3(GND_net), 
            .O(n17420));   // coms.v(229[15:344])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_836 (.I0(data_out_5__5__N_950), .I1(n8767), .I2(GND_net), 
            .I3(GND_net), .O(n17457));   // coms.v(116[16:91])
    defparam i1_2_lut_adj_836.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), 
            .E(VCC_net), .D(n10308));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), 
            .E(VCC_net), .D(n10229));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_837 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[10][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n8995));   // coms.v(226[15:362])
    defparam i1_2_lut_adj_837.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), 
            .E(VCC_net), .D(n10226));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_4_lut (.I0(n17641), .I1(n17457), .I2(n8964), .I3(n17525), 
            .O(n17415));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_838 (.I0(n9043), .I1(n8886), .I2(GND_net), .I3(GND_net), 
            .O(n17535));   // coms.v(177[16:29])
    defparam i1_2_lut_adj_838.LUT_INIT = 16'h6666;
    SB_DFF byte_transmit_counter__i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
           .D(n16856));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i53 (.Q(\data_in[6]_c [4]), .C(CLK_c), .D(n10376));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i52 (.Q(\data_in[6][3] ), .C(CLK_c), .D(n10375));   // coms.v(402[9] 410[5])
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), 
            .E(VCC_net), .D(n10222));   // coms.v(428[12] 532[6])
    SB_DFFE \data_out_10[[5__3512  (.Q(\data_out[10] [5]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__5__N_132));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i51 (.Q(\data_in[6][2] ), .C(CLK_c), .D(n10374));   // coms.v(402[9] 410[5])
    SB_LUT4 data_out_5__7__I_0_3654_2_lut (.I0(data_out_7__7__N_519), .I1(data_out_7__6__N_530), 
            .I2(GND_net), .I3(GND_net), .O(data_out_7__1__N_626));   // coms.v(114[16:29])
    defparam data_out_5__7__I_0_3654_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_839 (.I0(\data_in_frame[9] [1]), .I1(n17504), .I2(n9240), 
            .I3(n17535), .O(n17537));   // coms.v(236[16:315])
    defparam i3_4_lut_adj_839.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_840 (.I0(\data_out[0][1] ), .I1(\data_out[0][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n8777));
    defparam i1_2_lut_adj_840.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_841 (.I0(n2561), .I1(n8056), .I2(n17544), .I3(n2566), 
            .O(n19_c));
    defparam i3_4_lut_adj_841.LUT_INIT = 16'hde7b;
    SB_LUT4 i7720_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n9519), .I3(data_out_5__5__N_950), .O(n10136));
    defparam i7720_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 byte_transmit_counter2_1__bdd_4_lut (.I0(byte_transmit_counter2[1]), 
            .I1(n17955), .I2(n5_adj_2425), .I3(byte_transmit_counter2[2]), 
            .O(n18456));
    defparam byte_transmit_counter2_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_842 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9148));   // coms.v(225[15:370])
    defparam i1_2_lut_adj_842.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i50 (.Q(\data_in[6]_c [1]), .C(CLK_c), .D(n10373));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i49 (.Q(\data_in[6][0] ), .C(CLK_c), .D(n10372));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i48 (.Q(\data_in[5] [7]), .C(CLK_c), .D(n10371));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i47 (.Q(\data_in[5] [6]), .C(CLK_c), .D(n10370));   // coms.v(402[9] 410[5])
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), 
            .E(VCC_net), .D(n10219));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i46 (.Q(\data_in[5] [5]), .C(CLK_c), .D(n10369));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i45 (.Q(\data_in[5] [4]), .C(CLK_c), .D(n10368));   // coms.v(402[9] 410[5])
    SB_LUT4 i7722_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n9519), .I3(\data_out[0] [6]), .O(n10138));
    defparam i7722_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 i1_2_lut_adj_843 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17482));   // coms.v(235[16:323])
    defparam i1_2_lut_adj_843.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i44 (.Q(\data_in[5] [3]), .C(CLK_c), .D(n10367));   // coms.v(402[9] 410[5])
    SB_DFFE \data_out_10[[4__3513  (.Q(\data_out[10] [4]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__4__N_147));   // coms.v(274[12] 374[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), 
            .E(VCC_net), .D(n10216));   // coms.v(428[12] 532[6])
    SB_DFF tx_active_prev_3508 (.Q(tx_active_prev), .C(CLK_c), .D(tx_active));   // coms.v(274[12] 374[6])
    SB_DFFSR tx_transmit_3509 (.Q(tx_transmit), .C(CLK_c), .D(n17339), 
            .R(n4430));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[7__3534  (.Q(\data_out[7] [7]), .C(CLK_c), .E(n9518), 
            .D(n1774[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[6__3535  (.Q(\data_out[7] [6]), .C(CLK_c), .E(n9518), 
            .D(n1809[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[5__3536  (.Q(\data_out[7] [5]), .C(CLK_c), .E(n9518), 
            .D(n1844[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[4__3537  (.Q(\data_out[7] [4]), .C(CLK_c), .E(n9518), 
            .D(n1879[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[3__3538  (.Q(\data_out[7] [3]), .C(CLK_c), .E(n9518), 
            .D(n1914[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[2__3539  (.Q(\data_out[7] [2]), .C(CLK_c), .E(n9518), 
            .D(n1949[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[1__3540  (.Q(\data_out[7] [1]), .C(CLK_c), .E(n9518), 
            .D(n1984[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_7[[0__3541  (.Q(\data_out[7] [0]), .C(CLK_c), .E(n9518), 
            .D(n2019[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[7__3542  (.Q(\data_out[6] [7]), .C(CLK_c), .E(n9519), 
            .D(n2054[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[6__3543  (.Q(\data_out[6] [6]), .C(CLK_c), .E(n9519), 
            .D(n2089[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[5__3544  (.Q(\data_out[6] [5]), .C(CLK_c), .E(n9519), 
            .D(n2124[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[4__3545  (.Q(\data_out[6] [4]), .C(CLK_c), .E(n9519), 
            .D(n2159[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[3__3546  (.Q(\data_out[6] [3]), .C(CLK_c), .E(n9519), 
            .D(n2194[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[2__3547  (.Q(\data_out[6] [2]), .C(CLK_c), .E(n9519), 
            .D(n2229[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[1__3548  (.Q(\data_out[6] [1]), .C(CLK_c), .E(n9519), 
            .D(n2264[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_6[[0__3549  (.Q(\data_out[6] [0]), .C(CLK_c), .E(n9519), 
            .D(n2299[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[7__3550  (.Q(data_out_7__7__N_519), .C(CLK_c), 
            .E(n9519), .D(n2334[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[6__3551  (.Q(data_out_7__6__N_530), .C(CLK_c), 
            .E(n9519), .D(n2369[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[5__3552  (.Q(data_out_7__5__N_543), .C(CLK_c), 
            .E(n9519), .D(n2404[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[4__3553  (.Q(data_out_7__4__N_556), .C(CLK_c), 
            .E(n9519), .D(n2439[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[3__3554  (.Q(\data_out[5] [3]), .C(CLK_c), .E(n9519), 
            .D(n2474[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[2__3555  (.Q(\data_out[5] [2]), .C(CLK_c), .E(n9519), 
            .D(n2509[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[1__3556  (.Q(\data_out[5] [1]), .C(CLK_c), .E(n9519), 
            .D(n2544[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_5[[0__3557  (.Q(data_out_6__3__N_788), .C(CLK_c), 
            .E(n9519), .D(n2579[0]));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_1[[1__3588  (.Q(\data_out[1] [1]), .C(CLK_c), .E(n9519), 
            .D(n3203[0]));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i1 (.Q(\data_out_frame2[0] [0]), .C(CLK_c), 
           .D(n9685));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), 
            .E(VCC_net), .D(n10213));   // coms.v(428[12] 532[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
            .D(n17214), .S(n1_c));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_844 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_c));   // coms.v(235[16:323])
    defparam i1_2_lut_adj_844.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_845 (.I0(\data_in_frame[9] [0]), .I1(n17585), .I2(n17482), 
            .I3(n6_c), .O(n17587));   // coms.v(235[16:323])
    defparam i4_4_lut_adj_845.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_2426));   // coms.v(383[12:25])
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), 
            .E(VCC_net), .D(n10631));   // coms.v(428[12] 532[6])
    SB_LUT4 i6_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n9631));
    defparam i6_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 add_3777_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n16314), .O(n7260[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), 
            .E(VCC_net), .D(n10210));   // coms.v(428[12] 532[6])
    SB_LUT4 i5_4_lut (.I0(n2568), .I1(n2564), .I2(n9355), .I3(n17538), 
            .O(n21));
    defparam i5_4_lut.LUT_INIT = 16'hde7b;
    SB_LUT4 add_3777_7_lut (.I0(n29), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n16309), .O(n18012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3777_4 (.CI(n16306), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n16307));
    SB_LUT4 i4_4_lut_adj_847 (.I0(n20_adj_2427), .I1(n23_adj_2426), .I2(\data_in_frame[0] [1]), 
            .I3(\data_in_frame[5] [3]), .O(n10_adj_2428));   // coms.v(128[17:38])
    defparam i4_4_lut_adj_847.LUT_INIT = 16'h6996;
    SB_LUT4 i15663_4_lut (.I0(n17611), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n8777), .I3(n17659), .O(n17918));   // coms.v(277[4] 373[11])
    defparam i15663_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(data_out_5__7__N_931), .I1(\data_out[2] [3]), 
            .I2(data_out_6__6__N_729), .I3(\data_out[2][0] ), .O(n17641));   // coms.v(62[15:196])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(data_out_5__7__N_931), .I1(\data_out[2] [3]), 
            .I2(data_out_7__5__N_543), .I3(\data_out[0][3] ), .O(n17499));   // coms.v(62[15:196])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_848 (.I0(n8674), .I1(n10_adj_2428), .I2(\data_in_frame[1] [7]), 
            .I3(GND_net), .O(n9324));   // coms.v(128[17:38])
    defparam i5_3_lut_adj_848.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_1__bdd_4_lut_15987 (.I0(byte_transmit_counter2[1]), 
            .I1(n11), .I2(n12_c), .I3(byte_transmit_counter2[2]), .O(n18444));
    defparam byte_transmit_counter2_1__bdd_4_lut_15987.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[8] [1]), .I3(GND_net), .O(n9144));   // coms.v(229[15:344])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_849 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2429));   // coms.v(178[16:29])
    defparam i1_2_lut_adj_849.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_850 (.I0(n9151), .I1(\data_in_frame[6] [7]), .I2(n9144), 
            .I3(n6_adj_2429), .O(n17588));   // coms.v(178[16:29])
    defparam i4_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_851 (.I0(n17588), .I1(\data_in_frame[10] [5]), 
            .I2(n17433), .I3(GND_net), .O(n17590));   // coms.v(178[16:29])
    defparam i2_3_lut_adj_851.LUT_INIT = 16'h9696;
    SB_DFF \UART_TRANSMITTER.state_i0_i0  (.Q(\UART_TRANSMITTER.state[0] ), 
           .C(CLK_c), .D(n16864));   // coms.v(274[12] 374[6])
    SB_LUT4 i1_2_lut_adj_852 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9240));   // coms.v(236[16:315])
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_CARRY add_3777_12 (.CI(n16314), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n16315));
    SB_DFFE delay_counter_i0_i0 (.Q(\delay_counter[0] ), .C(CLK_c), .E(VCC_net), 
            .D(n10196));   // coms.v(274[12] 374[6])
    SB_LUT4 mux_661_i1_4_lut (.I0(n17918), .I1(\rand_setpoint[9] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1984[0]));   // coms.v(277[4] 373[11])
    defparam mux_661_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2_3_lut_adj_853 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n9043));   // coms.v(177[16:29])
    defparam i2_3_lut_adj_853.LUT_INIT = 16'h9696;
    SB_LUT4 n18444_bdd_4_lut (.I0(n18444), .I1(n9), .I2(n8_c), .I3(byte_transmit_counter2[2]), 
            .O(n18447));
    defparam n18444_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n10188));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), 
            .E(VCC_net), .D(n10305));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_adj_854 (.I0(n17647), .I1(n8890), .I2(n2567), .I3(GND_net), 
            .O(n17648));   // coms.v(167[15:498])
    defparam i2_3_lut_adj_854.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_855 (.I0(\data_out[3][4] ), .I1(\data_out[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n17525));   // coms.v(62[15:196])
    defparam i1_2_lut_adj_855.LUT_INIT = 16'h6666;
    SB_DFFE \data_out_10[[3__3514  (.Q(\data_out[10] [3]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__3__N_163));   // coms.v(274[12] 374[6])
    SB_CARRY add_3777_7 (.CI(n16309), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n16310));
    SB_LUT4 i3_4_lut_adj_856 (.I0(\data_out[2][0] ), .I1(\data_out[0][0] ), 
            .I2(\data_out[0][1] ), .I3(n17525), .O(n17644));   // coms.v(63[15:74])
    defparam i3_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_857 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n9317));   // coms.v(231[15:344])
    defparam i2_3_lut_adj_857.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_858 (.I0(\data_out[5] [2]), .I1(data_out_6__3__N_781), 
            .I2(data_out_7__6__N_530), .I3(n17644), .O(data_out_7__2__N_574));   // coms.v(63[15:74])
    defparam i3_4_lut_adj_858.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i43 (.Q(\data_in[5] [2]), .C(CLK_c), .D(n10366));   // coms.v(402[9] 410[5])
    SB_LUT4 i15760_2_lut (.I0(\rand_setpoint[10] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17921));   // coms.v(277[4] 373[11])
    defparam i15760_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3777_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n16313), .O(n7260[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_635_i1_4_lut (.I0(data_out_7__2__N_574), .I1(n17921), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1949[0]));   // coms.v(277[4] 373[11])
    defparam mux_635_i1_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_adj_859 (.I0(\data_out[0][1] ), .I1(\data_out[1][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n8600));   // coms.v(64[15:74])
    defparam i1_2_lut_adj_859.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_860 (.I0(n2560), .I1(n2572), .I2(n17582), .I3(n17588), 
            .O(n18));
    defparam i2_4_lut_adj_860.LUT_INIT = 16'h7bde;
    SB_LUT4 i4_4_lut_adj_861 (.I0(n9176), .I1(\data_in_frame[0] [6]), .I2(\data_in_frame[0] [5]), 
            .I3(\data_in_frame[4] [4]), .O(n10_adj_2430));   // coms.v(383[12:25])
    defparam i4_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i71 (.Q(\data_in[8] [6]), .C(CLK_c), .D(n10394));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i70 (.Q(\data_in[8] [5]), .C(CLK_c), .D(n10393));   // coms.v(402[9] 410[5])
    SB_LUT4 i12_4_lut_adj_862 (.I0(n23), .I1(n17536), .I2(n2571), .I3(n17547), 
            .O(n28));
    defparam i12_4_lut_adj_862.LUT_INIT = 16'hfbbf;
    SB_LUT4 i2_3_lut_adj_863 (.I0(data_out_6__3__N_781), .I1(\data_out[5] [3]), 
            .I2(n8600), .I3(GND_net), .O(n17635));   // coms.v(174[15:122])
    defparam i2_3_lut_adj_863.LUT_INIT = 16'h9696;
    SB_LUT4 i15674_3_lut (.I0(data_out_7__7__N_519), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n17635), .I3(GND_net), .O(n17922));   // coms.v(277[4] 373[11])
    defparam i15674_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 add_3776_9_lut (.I0(GND_net), .I1(\byte_transmit_counter[7] ), 
            .I2(GND_net), .I3(n16356), .O(tx_transmit_N_2239[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3776_8_lut (.I0(GND_net), .I1(\byte_transmit_counter[6] ), 
            .I2(GND_net), .I3(n16355), .O(tx_transmit_N_2239[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_864 (.I0(n9254), .I1(n19), .I2(n8725), .I3(n9317), 
            .O(n17594));   // coms.v(231[15:344])
    defparam i3_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 add_3777_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n16308), .O(n7260[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i34 (.Q(\data_in[4] [1]), .C(CLK_c), .D(n10148));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_adj_865 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[1][1] ), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n17485));   // coms.v(452[9:67])
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 mux_609_i1_4_lut (.I0(n17922), .I1(\rand_setpoint[11] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1914[0]));   // coms.v(277[4] 373[11])
    defparam mux_609_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_3777_11 (.CI(n16313), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n16314));
    SB_LUT4 i15673_2_lut (.I0(\rand_setpoint[12] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17931));   // coms.v(277[4] 373[11])
    defparam i15673_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3777_10_lut (.I0(n29), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n16312), .O(n18011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3777_3 (.CI(n16305), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n16306));
    SB_LUT4 mux_583_i1_4_lut (.I0(data_out_7__4__N_550), .I1(n17931), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1879[0]));   // coms.v(277[4] 373[11])
    defparam mux_583_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i10_4_lut (.I0(n19_c), .I1(n17592), .I2(n2575), .I3(n8890), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i15690_2_lut (.I0(\rand_setpoint[13] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17925));   // coms.v(277[4] 373[11])
    defparam i15690_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n10144));   // coms.v(402[9] 410[5])
    SB_LUT4 n18372_bdd_4_lut (.I0(n18372), .I1(n6_adj_2432), .I2(n18082), 
            .I3(byte_transmit_counter2[3]), .O(n18375));
    defparam n18372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut (.I0(byte_transmit_counter2[2]), 
            .I1(n17773), .I2(n17779), .I3(byte_transmit_counter2[3]), 
            .O(n18432));
    defparam byte_transmit_counter2_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY add_3776_8 (.CI(n16355), .I0(\byte_transmit_counter[6] ), .I1(GND_net), 
            .CO(n16356));
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), 
            .E(VCC_net), .D(n10622));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), 
            .E(VCC_net), .D(n10619));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i37 (.Q(\data_in[4]_c [4]), .C(CLK_c), .D(n10143));   // coms.v(402[9] 410[5])
    SB_DFF \FRAME_MATCHER.next_state_i1  (.Q(\FRAME_MATCHER.next_state[1] ), 
           .C(CLK_c), .D(n6));   // coms.v(428[12] 532[6])
    SB_CARRY add_3777_10 (.CI(n16312), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n16313));
    SB_LUT4 i11_4_lut_adj_866 (.I0(n21), .I1(n2562), .I2(n17481), .I3(n17541), 
            .O(n27));
    defparam i11_4_lut_adj_866.LUT_INIT = 16'hfbfe;
    SB_DFF \UART_TRANSMITTER.state_i0_i2  (.Q(\UART_TRANSMITTER.state[2] ), 
           .C(CLK_c), .D(n38));   // coms.v(274[12] 374[6])
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), 
            .E(VCC_net), .D(n10614));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), 
            .E(VCC_net), .D(n10611));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), 
           .D(n10608));   // coms.v(428[12] 532[6])
    SB_LUT4 add_3776_7_lut (.I0(GND_net), .I1(\byte_transmit_counter[5] ), 
            .I2(GND_net), .I3(n16354), .O(tx_transmit_N_2239[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), 
           .D(n10350));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), 
           .D(n10356));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i153 (.Q(\data_out_frame2[19][0] ), .C(CLK_c), 
           .D(n10604));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i152 (.Q(\data_out_frame2[18] [7]), .C(CLK_c), 
           .D(n10603));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i151 (.Q(\data_out_frame2[18] [6]), .C(CLK_c), 
           .D(n10602));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i150 (.Q(\data_out_frame2[18] [5]), .C(CLK_c), 
           .D(n10601));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i149 (.Q(\data_out_frame2[18] [4]), .C(CLK_c), 
           .D(n10600));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i148 (.Q(\data_out_frame2[18] [3]), .C(CLK_c), 
           .D(n10599));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i147 (.Q(\data_out_frame2[18] [2]), .C(CLK_c), 
           .D(n10598));   // coms.v(428[12] 532[6])
    SB_LUT4 i9_4_lut_adj_867 (.I0(n2570), .I1(n18), .I2(n17648), .I3(n17585), 
            .O(n25));
    defparam i9_4_lut_adj_867.LUT_INIT = 16'hdfef;
    SB_DFF byte_transmit_counter__i6 (.Q(\byte_transmit_counter[6] ), .C(CLK_c), 
           .D(n8));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i7 (.Q(\byte_transmit_counter[7] ), .C(CLK_c), 
           .D(n8_adj_3));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i146 (.Q(\data_out_frame2[18] [1]), .C(CLK_c), 
           .D(n10597));   // coms.v(428[12] 532[6])
    SB_LUT4 n18432_bdd_4_lut (.I0(n18432), .I1(n6_adj_2436), .I2(n18074), 
            .I3(byte_transmit_counter2[3]), .O(n18435));
    defparam n18432_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_557_i1_4_lut (.I0(n17499), .I1(n17925), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1844[0]));   // coms.v(277[4] 373[11])
    defparam mux_557_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_3_lut (.I0(\data_out_frame2[0] [4]), .I1(n14631), .I2(n142), 
            .I3(GND_net), .O(n9671));   // coms.v(422[11:16])
    defparam i1_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i2_3_lut_adj_868 (.I0(data_out_7__6__N_530), .I1(data_out_6__6__N_729), 
            .I2(\data_out[0][5] ), .I3(GND_net), .O(n17465));   // coms.v(173[15:115])
    defparam i2_3_lut_adj_868.LUT_INIT = 16'h9696;
    SB_LUT4 i15763_2_lut (.I0(\rand_setpoint[14] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17906));   // coms.v(277[4] 373[11])
    defparam i15763_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_531_i1_4_lut (.I0(n17465), .I1(n17906), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1809[0]));   // coms.v(277[4] 373[11])
    defparam mux_531_i1_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_3_lut_adj_869 (.I0(\data_out_frame2[0] [3]), .I1(n14631), 
            .I2(n142), .I3(GND_net), .O(n9674));   // coms.v(422[11:16])
    defparam i1_3_lut_adj_869.LUT_INIT = 16'hcece;
    SB_LUT4 select_220_Select_1_i1_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [2]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.next_state[1] ), .O(n1_adj_2437));
    defparam select_220_Select_1_i1_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), 
            .E(VCC_net), .D(n10649));   // coms.v(428[12] 532[6])
    SB_LUT4 n18456_bdd_4_lut_4_lut (.I0(byte_transmit_counter2[0]), .I1(\data_out_frame2[0] [4]), 
            .I2(byte_transmit_counter2[2]), .I3(n18456), .O(n18459));
    defparam n18456_bdd_4_lut_4_lut.LUT_INIT = 16'hfa04;
    SB_LUT4 i1_4_lut_adj_870 (.I0(\FRAME_MATCHER.state [2]), .I1(n31), .I2(n5_adj_2438), 
            .I3(\FRAME_MATCHER.state [1]), .O(n136));
    defparam i1_4_lut_adj_870.LUT_INIT = 16'hfaee;
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), 
            .E(VCC_net), .D(n10652));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_4_lut_adj_871 (.I0(data_out_5__7__N_931), .I1(\data_out[3][6] ), 
            .I2(data_out_7__4__N_556), .I3(n17400), .O(data_out_7__4__N_550));   // coms.v(169[15:130])
    defparam i2_3_lut_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), 
            .E(VCC_net), .D(n10655));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), 
            .E(VCC_net), .D(n10659));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), 
            .E(VCC_net), .D(n10662));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), 
           .D(n10663));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), 
           .D(n10314));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), 
           .D(n10262));   // coms.v(428[12] 532[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), 
            .E(VCC_net), .D(n10671));   // coms.v(428[12] 532[6])
    SB_DFF delay_counter_i0_i14 (.Q(\delay_counter[14] ), .C(CLK_c), .D(n10674));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i13 (.Q(\delay_counter[13] ), .C(CLK_c), .D(n10675));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .D(n10676));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .D(n10071));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .D(n10068));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .D(n10065));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .D(n10680));   // coms.v(274[12] 374[6])
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), 
            .E(VCC_net), .D(n10683));   // coms.v(428[12] 532[6])
    SB_DFF delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .D(n10059));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .D(n10056));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .D(n10686));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .D(n10050));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .D(n10047));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .D(n10042));   // coms.v(274[12] 374[6])
    SB_DFF delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .D(n10037));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n10691));   // coms.v(402[9] 410[5])
    SB_DFF \UART_TRANSMITTER.state_i0_i1  (.Q(\UART_TRANSMITTER.state[1] ), 
           .C(CLK_c), .D(n16870));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
           .D(n16858));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i2 (.Q(\byte_transmit_counter[2] ), .C(CLK_c), 
           .D(n8_adj_4));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i3 (.Q(\byte_transmit_counter[3] ), .C(CLK_c), 
           .D(n8_adj_5));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i4 (.Q(\byte_transmit_counter[4] ), .C(CLK_c), 
           .D(n8_adj_6));   // coms.v(274[12] 374[6])
    SB_DFF byte_transmit_counter__i5 (.Q(\byte_transmit_counter[5] ), .C(CLK_c), 
           .D(n8_adj_7));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i39 (.Q(\data_in[4]_c [6]), .C(CLK_c), .D(n10302));   // coms.v(402[9] 410[5])
    SB_LUT4 i12304_4_lut (.I0(n1_adj_2443), .I1(n136), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n157), .O(n14631));   // coms.v(422[11:16])
    defparam i12304_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i15683_3_lut (.I0(data_out_7__7__N_519), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(data_out_6__7__N_675), .I3(GND_net), .O(n17928));   // coms.v(277[4] 373[11])
    defparam i15683_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i1_3_lut_adj_872 (.I0(\data_out_frame2[0] [2]), .I1(n14631), 
            .I2(n142), .I3(GND_net), .O(n9677));   // coms.v(422[11:16])
    defparam i1_3_lut_adj_872.LUT_INIT = 16'hcece;
    SB_LUT4 mux_505_i1_4_lut (.I0(n17928), .I1(\rand_setpoint[15] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1774[0]));   // coms.v(277[4] 373[11])
    defparam mux_505_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_3_lut (.I0(data_out_5__7__N_931), .I1(\data_out[3][6] ), 
            .I2(\data_out[3][5] ), .I3(GND_net), .O(data_out_6__3__N_781));   // coms.v(169[15:130])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out[6] [6]), 
            .I1(\data_out[7] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2444));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_873 (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n97), .I3(GND_net), .O(n16_adj_2445));   // coms.v(277[4] 373[11])
    defparam i1_3_lut_adj_873.LUT_INIT = 16'haeae;
    SB_DFF data_out_frame2_0___i145 (.Q(\data_out_frame2[18] [0]), .C(CLK_c), 
           .D(n10596));   // coms.v(428[12] 532[6])
    SB_LUT4 i15698_2_lut (.I0(data_out_7__6__N_530), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17949));
    defparam i15698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_874 (.I0(n149), .I1(tx_transmit_N_2239[3]), .I2(n2649[0]), 
            .I3(n16_adj_2445), .O(n19_adj_2446));   // coms.v(277[4] 373[11])
    defparam i1_4_lut_adj_874.LUT_INIT = 16'h7350;
    SB_DFF data_out_frame2_0___i144 (.Q(\data_out_frame2[17] [7]), .C(CLK_c), 
           .D(n10595));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_4_lut_adj_875 (.I0(\UART_TRANSMITTER.state[0] ), .I1(n13415), 
            .I2(n19_adj_2446), .I3(n8550), .O(n17339));   // coms.v(277[4] 373[11])
    defparam i1_4_lut_adj_875.LUT_INIT = 16'h0010;
    SB_DFF data_out_frame2_0___i143 (.Q(\data_out_frame2[17] [6]), .C(CLK_c), 
           .D(n10594));   // coms.v(428[12] 532[6])
    SB_LUT4 add_3777_2_lut (.I0(GND_net), .I1(\delay_counter[0] ), .I2(GND_net), 
            .I3(VCC_net), .O(n7260[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_876 (.I0(n17556), .I1(data_out_6__7__N_675), .I2(n17492), 
            .I3(GND_net), .O(data_out_10__7__N_101));   // coms.v(174[15:122])
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i69 (.Q(\data_in[8] [4]), .C(CLK_c), .D(n10392));   // coms.v(402[9] 410[5])
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n5_adj_2438));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_0___i68 (.Q(\data_in[8] [3]), .C(CLK_c), .D(n10391));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15945 (.I0(byte_transmit_counter[1]), 
            .I1(n17941), .I2(n5_adj_2447), .I3(\byte_transmit_counter[2] ), 
            .O(n18396));
    defparam byte_transmit_counter_1__bdd_4_lut_15945.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_877 (.I0(n17445), .I1(n17620), .I2(n17510), .I3(n17638), 
            .O(data_out_9__1__N_462));   // coms.v(180[16:109])
    defparam i3_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_878 (.I0(\data_out[6] [0]), .I1(\data_out[7] [7]), 
            .I2(\data_out[7] [6]), .I3(GND_net), .O(n8950));   // coms.v(171[15:115])
    defparam i2_3_lut_adj_878.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out[6] [4]), 
            .I1(\data_out[7] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2447));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i115 (.Q(\data_in[14] [2]), .C(CLK_c), .D(n10438));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i114 (.Q(\data_in[14] [1]), .C(CLK_c), .D(n10437));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i113 (.Q(\data_in[14] [0]), .C(CLK_c), .D(n10436));   // coms.v(402[9] 410[5])
    SB_LUT4 i15689_2_lut (.I0(data_out_7__4__N_556), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17941));
    defparam i15689_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i112 (.Q(\data_in[13] [7]), .C(CLK_c), .D(n10435));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i111 (.Q(\data_in[13] [6]), .C(CLK_c), .D(n10434));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i110 (.Q(\data_in[13] [5]), .C(CLK_c), .D(n10433));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i142 (.Q(\data_out_frame2[17] [5]), .C(CLK_c), 
           .D(n10593));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i141 (.Q(\data_out_frame2[17] [4]), .C(CLK_c), 
           .D(n10592));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i140 (.Q(\data_out_frame2[17] [3]), .C(CLK_c), 
           .D(n10591));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_adj_879 (.I0(data_out_6__2__N_804), .I1(n8922), .I2(\data_out[1] [1]), 
            .I3(GND_net), .O(data_out_9__2__N_446));   // coms.v(181[16:29])
    defparam i2_3_lut_adj_879.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_880 (.I0(\data_out[7] [2]), .I1(\data_out[7] [3]), 
            .I2(data_out_7__4__N_550), .I3(n8950), .O(data_out_10__4__N_147));   // coms.v(171[15:115])
    defparam i3_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i13621_3_lut (.I0(\data_in[8] [4]), .I1(\data_in[9] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10392));   // coms.v(377[7:20])
    defparam i13621_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame2_0___i139 (.Q(\data_out_frame2[17] [2]), .C(CLK_c), 
           .D(n10590));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i138 (.Q(\data_out_frame2[17] [1]), .C(CLK_c), 
           .D(n10589));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i137 (.Q(\data_out_frame2[17] [0]), .C(CLK_c), 
           .D(n10588));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i136 (.Q(\data_out_frame2[16] [7]), .C(CLK_c), 
           .D(n10587));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i135 (.Q(\data_out_frame2[16] [6]), .C(CLK_c), 
           .D(n10586));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i134 (.Q(\data_out_frame2[16] [5]), .C(CLK_c), 
           .D(n10585));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i133 (.Q(\data_out_frame2[16] [4]), .C(CLK_c), 
           .D(n10584));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i132 (.Q(\data_out_frame2[16] [3]), .C(CLK_c), 
           .D(n10583));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i131 (.Q(\data_out_frame2[16] [2]), .C(CLK_c), 
           .D(n10582));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i130 (.Q(\data_out_frame2[16] [1]), .C(CLK_c), 
           .D(n10581));   // coms.v(428[12] 532[6])
    SB_LUT4 i15794_2_lut (.I0(\data_out[0][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18094));
    defparam i15794_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame2_0___i129 (.Q(\data_out_frame2[16] [0]), .C(CLK_c), 
           .D(n10580));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i128 (.Q(\data_out_frame2[15] [7]), .C(CLK_c), 
           .D(n10579));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i127 (.Q(\data_out_frame2[15] [6]), .C(CLK_c), 
           .D(n10578));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i126 (.Q(\data_out_frame2[15] [5]), .C(CLK_c), 
           .D(n10577));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i125 (.Q(\data_out_frame2[15] [4]), .C(CLK_c), 
           .D(n10576));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i124 (.Q(\data_out_frame2[15] [3]), .C(CLK_c), 
           .D(n10575));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i123 (.Q(\data_out_frame2[15] [2]), .C(CLK_c), 
           .D(n10574));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i67 (.Q(\data_in[8] [2]), .C(CLK_c), .D(n10390));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i109 (.Q(\data_in[13] [4]), .C(CLK_c), .D(n10432));   // coms.v(402[9] 410[5])
    SB_LUT4 i13631_3_lut (.I0(\data_in[5] [4]), .I1(\data_in[6]_c [4]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10368));   // coms.v(377[7:20])
    defparam i13631_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i108 (.Q(\data_in[13] [3]), .C(CLK_c), .D(n10431));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i107 (.Q(\data_in[13] [2]), .C(CLK_c), .D(n10430));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i122 (.Q(\data_out_frame2[15] [1]), .C(CLK_c), 
           .D(n10573));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i121 (.Q(\data_out_frame2[15] [0]), .C(CLK_c), 
           .D(n10572));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i120 (.Q(\data_out_frame2[14] [7]), .C(CLK_c), 
           .D(n10571));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i66 (.Q(\data_in[8] [1]), .C(CLK_c), .D(n10389));   // coms.v(402[9] 410[5])
    SB_LUT4 i15744_2_lut (.I0(\data_out[2] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18095));
    defparam i15744_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i106 (.Q(\data_in[13] [1]), .C(CLK_c), .D(n10429));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i105 (.Q(\data_in[13] [0]), .C(CLK_c), .D(n10428));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i104 (.Q(\data_in[12] [7]), .C(CLK_c), .D(n10427));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i103 (.Q(\data_in[12] [6]), .C(CLK_c), .D(n10426));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i102 (.Q(\data_in[12] [5]), .C(CLK_c), .D(n10425));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i101 (.Q(\data_in[12] [4]), .C(CLK_c), .D(n10424));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i119 (.Q(\data_out_frame2[14] [6]), .C(CLK_c), 
           .D(n10570));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i118 (.Q(\data_out_frame2[14] [5]), .C(CLK_c), 
           .D(n10569));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i117 (.Q(\data_out_frame2[14] [4]), .C(CLK_c), 
           .D(n10568));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i116 (.Q(\data_out_frame2[14] [3]), .C(CLK_c), 
           .D(n10567));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i115 (.Q(\data_out_frame2[14] [2]), .C(CLK_c), 
           .D(n10566));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i114 (.Q(\data_out_frame2[14] [1]), .C(CLK_c), 
           .D(n10565));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i113 (.Q(\data_out_frame2[14] [0]), .C(CLK_c), 
           .D(n10564));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i100 (.Q(\data_in[12] [3]), .C(CLK_c), .D(n10423));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i112 (.Q(\data_out_frame2[13] [7]), .C(CLK_c), 
           .D(n10563));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i111 (.Q(\data_out_frame2[13] [6]), .C(CLK_c), 
           .D(n10562));   // coms.v(428[12] 532[6])
    SB_CARRY add_3776_7 (.CI(n16354), .I0(\byte_transmit_counter[5] ), .I1(GND_net), 
            .CO(n16355));
    SB_LUT4 i2_3_lut_adj_881 (.I0(\data_out[8] [1]), .I1(\data_out[8] [2]), 
            .I2(\data_out[6] [3]), .I3(GND_net), .O(n17556));   // coms.v(174[15:122])
    defparam i2_3_lut_adj_881.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_882 (.I0(\data_out[2][0] ), .I1(data_out_6__6__N_729), 
            .I2(\data_out[0][3] ), .I3(GND_net), .O(n17400));   // coms.v(62[15:196])
    defparam i1_2_lut_3_lut_adj_882.LUT_INIT = 16'h9696;
    SB_LUT4 add_3776_6_lut (.I0(GND_net), .I1(\byte_transmit_counter[4] ), 
            .I2(GND_net), .I3(n16353), .O(tx_transmit_N_2239[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_6 (.CI(n16353), .I0(\byte_transmit_counter[4] ), .I1(GND_net), 
            .CO(n16354));
    SB_DFF data_out_frame2_0___i110 (.Q(\data_out_frame2[13] [5]), .C(CLK_c), 
           .D(n10561));   // coms.v(428[12] 532[6])
    SB_LUT4 add_3776_5_lut (.I0(GND_net), .I1(\byte_transmit_counter[3] ), 
            .I2(GND_net), .I3(n16352), .O(tx_transmit_N_2239[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3777_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n16311), .O(n7260[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_883 (.I0(\data_out[8] [6]), .I1(n17556), .I2(\data_out[6] [7]), 
            .I3(n6_adj_2448), .O(data_out_9__3__N_430));   // coms.v(174[15:122])
    defparam i4_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_884 (.I0(n9306), .I1(\data_in_frame[5] [2]), .I2(n8867), 
            .I3(n17406), .O(n12_adj_2449));   // coms.v(128[17:38])
    defparam i5_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_CARRY add_3776_5 (.CI(n16352), .I0(\byte_transmit_counter[3] ), .I1(GND_net), 
            .CO(n16353));
    SB_DFF data_out_frame2_0___i109 (.Q(\data_out_frame2[13] [4]), .C(CLK_c), 
           .D(n10560));   // coms.v(428[12] 532[6])
    SB_DFF \data_out_0[[0__3597  (.Q(\data_out[0][0] ), .C(CLK_c), .D(n10142));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_0[[1__3596  (.Q(\data_out[0][1] ), .C(CLK_c), .D(n10141));   // coms.v(274[12] 374[6])
    SB_LUT4 i4_4_lut_adj_885 (.I0(n8687), .I1(\data_in_frame[2] [6]), .I2(n2590), 
            .I3(\data_in_frame[5] [2]), .O(n10_adj_2450));   // coms.v(517[9:65])
    defparam i4_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i99 (.Q(\data_in[12] [2]), .C(CLK_c), .D(n10422));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_adj_886 (.I0(\data_in_frame[5] [7]), .I1(n8695), .I2(GND_net), 
            .I3(GND_net), .O(n8064));   // coms.v(120[16:83])
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_887 (.I0(n17470), .I1(n10_adj_2450), .I2(n17532), 
            .I3(GND_net), .O(n17534));   // coms.v(517[9:65])
    defparam i5_3_lut_adj_887.LUT_INIT = 16'h9696;
    SB_LUT4 i9089_3_lut (.I0(\data_in[6]_c [1]), .I1(\data_in[7]_c [1]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10373));   // coms.v(377[7:20])
    defparam i9089_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i98 (.Q(\data_in[12] [1]), .C(CLK_c), .D(n10421));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i108 (.Q(\data_out_frame2[13] [3]), .C(CLK_c), 
           .D(n10559));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i42 (.Q(\data_in[5] [1]), .C(CLK_c), .D(n10365));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame2[6] [4]), 
            .I1(\data_out_frame2[7] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2425));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15709_2_lut (.I0(\data_out_frame2[5] [4]), .I1(byte_transmit_counter2[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17955));
    defparam i15709_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_888 (.I0(\data_out[8] [0]), .I1(\data_out[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17638));   // coms.v(172[15:100])
    defparam i1_2_lut_adj_888.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_889 (.I0(\UART_TRANSMITTER.state[1] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2614[0]));   // coms.v(274[12] 374[6])
    defparam i1_2_lut_adj_889.LUT_INIT = 16'h8888;
    SB_LUT4 i15_2_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n9365));   // coms.v(383[12:25])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \data_out_10[[2__3515  (.Q(\data_out[10] [2]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__2__N_179));   // coms.v(274[12] 374[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_16021 (.I0(byte_transmit_counter[1]), 
            .I1(n18017), .I2(n5), .I3(\byte_transmit_counter[2] ), .O(n18426));
    defparam byte_transmit_counter_1__bdd_4_lut_16021.LUT_INIT = 16'he4aa;
    SB_DFF \data_out_0[[3__3594  (.Q(\data_out[0][3] ), .C(CLK_c), .D(n10140));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i41 (.Q(\data_in[5] [0]), .C(CLK_c), .D(n10364));   // coms.v(402[9] 410[5])
    SB_LUT4 i10642_3_lut (.I0(\data_in[4]_c [6]), .I1(\data_in[5] [6]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10302));   // coms.v(377[7:20])
    defparam i10642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_890 (.I0(\data_out[7] [3]), .I1(\data_out[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2451));   // coms.v(172[15:100])
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_891 (.I0(\data_out[6] [1]), .I1(n17638), .I2(n17499), 
            .I3(n6_adj_2451), .O(data_out_10__5__N_132));   // coms.v(172[15:100])
    defparam i4_4_lut_adj_891.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_892 (.I0(\data_out[0][5] ), .I1(\data_out[0] [6]), 
            .I2(\data_out[1] [1]), .I3(\data_out[1][2] ), .O(n8767));
    defparam i1_2_lut_3_lut_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_893 (.I0(n8062), .I1(n2599), .I2(n2587), .I3(n8751), 
            .O(n20_adj_2452));
    defparam i4_4_lut_adj_893.LUT_INIT = 16'hb7ed;
    SB_LUT4 i8_4_lut (.I0(n11_adj_2453), .I1(n2598), .I2(n12_adj_2449), 
            .I3(n17522), .O(n24_adj_2454));
    defparam i8_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 n18426_bdd_4_lut (.I0(n18426), .I1(n2), .I2(n18089), .I3(\byte_transmit_counter[2] ), 
            .O(n18429));
    defparam n18426_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_in_frame[1] [2]), .I1(n9306), .I2(GND_net), 
            .I3(GND_net), .O(n17424));   // coms.v(71[16:29])
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_CARRY add_3777_6 (.CI(n16308), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n16309));
    SB_DFF data_out_frame2_0___i107 (.Q(\data_out_frame2[13] [2]), .C(CLK_c), 
           .D(n10558));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i106 (.Q(\data_out_frame2[13] [1]), .C(CLK_c), 
           .D(n10557));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i105 (.Q(\data_out_frame2[13] [0]), .C(CLK_c), 
           .D(n10556));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i104 (.Q(\data_out_frame2[12] [7]), .C(CLK_c), 
           .D(n10555));   // coms.v(428[12] 532[6])
    SB_DFFSS tx2_transmit_3602 (.Q(r_SM_Main_2__N_2326[0]), .C(CLK_c), .D(n1_adj_2455), 
            .S(n142));   // coms.v(428[12] 532[6])
    SB_DFFE \data_out_10[[1__3516  (.Q(\data_out[10] [1]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__1__N_196));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_0[[5__3592  (.Q(\data_out[0][5] ), .C(CLK_c), .D(n10139));   // coms.v(274[12] 374[6])
    SB_LUT4 i2_3_lut_4_lut_adj_895 (.I0(\data_out[0][5] ), .I1(\data_out[0] [6]), 
            .I2(data_out_6__7__N_678), .I3(\data_out[2] [3]), .O(data_out_6__7__N_675));
    defparam i2_3_lut_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_DFF \data_out_0[[6__3591  (.Q(\data_out[0] [6]), .C(CLK_c), .D(n10138));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i103 (.Q(\data_out_frame2[12] [6]), .C(CLK_c), 
           .D(n10554));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_896 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9039));   // coms.v(76[16:93])
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i102 (.Q(\data_out_frame2[12] [5]), .C(CLK_c), 
           .D(n10553));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i101 (.Q(\data_out_frame2[12] [4]), .C(CLK_c), 
           .D(n10552));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i100 (.Q(\data_out_frame2[12] [3]), .C(CLK_c), 
           .D(n10551));   // coms.v(428[12] 532[6])
    SB_LUT4 add_3776_4_lut (.I0(GND_net), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n16351), .O(tx_transmit_N_2239[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13627_3_lut (.I0(\data_in[6]_c [4]), .I1(\data_in[7]_c [4]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10376));   // coms.v(377[7:20])
    defparam i13627_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame2_0___i99 (.Q(\data_out_frame2[12] [2]), .C(CLK_c), 
           .D(n10550));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i98 (.Q(\data_out_frame2[12] [1]), .C(CLK_c), 
           .D(n10549));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i97 (.Q(\data_out_frame2[12] [0]), .C(CLK_c), 
           .D(n10548));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i97 (.Q(\data_in[12] [0]), .C(CLK_c), .D(n10420));   // coms.v(402[9] 410[5])
    SB_LUT4 i12_4_lut_adj_897 (.I0(byte_transmit_counter[1]), .I1(tx_transmit_N_2239_c[1]), 
            .I2(n9631), .I3(n17349), .O(n16858));   // coms.v(19[11:32])
    defparam i12_4_lut_adj_897.LUT_INIT = 16'h0aca;
    SB_DFFE \data_out_10[[0__3517  (.Q(\data_out[10] [0]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__0__N_259));   // coms.v(274[12] 374[6])
    SB_LUT4 i4_3_lut_4_lut (.I0(n2839), .I1(n8874), .I2(n8_adj_2459), 
            .I3(n2604), .O(n11_adj_2460));   // coms.v(517[9:65])
    defparam i4_3_lut_4_lut.LUT_INIT = 16'hf9f6;
    SB_DFF \data_out_1[[2__3587  (.Q(\data_out[1][2] ), .C(CLK_c), .D(n10137));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_1[[4__3585  (.Q(data_out_5__5__N_950), .C(CLK_c), .D(n10136));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i40 (.Q(\data_in[4][7] ), .C(CLK_c), .D(n10363));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i62 (.Q(\data_in[7][5] ), .C(CLK_c), .D(n10385));   // coms.v(402[9] 410[5])
    SB_LUT4 i6_4_lut (.I0(n2593), .I1(n2597), .I2(n8886), .I3(n17529), 
            .O(n22_adj_2461));
    defparam i6_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF \data_out_1[[6__3583  (.Q(\data_out[1][6] ), .C(CLK_c), .D(n10135));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_1[[7__3582  (.Q(\data_out[1][7] ), .C(CLK_c), .D(n10134));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_2[[0__3581  (.Q(\data_out[2][0] ), .C(CLK_c), .D(n10133));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_2[[2__3579  (.Q(data_out_6__6__N_729), .C(CLK_c), .D(n10132));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_2[[3__3578  (.Q(\data_out[2] [3]), .C(CLK_c), .D(n10131));   // coms.v(274[12] 374[6])
    SB_LUT4 i2_3_lut_adj_898 (.I0(n8658), .I1(n9039), .I2(\data_in_frame[3] [5]), 
            .I3(GND_net), .O(n17575));   // coms.v(452[9:67])
    defparam i2_3_lut_adj_898.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_899 (.I0(n2595), .I1(n2589), .I2(n9054), .I3(n9103), 
            .O(n23_adj_2462));
    defparam i7_4_lut_adj_899.LUT_INIT = 16'h7bde;
    SB_DFF \data_out_2[[5__3576  (.Q(data_out_6__7__N_678), .C(CLK_c), .D(n10130));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_2[[7__3574  (.Q(data_out_6__1__N_850), .C(CLK_c), .D(n10129));   // coms.v(274[12] 374[6])
    SB_LUT4 i11030_2_lut (.I0(tx_active), .I1(tx_transmit), .I2(GND_net), 
            .I3(GND_net), .O(n13415));
    defparam i11030_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15824_3_lut (.I0(\data_out_frame2[0] [2]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n18084));
    defparam i15824_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15970 (.I0(byte_transmit_counter2[2]), 
            .I1(n17785), .I2(n17788), .I3(byte_transmit_counter2[3]), 
            .O(n18420));
    defparam byte_transmit_counter2_2__bdd_4_lut_15970.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame2[6] [2]), 
            .I1(\data_out_frame2[7] [2]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2463));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18420_bdd_4_lut (.I0(n18420), .I1(n6_adj_2464), .I2(n18076), 
            .I3(byte_transmit_counter2[3]), .O(n18423));
    defparam n18420_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i96 (.Q(\data_out_frame2[11] [7]), .C(CLK_c), 
           .D(n10547));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17430));   // coms.v(452[9:67])
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i96 (.Q(\data_in[11] [7]), .C(CLK_c), .D(n10419));   // coms.v(402[9] 410[5])
    SB_DFF \data_out_3[[0__3573  (.Q(data_out_6__2__N_804), .C(CLK_c), .D(n10128));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i95 (.Q(\data_out_frame2[11] [6]), .C(CLK_c), 
           .D(n10546));   // coms.v(428[12] 532[6])
    SB_LUT4 i5_4_lut_adj_901 (.I0(n8064), .I1(n2596), .I2(n2584), .I3(n9151), 
            .O(n21_adj_2465));
    defparam i5_4_lut_adj_901.LUT_INIT = 16'hb7ed;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame2[5] [2]), 
            .I1(n5_adj_2463), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2466));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_in_0___i95 (.Q(\data_in[11] [6]), .C(CLK_c), .D(n10418));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i94 (.Q(\data_out_frame2[11] [5]), .C(CLK_c), 
           .D(n10545));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i94 (.Q(\data_in[11] [5]), .C(CLK_c), .D(n10417));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i93 (.Q(\data_out_frame2[11] [4]), .C(CLK_c), 
           .D(n10544));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i93 (.Q(\data_in[11] [4]), .C(CLK_c), .D(n10416));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i92 (.Q(\data_out_frame2[11] [3]), .C(CLK_c), 
           .D(n10543));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i92 (.Q(\data_in[11] [3]), .C(CLK_c), .D(n10415));   // coms.v(402[9] 410[5])
    SB_DFF \data_out_3[[2__3571  (.Q(data_out_5__4__N_959), .C(CLK_c), .D(n10127));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i91 (.Q(\data_out_frame2[11] [2]), .C(CLK_c), 
           .D(n10542));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i91 (.Q(\data_in[11] [2]), .C(CLK_c), .D(n10414));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i90 (.Q(\data_out_frame2[11] [1]), .C(CLK_c), 
           .D(n10541));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i90 (.Q(\data_in[11] [1]), .C(CLK_c), .D(n10413));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i89 (.Q(\data_out_frame2[11] [0]), .C(CLK_c), 
           .D(n10540));   // coms.v(428[12] 532[6])
    SB_LUT4 i13628_3_lut (.I0(\data_in[3] [4]), .I1(\data_in[4]_c [4]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10103));   // coms.v(377[7:20])
    defparam i13628_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i89 (.Q(\data_in[11] [0]), .C(CLK_c), .D(n10412));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i88 (.Q(\data_out_frame2[10] [7]), .C(CLK_c), 
           .D(n10539));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i88 (.Q(\data_in[10] [7]), .C(CLK_c), .D(n10411));   // coms.v(402[9] 410[5])
    SB_DFF \data_out_3[[4__3569  (.Q(\data_out[3][4] ), .C(CLK_c), .D(n10126));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i87 (.Q(\data_out_frame2[10] [6]), .C(CLK_c), 
           .D(n10538));   // coms.v(428[12] 532[6])
    SB_LUT4 i241_2_lut (.I0(tx_active), .I1(tx_active_prev), .I2(GND_net), 
            .I3(GND_net), .O(n251));   // coms.v(293[9:37])
    defparam i241_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_out_frame2_0___i86 (.Q(\data_out_frame2[10] [5]), .C(CLK_c), 
           .D(n10537));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i87 (.Q(\data_in[10] [6]), .C(CLK_c), .D(n10410));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i85 (.Q(\data_out_frame2[10] [4]), .C(CLK_c), 
           .D(n10536));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i86 (.Q(\data_in[10] [5]), .C(CLK_c), .D(n10409));   // coms.v(402[9] 410[5])
    SB_DFFE \data_out_9[[7__3518  (.Q(\data_out[9] [7]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__7__N_323));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i84 (.Q(\data_out_frame2[10] [3]), .C(CLK_c), 
           .D(n10535));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i85 (.Q(\data_in[10] [4]), .C(CLK_c), .D(n10408));   // coms.v(402[9] 410[5])
    SB_DFF \data_out_3[[5__3568  (.Q(\data_out[3][5] ), .C(CLK_c), .D(n10125));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i83 (.Q(\data_out_frame2[10] [2]), .C(CLK_c), 
           .D(n10534));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i82 (.Q(\data_out_frame2[10] [1]), .C(CLK_c), 
           .D(n10533));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i84 (.Q(\data_in[10] [3]), .C(CLK_c), .D(n10407));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i81 (.Q(\data_out_frame2[10] [0]), .C(CLK_c), 
           .D(n10532));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i83 (.Q(\data_in[10] [2]), .C(CLK_c), .D(n10406));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i80 (.Q(\data_out_frame2[9] [7]), .C(CLK_c), 
           .D(n10531));   // coms.v(428[12] 532[6])
    SB_LUT4 n18396_bdd_4_lut (.I0(n18396), .I1(n18093), .I2(n18092), .I3(\byte_transmit_counter[2] ), 
            .O(n18399));
    defparam n18396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i79 (.Q(\data_out_frame2[9] [6]), .C(CLK_c), 
           .D(n10530));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i82 (.Q(\data_in[10] [1]), .C(CLK_c), .D(n10405));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i78 (.Q(\data_out_frame2[9] [5]), .C(CLK_c), 
           .D(n10529));   // coms.v(428[12] 532[6])
    SB_LUT4 i3_4_lut_adj_902 (.I0(n2591), .I1(n9324), .I2(n8751), .I3(n17532), 
            .O(n17533));   // coms.v(517[9:65])
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i77 (.Q(\data_out_frame2[9] [4]), .C(CLK_c), 
           .D(n10528));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i76 (.Q(\data_out_frame2[9] [3]), .C(CLK_c), 
           .D(n10527));   // coms.v(428[12] 532[6])
    SB_DFF \data_out_3[[6__3567  (.Q(\data_out[3][6] ), .C(CLK_c), .D(n10124));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i75 (.Q(\data_out_frame2[9] [2]), .C(CLK_c), 
           .D(n10526));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i74 (.Q(\data_out_frame2[9] [1]), .C(CLK_c), 
           .D(n10525));   // coms.v(428[12] 532[6])
    SB_DFF \data_out_3[[7__3566  (.Q(data_out_5__7__N_931), .C(CLK_c), .D(n10123));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0]_c [0]), .C(CLK_c), .D(n10122));   // coms.v(402[9] 410[5])
    SB_LUT4 i13953_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[4][0] ), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10107));   // coms.v(377[7:20])
    defparam i13953_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3776_4 (.CI(n16351), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n16352));
    SB_DFF data_out_frame2_0___i73 (.Q(\data_out_frame2[9] [0]), .C(CLK_c), 
           .D(n10524));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_adj_903 (.I0(n2839), .I1(n8874), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n9151));   // coms.v(517[9:65])
    defparam i1_2_lut_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_904 (.I0(\data_out[5] [2]), .I1(data_out_5__5__N_950), 
            .I2(\data_out[3][5] ), .I3(GND_net), .O(n6_adj_2467));   // coms.v(113[16:37])
    defparam i1_2_lut_3_lut_adj_904.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_905 (.I0(tx_transmit_N_2239[6]), .I1(tx_transmit_N_2239[4]), 
            .I2(tx_transmit_N_2239[5]), .I3(tx_transmit_N_2239[7]), .O(n8550));   // coms.v(330[10:53])
    defparam i3_4_lut_adj_905.LUT_INIT = 16'hfffe;
    SB_LUT4 i13959_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10111));   // coms.v(377[7:20])
    defparam i13959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_906 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(n9345), .I3(GND_net), .O(n17532));   // coms.v(128[17:30])
    defparam i1_2_lut_3_lut_adj_906.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame2_0___i72 (.Q(\data_out_frame2[8] [7]), .C(CLK_c), 
           .D(n10523));   // coms.v(428[12] 532[6])
    SB_LUT4 i4_3_lut_4_lut_adj_907 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(n8666), .I3(n17605), .O(n11_adj_2453));   // coms.v(128[17:30])
    defparam i4_3_lut_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n10121));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i71 (.Q(\data_out_frame2[8] [6]), .C(CLK_c), 
           .D(n10522));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_908 (.I0(tx_transmit_N_2239[3]), .I1(n8550), .I2(GND_net), 
            .I3(GND_net), .O(n121));   // coms.v(294[31:54])
    defparam i1_2_lut_adj_908.LUT_INIT = 16'heeee;
    SB_DFFE \data_out_9[[6__3519  (.Q(\data_out[9] [6]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__6__N_386));   // coms.v(274[12] 374[6])
    SB_DFF data_out_frame2_0___i70 (.Q(\data_out_frame2[8] [5]), .C(CLK_c), 
           .D(n10521));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i69 (.Q(\data_out_frame2[8] [4]), .C(CLK_c), 
           .D(n10520));   // coms.v(428[12] 532[6])
    SB_LUT4 i13958_3_lut (.I0(\data_in[3][7] ), .I1(\data_in[4][7] ), .I2(rx_data_ready), 
            .I3(GND_net), .O(n9939));   // coms.v(377[7:20])
    defparam i13958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_909 (.I0(n2594), .I1(n8061), .I2(n9100), .I3(n2588), 
            .O(n18_adj_2468));
    defparam i2_4_lut_adj_909.LUT_INIT = 16'hde7b;
    SB_LUT4 i10_4_lut_adj_910 (.I0(n2586), .I1(n20_adj_2452), .I2(n17534), 
            .I3(n8857), .O(n26_adj_2469));
    defparam i10_4_lut_adj_910.LUT_INIT = 16'hfdfe;
    SB_LUT4 i11059_2_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n2649[0]));   // coms.v(277[4] 373[11])
    defparam i11059_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i81 (.Q(\data_in[10] [0]), .C(CLK_c), .D(n10404));   // coms.v(402[9] 410[5])
    SB_LUT4 i13630_3_lut (.I0(\data_in[7]_c [4]), .I1(\data_in[8] [4]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10384));   // coms.v(377[7:20])
    defparam i13630_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i12 (.Q(\data_in[1]_c [3]), .C(CLK_c), .D(n10120));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i68 (.Q(\data_out_frame2[8] [3]), .C(CLK_c), 
           .D(n10519));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i67 (.Q(\data_out_frame2[8] [2]), .C(CLK_c), 
           .D(n10518));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i80 (.Q(\data_in[9] [7]), .C(CLK_c), .D(n10403));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i66 (.Q(\data_out_frame2[8] [1]), .C(CLK_c), 
           .D(n10517));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i65 (.Q(\data_out_frame2[8] [0]), .C(CLK_c), 
           .D(n10516));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i64 (.Q(\data_out_frame2[7] [7]), .C(CLK_c), 
           .D(n10515));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1][4] ), .C(CLK_c), .D(n10119));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_4_lut_adj_911 (.I0(\data_out[8] [5]), .I1(n8970), .I2(\data_out[7] [2]), 
            .I3(n17600), .O(data_out_9__6__N_386));   // coms.v(181[16:29])
    defparam i2_3_lut_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_912 (.I0(delay_counter[4]), .I1(delay_counter[1]), 
            .I2(delay_counter[3]), .I3(delay_counter[2]), .O(n17387));
    defparam i3_4_lut_adj_912.LUT_INIT = 16'hfffe;
    SB_DFF data_in_0___i14 (.Q(\data_in[1][5] ), .C(CLK_c), .D(n10118));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_4_lut_adj_913 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[2] [6]), .O(n17467));   // coms.v(230[15:344])
    defparam i2_3_lut_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n21_adj_2465), .I1(n23_adj_2462), .I2(n22_adj_2461), 
            .I3(n24_adj_2454), .O(n30));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_0___i79 (.Q(\data_in[9] [6]), .C(CLK_c), .D(n10402));   // coms.v(402[9] 410[5])
    SB_LUT4 i13438_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3][2] ), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10113));   // coms.v(377[7:20])
    defparam i13438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[9] [5]), .I1(n17433), .I2(n10_adj_2470), 
            .I3(n17409), .O(n17618));   // coms.v(235[16:323])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_914 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[4] [2]), 
            .I2(n17442), .I3(n17507), .O(n8687));   // coms.v(230[15:344])
    defparam i2_3_lut_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i9439_3_lut (.I0(delay_counter[5]), .I1(n18012), .I2(n1314), 
            .I3(GND_net), .O(n10686));
    defparam i9439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_915 (.I0(n8550), .I1(tx_transmit_N_2239[3]), .I2(n149), 
            .I3(GND_net), .O(n119));
    defparam i1_3_lut_adj_915.LUT_INIT = 16'heaea;
    SB_LUT4 add_3776_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n16350), .O(tx_transmit_N_2239_c[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_916 (.I0(n17), .I1(n30), .I2(n26_adj_2469), 
            .I3(n18_adj_2468), .O(n1_adj_2443));
    defparam i15_4_lut_adj_916.LUT_INIT = 16'hfffe;
    SB_LUT4 i13963_3_lut (.I0(\data_in[2]_c [0]), .I1(\data_in[3] [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10115));   // coms.v(377[7:20])
    defparam i13963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n81), .I1(n157), .I2(n142), .I3(\data_out_frame2[0] [7]), 
            .O(n9662));   // coms.v(422[11:16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h4f44;
    SB_DFFE \data_out_9[[5__3520  (.Q(\data_out[9] [5]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__5__N_401));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1][6] ), .C(CLK_c), .D(n10117));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_4_lut_adj_917 (.I0(n97), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n121), .I3(n8529), .O(n16450));
    defparam i2_4_lut_adj_917.LUT_INIT = 16'h3200;
    SB_LUT4 i1_3_lut_4_lut_adj_918 (.I0(n81), .I1(n157), .I2(n142), .I3(\data_out_frame2[0] [6]), 
            .O(n9665));   // coms.v(422[11:16])
    defparam i1_3_lut_4_lut_adj_918.LUT_INIT = 16'h4f44;
    SB_LUT4 i1_3_lut_4_lut_adj_919 (.I0(n81), .I1(n157), .I2(n142), .I3(\data_out_frame2[0] [5]), 
            .O(n9668));   // coms.v(422[11:16])
    defparam i1_3_lut_4_lut_adj_919.LUT_INIT = 16'h4f44;
    SB_LUT4 i1_4_lut_adj_920 (.I0(n16450), .I1(n119), .I2(n17387), .I3(n8486), 
            .O(n4));
    defparam i1_4_lut_adj_920.LUT_INIT = 16'haeaa;
    SB_LUT4 i9443_3_lut (.I0(delay_counter[8]), .I1(n18011), .I2(n1314), 
            .I3(GND_net), .O(n10680));
    defparam i9443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_921 (.I0(\data_in_frame[9] [5]), .I1(n17433), 
            .I2(n17594), .I3(GND_net), .O(n17619));   // coms.v(235[16:323])
    defparam i1_2_lut_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_922 (.I0(n81), .I1(n157), .I2(n142), .I3(\data_out_frame2[0] [1]), 
            .O(n9680));   // coms.v(422[11:16])
    defparam i1_3_lut_4_lut_adj_922.LUT_INIT = 16'h4f44;
    SB_DFFE \data_out_9[[4__3521  (.Q(\data_out[9] [4]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__4__N_414));   // coms.v(274[12] 374[6])
    SB_LUT4 i1_3_lut_4_lut_adj_923 (.I0(n81), .I1(n157), .I2(n142), .I3(\data_out_frame2[0] [0]), 
            .O(n9685));   // coms.v(422[11:16])
    defparam i1_3_lut_4_lut_adj_923.LUT_INIT = 16'h4f44;
    SB_LUT4 i15304_4_lut (.I0(delay_counter[9]), .I1(delay_counter[7]), 
            .I2(delay_counter[11]), .I3(delay_counter[6]), .O(n17753));
    defparam i15304_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15306_4_lut (.I0(delay_counter[5]), .I1(delay_counter[12]), 
            .I2(delay_counter[10]), .I3(delay_counter[8]), .O(n17755));
    defparam i15306_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame2_0___i63 (.Q(\data_out_frame2[7] [6]), .C(CLK_c), 
           .D(n10514));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i78 (.Q(\data_in[9] [5]), .C(CLK_c), .D(n10401));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i16 (.Q(\data_in[1][7] ), .C(CLK_c), .D(n10116));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i62 (.Q(\data_out_frame2[7] [5]), .C(CLK_c), 
           .D(n10513));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i77 (.Q(\data_in[9] [4]), .C(CLK_c), .D(n10400));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i61 (.Q(\data_out_frame2[7] [4]), .C(CLK_c), 
           .D(n10512));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i76 (.Q(\data_in[9] [3]), .C(CLK_c), .D(n10399));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_3_lut_adj_924 (.I0(n17312), .I1(n17755), .I2(n17753), .I3(GND_net), 
            .O(n17349));
    defparam i1_3_lut_adj_924.LUT_INIT = 16'h0202;
    SB_DFF data_in_0___i17 (.Q(\data_in[2]_c [0]), .C(CLK_c), .D(n10115));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i2 (.Q(\data_in[0][1] ), .C(CLK_c), .D(n9938));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i18 (.Q(\data_in[2][1] ), .C(CLK_c), .D(n10114));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n10113));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i60 (.Q(\data_out_frame2[7] [3]), .C(CLK_c), 
           .D(n10511));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i59 (.Q(\data_out_frame2[7] [2]), .C(CLK_c), 
           .D(n10510));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i58 (.Q(\data_out_frame2[7] [1]), .C(CLK_c), 
           .D(n10509));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i75 (.Q(\data_in[9] [2]), .C(CLK_c), .D(n10398));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i20 (.Q(\data_in[2][3] ), .C(CLK_c), .D(n10112));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i57 (.Q(\data_out_frame2[7] [0]), .C(CLK_c), 
           .D(n10508));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i74 (.Q(\data_in[9] [1]), .C(CLK_c), .D(n10397));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n10111));   // coms.v(402[9] 410[5])
    SB_LUT4 i3_4_lut_adj_925 (.I0(\data_out[8] [7]), .I1(n9091), .I2(n9087), 
            .I3(n17398), .O(data_out_9__4__N_414));   // coms.v(125[17:62])
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter2_2272__i7 (.Q(byte_transmit_counter2[7]), 
            .C(CLK_c), .E(n9605), .D(n37[7]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_DFF data_out_frame2_0___i56 (.Q(\data_out_frame2[6] [7]), .C(CLK_c), 
           .D(n10507));   // coms.v(428[12] 532[6])
    SB_DFFESR byte_transmit_counter2_2272__i6 (.Q(byte_transmit_counter2[6]), 
            .C(CLK_c), .E(n9605), .D(n37[6]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_LUT4 i12308_3_lut (.I0(n1_adj_2443), .I1(n5_adj_2438), .I2(\FRAME_MATCHER.state [0]), 
            .I3(GND_net), .O(n81));   // coms.v(422[11:16])
    defparam i12308_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame2_0___i55 (.Q(\data_out_frame2[6] [6]), .C(CLK_c), 
           .D(n10506));   // coms.v(428[12] 532[6])
    SB_DFFESR byte_transmit_counter2_2272__i5 (.Q(byte_transmit_counter2[5]), 
            .C(CLK_c), .E(n9605), .D(n37[5]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_DFF data_out_frame2_0___i54 (.Q(\data_out_frame2[6] [5]), .C(CLK_c), 
           .D(n10505));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2][5] ), .C(CLK_c), .D(n10110));   // coms.v(402[9] 410[5])
    SB_LUT4 i12_4_lut_adj_926 (.I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2239_c[0]), 
            .I2(n9631), .I3(n17349), .O(n16856));   // coms.v(19[11:32])
    defparam i12_4_lut_adj_926.LUT_INIT = 16'h0aca;
    SB_LUT4 i9040_3_lut (.I0(\data_in[1][6] ), .I1(\data_in[2][6] ), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10117));   // coms.v(377[7:20])
    defparam i9040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_927 (.I0(n1396), .I1(n15927), .I2(GND_net), .I3(GND_net), 
            .O(n9984));
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h4444;
    SB_DFFESR byte_transmit_counter2_2272__i4 (.Q(byte_transmit_counter2[4]), 
            .C(CLK_c), .E(n9605), .D(n37[4]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_DFF data_out_frame2_0___i53 (.Q(\data_out_frame2[6] [4]), .C(CLK_c), 
           .D(n10504));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i52 (.Q(\data_out_frame2[6] [3]), .C(CLK_c), 
           .D(n10503));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2][6] ), .C(CLK_c), .D(n10109));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_928 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[9] [3]), .I3(\data_in_frame[9] [5]), .O(n17418));   // coms.v(229[15:344])
    defparam i1_2_lut_3_lut_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_out[8] [4]), .I1(\data_out[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17620));   // coms.v(21[11:19])
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_930 (.I0(data_out_6__5__N_752), .I1(n17454), .I2(\data_out[6] [5]), 
            .I3(n17620), .O(data_out_9__5__N_401));   // coms.v(21[11:19])
    defparam i3_4_lut_adj_930.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_931 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [3]), 
            .I2(n8857), .I3(n9208), .O(n17541));   // coms.v(226[15:362])
    defparam i2_3_lut_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i24 (.Q(\data_in[2][7] ), .C(CLK_c), .D(n10108));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_adj_932 (.I0(\data_in[1] [2]), .I1(\data_in[1] [1]), 
            .I2(\data_in[3][6] ), .I3(GND_net), .O(n8572));   // coms.v(435[16:89])
    defparam i2_3_lut_adj_932.LUT_INIT = 16'hfbfb;
    SB_LUT4 i9441_3_lut (.I0(delay_counter[12]), .I1(n18009), .I2(n1314), 
            .I3(GND_net), .O(n10676));
    defparam i9441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17406));   // coms.v(71[16:45])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15930 (.I0(byte_transmit_counter2[2]), 
            .I1(n17815), .I2(n17818), .I3(byte_transmit_counter2[3]), 
            .O(n18372));
    defparam byte_transmit_counter2_2__bdd_4_lut_15930.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15921 (.I0(byte_transmit_counter2[2]), 
            .I1(n17824), .I2(n17827), .I3(byte_transmit_counter2[3]), 
            .O(n18366));
    defparam byte_transmit_counter2_2__bdd_4_lut_15921.LUT_INIT = 16'he4aa;
    SB_LUT4 i15249_2_lut (.I0(\data_in[0] [7]), .I1(\data_in[1]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17697));
    defparam i15249_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n10107));   // coms.v(402[9] 410[5])
    SB_LUT4 i5_4_lut_adj_934 (.I0(\data_in[2] [4]), .I1(\data_in[3][3] ), 
            .I2(\data_in[2][6] ), .I3(\data_in[2][1] ), .O(n12_adj_2472));   // coms.v(440[16:93])
    defparam i5_4_lut_adj_934.LUT_INIT = 16'hfffe;
    SB_LUT4 i15315_4_lut (.I0(\data_in[1][5] ), .I1(\data_in[0][4] ), .I2(\data_in[1]_c [0]), 
            .I3(n17697), .O(n17765));
    defparam i15315_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_935 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[10] [3]), .I3(GND_net), .O(n17433));   // coms.v(229[15:344])
    defparam i1_2_lut_3_lut_adj_935.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n17218));   // coms.v(446[4] 531[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i9437_3_lut (.I0(\delay_counter[13] ), .I1(n18008), .I2(n1314), 
            .I3(GND_net), .O(n10675));
    defparam i9437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_936 (.I0(n2839), .I1(\data_in_frame[3] [0]), .I2(\data_in_frame[4] [4]), 
            .I3(n17406), .O(n17656));   // coms.v(517[9:65])
    defparam i1_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i9397_3_lut (.I0(\delay_counter[14] ), .I1(n18105), .I2(n1314), 
            .I3(GND_net), .O(n10674));
    defparam i9397_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3776_3 (.CI(n16350), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n16351));
    SB_DFF data_in_0___i26 (.Q(\data_in[3][1] ), .C(CLK_c), .D(n10106));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i27 (.Q(\data_in[3][2] ), .C(CLK_c), .D(n10105));   // coms.v(402[9] 410[5])
    SB_LUT4 add_3776_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(n251), .I3(GND_net), .O(tx_transmit_N_2239_c[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_937 (.I0(n17765), .I1(n12_adj_2472), .I2(\data_in[0][2] ), 
            .I3(\data_in[3][1] ), .O(n8556));   // coms.v(440[16:93])
    defparam i6_4_lut_adj_937.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_4_lut_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n142), .I2(GND_net), 
            .I3(GND_net), .O(n17214));   // coms.v(446[4] 531[11])
    defparam i2_4_lut_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i28 (.Q(\data_in[3][3] ), .C(CLK_c), .D(n10104));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_adj_938 (.I0(\data_in_frame[1][1] ), .I1(n17656), .I2(GND_net), 
            .I3(GND_net), .O(n17529));   // coms.v(71[16:45])
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_LUT4 i15266_3_lut (.I0(\data_in[0][1] ), .I1(\data_in[2][5] ), .I2(\data_in[2][7] ), 
            .I3(GND_net), .O(n17715));
    defparam i15266_3_lut.LUT_INIT = 16'h8080;
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n10103));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_adj_939 (.I0(n17516), .I1(n8976), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n8886));
    defparam i2_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 i15907_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n142));   // coms.v(446[4] 531[11])
    defparam i15907_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i3869_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [7]), .I3(\data_in_frame[10] [7]), .O(n2560));   // coms.v(435[13] 445[7])
    defparam i3869_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_0___i30 (.Q(\data_in[3][5] ), .C(CLK_c), .D(n10102));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_in[3][7] ), .I1(\data_in[0]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2473));   // coms.v(440[16:93])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_941 (.I0(\data_in[2]_c [0]), .I1(n6_adj_2473), 
            .I2(n17715), .I3(\data_in[2] [2]), .O(n8_adj_2474));   // coms.v(440[16:93])
    defparam i3_4_lut_adj_941.LUT_INIT = 16'hdfff;
    SB_LUT4 i10279_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [6]), .I3(\data_in_frame[10][6] ), .O(n2561));   // coms.v(435[13] 445[7])
    defparam i10279_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_3776_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(n251), 
            .CO(n16350));
    SB_LUT4 i3889_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [5]), .I3(\data_in_frame[9] [5]), .O(n2570));   // coms.v(435[13] 445[7])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [5]), .I3(\data_in_frame[10] [5]), .O(n2562));   // coms.v(435[13] 445[7])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10201_3_lut (.I0(\data_in[1]_c [3]), .I1(\data_in[2][3] ), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10120));   // coms.v(377[7:20])
    defparam i10201_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i33 (.Q(\data_in[4][0] ), .C(CLK_c), .D(n10101));   // coms.v(402[9] 410[5])
    SB_DFFESR byte_transmit_counter2_2272__i3 (.Q(byte_transmit_counter2[3]), 
            .C(CLK_c), .E(n9605), .D(n37[3]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_DFFESR byte_transmit_counter2_2272__i2 (.Q(byte_transmit_counter2[2]), 
            .C(CLK_c), .E(n9605), .D(n37[2]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_DFF data_in_0___i38 (.Q(\data_in[4][5] ), .C(CLK_c), .D(n10100));   // coms.v(402[9] 410[5])
    SB_LUT4 n18366_bdd_4_lut (.I0(n18366), .I1(n6_adj_2466), .I2(n18084), 
            .I3(byte_transmit_counter2[3]), .O(n18369));
    defparam n18366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR byte_transmit_counter2_2272__i1 (.Q(byte_transmit_counter2[1]), 
            .C(CLK_c), .E(n9605), .D(n37[1]), .R(n9900));   // coms.v(489[6] 497[9])
    SB_LUT4 i46_2_lut (.I0(\data_in[1][7] ), .I1(\data_in[0]_c [3]), .I2(GND_net), 
            .I3(GND_net), .O(n28_adj_2475));
    defparam i46_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \data_out_8[[0__3533  (.Q(\data_out[8] [0]), .C(CLK_c), .D(n10361));   // coms.v(274[12] 374[6])
    SB_LUT4 i3875_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [4]), .I3(\data_in_frame[10] [4]), .O(n2563));   // coms.v(435[13] 445[7])
    defparam i3875_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3877_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [3]), .I3(\data_in_frame[10] [3]), .O(n2564));   // coms.v(435[13] 445[7])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [2]), .I3(\data_in_frame[10] [2]), .O(n2565));   // coms.v(435[13] 445[7])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_0___i35 (.Q(\data_in[4][2] ), .C(CLK_c), .D(n10099));   // coms.v(402[9] 410[5])
    SB_DFF data_out_frame2_0___i51 (.Q(\data_out_frame2[6] [2]), .C(CLK_c), 
           .D(n10502));   // coms.v(428[12] 532[6])
    SB_LUT4 i3881_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [1]), .I3(\data_in_frame[10] [1]), .O(n2566));   // coms.v(435[13] 445[7])
    defparam i3881_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3883_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[10] [0]), .I3(\data_in_frame[10] [0]), .O(n2567));   // coms.v(435[13] 445[7])
    defparam i3883_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_out_frame2_0___i50 (.Q(\data_out_frame2[6] [1]), .C(CLK_c), 
           .D(n10501));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i49 (.Q(\data_out_frame2[6] [0]), .C(CLK_c), 
           .D(n10500));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i48 (.Q(\data_out_frame2[5] [7]), .C(CLK_c), 
           .D(n10499));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i47 (.Q(\data_out_frame2[5] [6]), .C(CLK_c), 
           .D(n10498));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i46 (.Q(\data_out_frame2[5] [5]), .C(CLK_c), 
           .D(n10497));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i45 (.Q(\data_out_frame2[5] [4]), .C(CLK_c), 
           .D(n10496));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i44 (.Q(\data_out_frame2[5] [3]), .C(CLK_c), 
           .D(n10495));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i43 (.Q(\data_out_frame2[5] [2]), .C(CLK_c), 
           .D(n10494));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i42 (.Q(\data_out_frame2[5] [1]), .C(CLK_c), 
           .D(n10493));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i41 (.Q(\data_out_frame2[5] [0]), .C(CLK_c), 
           .D(n10492));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i168 (.Q(\data_in[20] [7]), .C(CLK_c), .D(n10491));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i167 (.Q(\data_in[20] [6]), .C(CLK_c), .D(n10490));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i166 (.Q(\data_in[20] [5]), .C(CLK_c), .D(n10489));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i165 (.Q(\data_in[20] [4]), .C(CLK_c), .D(n10488));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i164 (.Q(\data_in[20] [3]), .C(CLK_c), .D(n10487));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i163 (.Q(\data_in[20] [2]), .C(CLK_c), .D(n10486));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i162 (.Q(\data_in[20] [1]), .C(CLK_c), .D(n10485));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i161 (.Q(\data_in[20] [0]), .C(CLK_c), .D(n10484));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i160 (.Q(\data_in[19] [7]), .C(CLK_c), .D(n10483));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i159 (.Q(\data_in[19] [6]), .C(CLK_c), .D(n10482));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i158 (.Q(\data_in[19] [5]), .C(CLK_c), .D(n10481));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i157 (.Q(\data_in[19] [4]), .C(CLK_c), .D(n10480));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i156 (.Q(\data_in[19] [3]), .C(CLK_c), .D(n10479));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i155 (.Q(\data_in[19] [2]), .C(CLK_c), .D(n10478));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i154 (.Q(\data_in[19] [1]), .C(CLK_c), .D(n10477));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i153 (.Q(\data_in[19] [0]), .C(CLK_c), .D(n10476));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i152 (.Q(\data_in[18] [7]), .C(CLK_c), .D(n10475));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i151 (.Q(\data_in[18] [6]), .C(CLK_c), .D(n10474));   // coms.v(402[9] 410[5])
    SB_DFFE \data_out_9[[3__3522  (.Q(\data_out[9] [3]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__3__N_430));   // coms.v(274[12] 374[6])
    SB_LUT4 i3893_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [3]), .I3(\data_in_frame[9] [3]), .O(n2572));   // coms.v(435[13] 445[7])
    defparam i3893_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_0___i65 (.Q(\data_in[8] [0]), .C(CLK_c), .D(n10388));   // coms.v(402[9] 410[5])
    SB_LUT4 i9042_3_lut (.I0(\data_in[0]_c [0]), .I1(\data_in[1]_c [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10122));   // coms.v(377[7:20])
    defparam i9042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3897_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [1]), .I3(\data_in_frame[9] [1]), .O(n2574));   // coms.v(435[13] 445[7])
    defparam i3897_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n142), .O(n17216));
    defparam i2_3_lut_2_lut.LUT_INIT = 16'h00aa;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15916 (.I0(byte_transmit_counter2[2]), 
            .I1(n17833), .I2(n17836), .I3(byte_transmit_counter2[3]), 
            .O(n18360));
    defparam byte_transmit_counter2_2__bdd_4_lut_15916.LUT_INIT = 16'he4aa;
    SB_LUT4 i13614_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [6]), .I3(\data_in_frame[9][6] ), .O(n15927));   // coms.v(435[13] 445[7])
    defparam i13614_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n18390_bdd_4_lut (.I0(n18390), .I1(n18095), .I2(n18094), .I3(\byte_transmit_counter[2] ), 
            .O(n18393));
    defparam n18390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \data_out_9[[2__3523  (.Q(\data_out[9] [2]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__2__N_446));   // coms.v(274[12] 374[6])
    SB_LUT4 i1_2_lut_3_lut_adj_942 (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(n1396), .I3(GND_net), .O(n9419));   // coms.v(435[13] 445[7])
    defparam i1_2_lut_3_lut_adj_942.LUT_INIT = 16'hf4f4;
    SB_LUT4 i3885_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [7]), .I3(\data_in_frame[9] [7]), .O(n2568));   // coms.v(435[13] 445[7])
    defparam i3885_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10244_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [2]), .I3(\data_in_frame[9] [2]), .O(n2573));   // coms.v(435[13] 445[7])
    defparam i10244_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3899_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [0]), .I3(\data_in_frame[9] [0]), .O(n2575));   // coms.v(435[13] 445[7])
    defparam i3899_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13622_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[9] [4]), .I3(\data_in_frame[9] [4]), .O(n2571));   // coms.v(435[13] 445[7])
    defparam i13622_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_0___i150 (.Q(\data_in[18] [5]), .C(CLK_c), .D(n10473));   // coms.v(402[9] 410[5])
    SB_DFFE \data_out_9[[1__3524  (.Q(\data_out[9] [1]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__1__N_462));   // coms.v(274[12] 374[6])
    SB_DFFE \data_out_9[[0__3525  (.Q(\data_out[9] [0]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_9__0__N_475));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i149 (.Q(\data_in[18] [4]), .C(CLK_c), .D(n10472));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_4_lut_adj_943 (.I0(\data_in[3][5] ), .I1(n28_adj_2475), .I2(n8_adj_2474), 
            .I3(\data_in[1][6] ), .O(n8559));   // coms.v(440[16:93])
    defparam i1_4_lut_adj_943.LUT_INIT = 16'hfffb;
    SB_LUT4 i15742_2_lut (.I0(data_out_5__5__N_950), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18092));
    defparam i15742_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7621_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[1]), .I3(delay_counter[1]), 
            .O(n10037));
    defparam i7621_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i15743_2_lut (.I0(\data_out[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18093));
    defparam i15743_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i148 (.Q(\data_in[18] [3]), .C(CLK_c), .D(n10471));   // coms.v(402[9] 410[5])
    SB_LUT4 i7626_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[2]), .I3(delay_counter[2]), 
            .O(n10042));
    defparam i7626_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 add_3777_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n16307), .O(n7260[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \data_out_10[[7__3510  (.Q(\data_out[10] [7]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__7__N_101));   // coms.v(274[12] 374[6])
    SB_LUT4 i7631_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[3]), .I3(delay_counter[3]), 
            .O(n10047));
    defparam i7631_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i7634_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[4]), .I3(delay_counter[4]), 
            .O(n10050));
    defparam i7634_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i15784_2_lut (.I0(\data_out[0][5] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18091));
    defparam i15784_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15805_3_lut (.I0(\data_out_frame2[0] [0]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n18074));
    defparam i15805_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i2_3_lut (.I0(data_out_6__7__N_678), 
            .I1(\data_out[3][5] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2476));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \data_out_10[[6__3511  (.Q(\data_out[10] [6]), .C(CLK_c), .E(data_out_10__7__N_114), 
            .D(data_out_10__6__N_118));   // coms.v(274[12] 374[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame2[6] [0]), 
            .I1(\data_out_frame2[7] [0]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2477));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3777_2 (.CI(VCC_net), .I0(\delay_counter[0] ), .I1(GND_net), 
            .CO(n16305));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame2[5] [0]), 
            .I1(n5_adj_2477), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2436));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_in[0][6] ), .I1(n8556), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_2478));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'heeee;
    SB_LUT4 i7640_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[6]), .I3(delay_counter[6]), 
            .O(n10056));
    defparam i7640_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i15294_4_lut (.I0(\data_in[3][2] ), .I1(\data_in[0][5] ), .I2(\data_in[3] [4]), 
            .I3(\data_in[3] [0]), .O(n17743));
    defparam i15294_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_out_frame2_0___i2 (.Q(\data_out_frame2[0] [1]), .C(CLK_c), 
           .D(n9680));   // coms.v(428[12] 532[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15965 (.I0(byte_transmit_counter[1]), 
            .I1(n17949), .I2(n5_adj_2444), .I3(\byte_transmit_counter[2] ), 
            .O(n18414));
    defparam byte_transmit_counter_1__bdd_4_lut_15965.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_945 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17550));   // coms.v(452[9:67])
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i3 (.Q(\data_out_frame2[0] [2]), .C(CLK_c), 
           .D(n9677));   // coms.v(428[12] 532[6])
    SB_LUT4 i4_4_lut_adj_946 (.I0(\data_in[1][4] ), .I1(n17743), .I2(\data_in[2][3] ), 
            .I3(n6_adj_2478), .O(n8460));
    defparam i4_4_lut_adj_946.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_2_lut (.I0(n8460), .I1(n8559), .I2(GND_net), .I3(GND_net), 
            .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_947 (.I0(n7), .I1(\data_in[3][6] ), .I2(\data_in[1] [1]), 
            .I3(\data_in[1] [2]), .O(n63_adj_9));
    defparam i4_4_lut_adj_947.LUT_INIT = 16'hfbff;
    SB_LUT4 i15296_4_lut (.I0(\data_in[3][5] ), .I1(\data_in[1][6] ), .I2(\data_in[3][7] ), 
            .I3(\data_in[0]_c [0]), .O(n17745));
    defparam i15296_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7643_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[7]), .I3(delay_counter[7]), 
            .O(n10059));
    defparam i7643_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i7649_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[9]), .I3(delay_counter[9]), 
            .O(n10065));
    defparam i7649_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_DFF data_out_frame2_0___i4 (.Q(\data_out_frame2[0] [3]), .C(CLK_c), 
           .D(n9674));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i5 (.Q(\data_out_frame2[0] [4]), .C(CLK_c), 
           .D(n9671));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i6 (.Q(\data_out_frame2[0] [5]), .C(CLK_c), 
           .D(n9668));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i7 (.Q(\data_out_frame2[0] [6]), .C(CLK_c), 
           .D(n9665));   // coms.v(428[12] 532[6])
    SB_DFF data_out_frame2_0___i8 (.Q(\data_out_frame2[0] [7]), .C(CLK_c), 
           .D(n9662));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i154 (.Q(\data_out_frame2[19] [1]), .C(CLK_c), 
            .E(n9606), .D(n17619));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i155 (.Q(\data_out_frame2[19] [2]), .C(CLK_c), 
            .E(n9606), .D(n17480));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i156 (.Q(\data_out_frame2[19] [3]), .C(CLK_c), 
            .E(n9606), .D(n17590));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i157 (.Q(\data_out_frame2[19] [4]), .C(CLK_c), 
            .E(n9606), .D(n17548));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i158 (.Q(\data_out_frame2[19] [5]), .C(CLK_c), 
            .E(n9606), .D(n17587));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i159 (.Q(\data_out_frame2[19] [6]), .C(CLK_c), 
            .E(n9606), .D(n17537));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i160 (.Q(\data_out_frame2[19] [7]), .C(CLK_c), 
            .E(n9606), .D(n17420));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i161 (.Q(\data_out_frame2[20] [0]), .C(CLK_c), 
            .E(n9606), .D(n17649));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i162 (.Q(\data_out_frame2[20] [1]), .C(CLK_c), 
            .E(n9606), .D(n17618));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i163 (.Q(\data_out_frame2[20] [2]), .C(CLK_c), 
            .E(n9606), .D(n17490));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i164 (.Q(\data_out_frame2[20] [3]), .C(CLK_c), 
            .E(n9606), .D(n17540));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i165 (.Q(\data_out_frame2[20] [4]), .C(CLK_c), 
            .E(n9606), .D(n17593));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i166 (.Q(\data_out_frame2[20] [5]), .C(CLK_c), 
            .E(n9606), .D(n17543));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i167 (.Q(\data_out_frame2[20] [6]), .C(CLK_c), 
            .E(n9606), .D(n17545));   // coms.v(428[12] 532[6])
    SB_DFFE data_out_frame2_0___i168 (.Q(\data_out_frame2[20] [7]), .C(CLK_c), 
            .E(n9606), .D(n17584));   // coms.v(428[12] 532[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
            .D(n17216), .S(n1_adj_2437));   // coms.v(428[12] 532[6])
    SB_DFFSS \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
            .D(n17218), .S(n4_adj_2480));   // coms.v(428[12] 532[6])
    SB_DFF \data_out_8[[1__3532  (.Q(\data_out[8] [1]), .C(CLK_c), .D(n10360));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[2__3531  (.Q(\data_out[8] [2]), .C(CLK_c), .D(n10359));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[3__3530  (.Q(\data_out[8] [3]), .C(CLK_c), .D(n10358));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[4__3529  (.Q(\data_out[8] [4]), .C(CLK_c), .D(n10357));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[5__3528  (.Q(\data_out[8] [5]), .C(CLK_c), .D(n10353));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[6__3527  (.Q(\data_out[8] [6]), .C(CLK_c), .D(n10352));   // coms.v(274[12] 374[6])
    SB_DFF \data_out_8[[7__3526  (.Q(\data_out[8] [7]), .C(CLK_c), .D(n10351));   // coms.v(274[12] 374[6])
    SB_DFF data_in_0___i36 (.Q(\data_in[4][3] ), .C(CLK_c), .D(n10347));   // coms.v(402[9] 410[5])
    SB_LUT4 i7652_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[10]), .I3(delay_counter[10]), 
            .O(n10068));
    defparam i7652_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_DFF data_in_0___i9 (.Q(\data_in[1]_c [0]), .C(CLK_c), .D(n10342));   // coms.v(402[9] 410[5])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), 
           .D(n10266));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), 
           .D(n10269));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), 
           .D(n10272));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), 
           .D(n10276));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), 
           .D(n10279));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), 
           .D(n10333));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i147 (.Q(\data_in[18] [2]), .C(CLK_c), .D(n10470));   // coms.v(402[9] 410[5])
    SB_LUT4 add_3777_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n16305), .O(n7260[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i146 (.Q(\data_in[18] [1]), .C(CLK_c), .D(n10469));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i145 (.Q(\data_in[18] [0]), .C(CLK_c), .D(n10468));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i144 (.Q(\data_in[17] [7]), .C(CLK_c), .D(n10467));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i143 (.Q(\data_in[17] [6]), .C(CLK_c), .D(n10466));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i31 (.Q(\data_in[3][6] ), .C(CLK_c), .D(n10330));   // coms.v(402[9] 410[5])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), 
           .D(n10286));   // coms.v(428[12] 532[6])
    SB_LUT4 i7655_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[11]), .I3(delay_counter[11]), 
            .O(n10071));
    defparam i7655_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i3_4_lut_adj_948 (.I0(\data_in_frame[3] [6]), .I1(n17550), .I2(n17442), 
            .I3(n17553), .O(n8674));   // coms.v(383[12:25])
    defparam i3_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out[6] [5]), 
            .I1(\data_out[7] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2481));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15694_2_lut (.I0(data_out_7__5__N_543), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17943));
    defparam i15694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_949 (.I0(n8970), .I1(n17626), .I2(n17608), .I3(n17662), 
            .O(n12_adj_2482));   // coms.v(181[16:29])
    defparam i5_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_950 (.I0(n17665), .I1(n12_adj_2482), .I2(\data_out[8] [6]), 
            .I3(\data_out[7] [3]), .O(data_out_9__7__N_323));   // coms.v(181[16:29])
    defparam i6_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_951 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[6] [1]), .I3(GND_net), .O(n9208));   // coms.v(227[15:353])
    defparam i1_2_lut_3_lut_adj_951.LUT_INIT = 16'h9696;
    SB_LUT4 i7780_4_lut_4_lut (.I0(n1314), .I1(n29), .I2(n7260[0]), .I3(\delay_counter[0] ), 
            .O(n10196));
    defparam i7780_4_lut_4_lut.LUT_INIT = 16'hfb51;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17650));   // coms.v(230[15:344])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i15798_2_lut (.I0(\data_out[1][2] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18096));
    defparam i15798_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[9][6] ), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17559));   // coms.v(228[15:344])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_954 (.I0(n17629), .I1(n8725), .I2(n17467), .I3(GND_net), 
            .O(n8890));   // coms.v(69[15:74])
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i64 (.Q(\data_in[7][7] ), .C(CLK_c), .D(n10387));   // coms.v(402[9] 410[5])
    SB_CARRY add_3777_9 (.CI(n16311), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n16312));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i2_3_lut (.I0(data_out_6__6__N_729), 
            .I1(data_out_5__4__N_959), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2483));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_955 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(n8890), .I3(n17559), .O(n9135));   // coms.v(228[15:344])
    defparam i3_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 n18414_bdd_4_lut (.I0(n18414), .I1(n18090), .I2(n1_adj_2484), 
            .I3(\byte_transmit_counter[2] ), .O(n18417));
    defparam n18414_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_220_Select_0_i1_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [2]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.next_state[0] ), .O(n1_c));
    defparam select_220_Select_0_i1_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFF data_in_0___i63 (.Q(\data_in[7][6] ), .C(CLK_c), .D(n10386));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15960 (.I0(byte_transmit_counter2[2]), 
            .I1(n17794), .I2(n17797), .I3(byte_transmit_counter2[3]), 
            .O(n18408));
    defparam byte_transmit_counter2_2__bdd_4_lut_15960.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_956 (.I0(\data_in[2][7] ), .I1(n8572), .I2(\data_in[2] [2]), 
            .I3(n8460), .O(n16_adj_2485));   // coms.v(435[16:89])
    defparam i6_4_lut_adj_956.LUT_INIT = 16'hfffe;
    SB_LUT4 i15815_2_lut (.I0(\data_out[0][0] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18088));
    defparam i15815_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_957 (.I0(\data_in[2][5] ), .I1(\data_in[2]_c [0]), 
            .I2(\data_in[0][1] ), .I3(\data_in[1][7] ), .O(n17_adj_2486));   // coms.v(435[16:89])
    defparam i7_4_lut_adj_957.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [4]), 
            .I2(n9219), .I3(n8063), .O(n17544));   // coms.v(227[15:353])
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i2_3_lut (.I0(\data_out[2][0] ), 
            .I1(data_out_6__2__N_804), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2487));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out[6] [0]), 
            .I1(\data_out[7] [0]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2488));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_959 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(n10_adj_2430), .I3(\data_in_frame[2] [3]), .O(n8695));   // coms.v(383[12:25])
    defparam i5_3_lut_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i15728_2_lut (.I0(data_out_6__3__N_788), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17911));
    defparam i15728_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \FRAME_MATCHER.next_state_i0  (.Q(\FRAME_MATCHER.next_state[0] ), 
           .C(CLK_c), .D(n17092));   // coms.v(428[12] 532[6])
    SB_DFF data_in_0___i142 (.Q(\data_in[17] [5]), .C(CLK_c), .D(n10465));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_in_frame[5] [6]), .I1(n8687), .I2(GND_net), 
            .I3(GND_net), .O(n8063));   // coms.v(119[16:83])
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_961 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n9349));   // coms.v(452[9:67])
    defparam i2_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_962 (.I0(n9349), .I1(n30_adj_2489), .I2(n9334), 
            .I3(GND_net), .O(n17476));   // coms.v(452[9:67])
    defparam i2_3_lut_adj_962.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out[6] [3]), 
            .I1(\data_out[7] [3]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2490));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15801_2_lut (.I0(\data_out[5] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17937));
    defparam i15801_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_963 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(n8874), .I3(n9349), .O(n9368));   // coms.v(128[17:38])
    defparam i3_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_964 (.I0(n25_adj_2491), .I1(n17507), .I2(n9163), 
            .I3(n17602), .O(n12_adj_2492));   // coms.v(517[9:65])
    defparam i5_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_965 (.I0(n17656), .I1(n12_adj_2492), .I2(\data_in_frame[2] [2]), 
            .I3(\data_in_frame[0] [1]), .O(n9334));   // coms.v(517[9:65])
    defparam i6_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i15874_4_lut_4_lut_4_lut (.I0(\UART_TRANSMITTER.state[0] ), .I1(n4430), 
            .I2(GND_net), .I3(GND_net), .O(n9519));   // coms.v(277[4] 373[11])
    defparam i15874_4_lut_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_966 (.I0(n9334), .I1(n2600), .I2(n9365), .I3(n9368), 
            .O(n10_adj_2493));   // coms.v(76[16:93])
    defparam i4_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_967 (.I0(\data_in_frame[7][0] ), .I1(\data_in_frame[8] [6]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n9279));   // coms.v(224[15:379])
    defparam i1_2_lut_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_968 (.I0(n2597), .I1(n2601), .I2(n17575), .I3(n17516), 
            .O(n11_adj_2494));   // coms.v(452[9:67])
    defparam i3_4_lut_adj_968.LUT_INIT = 16'h7bde;
    SB_LUT4 i15831_3_lut (.I0(\data_out_frame2[0] [5]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n18080));
    defparam i15831_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i15819_3_lut (.I0(\data_out_frame2[0] [7]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n18076));
    defparam i15819_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame2[6] [5]), 
            .I1(\data_out_frame2[7] [5]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2495));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut (.I0(\data_out_frame2[5] [5]), 
            .I1(n5_adj_2495), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2496));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i2_3_lut_4_lut_adj_969 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[4] [4]), 
            .I2(n9043), .I3(n9283), .O(n6_adj_10));   // coms.v(383[12:25])
    defparam i2_3_lut_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n2593), .I1(n2595), .I2(n8687), .I3(n8674), 
            .O(n8_adj_2459));   // coms.v(452[9:67])
    defparam i1_4_lut_adj_970.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_971 (.I0(n2596), .I1(n2605), .I2(n8666), .I3(n17529), 
            .O(n10_adj_2498));   // coms.v(452[9:67])
    defparam i3_4_lut_adj_971.LUT_INIT = 16'hde7b;
    SB_LUT4 i7843_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1][7] ), 
            .I3(\data_in_frame[1] [7]), .O(n10259));
    defparam i7843_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out[6] [2]), 
            .I1(\data_out[7] [2]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2499));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_972 (.I0(n2607), .I1(n2602), .I2(n8751), .I3(n17513), 
            .O(n9_adj_2500));   // coms.v(452[9:67])
    defparam i2_4_lut_adj_972.LUT_INIT = 16'hde7b;
    SB_LUT4 i1_2_lut_3_lut_adj_973 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[4] [4]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n9058));   // coms.v(383[12:25])
    defparam i1_2_lut_3_lut_adj_973.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(tx2_transmit_N_2287), .O(n1_adj_2455));   // coms.v(428[12] 532[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i15731_2_lut (.I0(\data_out[5] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17936));
    defparam i15731_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_974 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n9219));   // coms.v(228[15:344])
    defparam i1_2_lut_3_lut_adj_974.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame2[6] [7]), 
            .I1(\data_out_frame2[7] [7]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2501));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut (.I0(\data_out_frame2[5] [7]), 
            .I1(n5_adj_2501), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2464));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i13629_3_lut (.I0(\data_in[4]_c [4]), .I1(\data_in[5] [4]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10143));   // coms.v(377[7:20])
    defparam i13629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15708_3_lut (.I0(\data_out_frame2[0] [1]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n18086));
    defparam i15708_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut_3_lut_adj_975 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[10][6] ), .I3(GND_net), .O(n6_adj_2502));   // coms.v(226[15:362])
    defparam i1_2_lut_3_lut_adj_975.LUT_INIT = 16'h9696;
    SB_LUT4 i7839_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1][6] ), 
            .I3(\data_in_frame[1] [6]), .O(n10255));
    defparam i7839_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_976 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[10] [7]), .I3(\data_in_frame[9] [1]), .O(n8989));   // coms.v(229[15:344])
    defparam i1_2_lut_3_lut_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame2[6] [1]), 
            .I1(\data_out_frame2[7] [1]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2503));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_977 (.I0(\data_in_frame[1] [7]), .I1(n9039), .I2(n2599), 
            .I3(n17476), .O(n17478));   // coms.v(76[16:93])
    defparam i3_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut (.I0(\data_out_frame2[5] [1]), 
            .I1(n5_adj_2503), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2504));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i7836_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1][5] ), 
            .I3(\data_in_frame[1] [5]), .O(n10252));
    defparam i7836_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_3_lut_adj_978 (.I0(n9204), .I1(\data_in_frame[5] [4]), 
            .I2(n8674), .I3(GND_net), .O(n17591));   // coms.v(226[15:362])
    defparam i1_2_lut_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_979 (.I0(n2594), .I1(n2603), .I2(n17569), .I3(n17424), 
            .O(n10_adj_2505));   // coms.v(452[9:67])
    defparam i2_4_lut_adj_979.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_4_lut_adj_980 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [6]), 
            .I2(n9144), .I3(n8064), .O(n17582));   // coms.v(229[15:344])
    defparam i2_3_lut_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_981 (.I0(n11_adj_2494), .I1(n2606), .I2(n17428), 
            .I3(n17522), .O(n14));   // coms.v(452[9:67])
    defparam i6_4_lut_adj_981.LUT_INIT = 16'hfbfe;
    SB_LUT4 n18408_bdd_4_lut (.I0(n18408), .I1(n6_adj_2506), .I2(n18078), 
            .I3(byte_transmit_counter2[3]), .O(n18411));
    defparam n18408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7895_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][6] ), 
            .I3(\data_in_frame[3] [6]), .O(n10311));
    defparam i7895_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_4_lut_adj_982 (.I0(n8867), .I1(n11_adj_2460), .I2(n9_adj_2500), 
            .I3(n10_adj_2498), .O(n17325));   // coms.v(452[9:67])
    defparam i1_4_lut_adj_982.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_983 (.I0(n17478), .I1(n17632), .I2(n2598), .I3(n17476), 
            .O(n9_adj_2507));   // coms.v(452[9:67])
    defparam i1_4_lut_adj_983.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_4_lut_adj_984 (.I0(n9_adj_2507), .I1(n17325), .I2(n14), 
            .I3(n10_adj_2505), .O(n31));   // coms.v(452[9:67])
    defparam i1_4_lut_adj_984.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_985 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(n17403), .I3(\data_in_frame[2] [6]), .O(n9283));   // coms.v(228[15:344])
    defparam i2_3_lut_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17614));   // coms.v(128[17:38])
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_2508));   // coms.v(383[12:25])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9186));   // coms.v(452[9:67])
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i7833_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1][4] ), 
            .I3(\data_in_frame[1] [4]), .O(n10249));
    defparam i7833_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i10211_3_lut (.I0(\data_in[0]_c [3]), .I1(\data_in[1]_c [3]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n9936));   // coms.v(377[7:20])
    defparam i10211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15817_3_lut (.I0(\data_out_frame2[0] [3]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n18082));
    defparam i15817_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1]_c [3]), 
            .I3(\data_in_frame[1] [3]), .O(n10242));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame2[6] [3]), 
            .I1(\data_out_frame2[7] [3]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2509));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7823_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[1] [2]), 
            .I3(\data_in_frame[1] [2]), .O(n10239));
    defparam i7823_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_4_lut_4_lut_adj_989 (.I0(n16468), .I1(n1396), .I2(\data_in[1] [1]), 
            .I3(\data_in_frame[1][1] ), .O(n10236));
    defparam i1_4_lut_4_lut_adj_989.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame2[5] [3]), 
            .I1(n5_adj_2509), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2432));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_in_0___i141 (.Q(\data_in[17] [4]), .C(CLK_c), .D(n10464));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i140 (.Q(\data_in[17] [3]), .C(CLK_c), .D(n10463));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i139 (.Q(\data_in[17] [2]), .C(CLK_c), .D(n10462));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i138 (.Q(\data_in[17] [1]), .C(CLK_c), .D(n10461));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i137 (.Q(\data_in[17] [0]), .C(CLK_c), .D(n10460));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i136 (.Q(\data_in[16] [7]), .C(CLK_c), .D(n10459));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i135 (.Q(\data_in[16] [6]), .C(CLK_c), .D(n10458));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i134 (.Q(\data_in[16] [5]), .C(CLK_c), .D(n10457));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_990 (.I0(data_out_5__4__N_959), .I1(data_out_6__2__N_804), 
            .I2(data_out_6__7__N_678), .I3(data_out_6__1__N_850), .O(n8964));   // coms.v(125[17:62])
    defparam i1_2_lut_3_lut_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i9091_3_lut (.I0(\data_in[4] [1]), .I1(\data_in[5] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10148));   // coms.v(377[7:20])
    defparam i9091_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i133 (.Q(\data_in[16] [4]), .C(CLK_c), .D(n10456));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i132 (.Q(\data_in[16] [3]), .C(CLK_c), .D(n10455));   // coms.v(402[9] 410[5])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), 
           .D(n10289));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), 
           .D(n10293));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), 
           .D(n10296));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_adj_991 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n17507));   // coms.v(517[9:65])
    defparam i1_2_lut_3_lut_adj_991.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut_adj_992 (.I0(n16468), .I1(n1396), .I2(\data_in[1]_c [0]), 
            .I3(\data_in_frame[1] [0]), .O(n10232));
    defparam i1_4_lut_4_lut_adj_992.LUT_INIT = 16'h3210;
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), 
           .D(n10299));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_993 (.I0(byte_transmit_counter2[0]), .I1(byte_transmit_counter2[1]), 
            .I2(GND_net), .I3(GND_net), .O(n134));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'heeee;
    SB_DFF data_in_0___i131 (.Q(\data_in[16] [2]), .C(CLK_c), .D(n10454));   // coms.v(402[9] 410[5])
    SB_LUT4 i2_3_lut_4_lut_adj_994 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[0] [1]), .I3(n17553), .O(n8658));   // coms.v(452[9:67])
    defparam i2_3_lut_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i7892_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][5] ), 
            .I3(\data_in_frame[3] [5]), .O(n10308));
    defparam i7892_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_3_lut_adj_995 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n9163));   // coms.v(452[9:67])
    defparam i1_2_lut_3_lut_adj_995.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_996 (.I0(n9058), .I1(\data_in_frame[4] [3]), 
            .I2(\data_in_frame[8] [3]), .I3(\data_in_frame[7] [7]), .O(n8725));   // coms.v(230[15:344])
    defparam i1_2_lut_3_lut_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut (.I0(n18603), .I1(\data_out_frame2[20] [0]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2510));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\data_out[8] [7]), .I1(\data_out[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17454));   // coms.v(21[11:19])
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i130 (.Q(\data_in[16] [1]), .C(CLK_c), .D(n10453));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i129 (.Q(\data_in[16] [0]), .C(CLK_c), .D(n10452));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i128 (.Q(\data_in[15] [7]), .C(CLK_c), .D(n10451));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i73 (.Q(\data_in[9] [0]), .C(CLK_c), .D(n10396));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut (.I0(n18435), .I1(n22_adj_2510), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[0]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7813_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[0] [7]), 
            .I3(\data_in_frame[0] [7]), .O(n10229));
    defparam i7813_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_3_lut_adj_998 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n17602));   // coms.v(517[9:65])
    defparam i1_2_lut_3_lut_adj_998.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_999 (.I0(\data_out[5] [2]), .I1(data_out_6__3__N_788), 
            .I2(\data_out[5] [1]), .I3(n17415), .O(n17659));   // coms.v(114[16:245])
    defparam i1_2_lut_3_lut_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\data_out[7] [2]), .I1(n17492), .I2(n17454), 
            .I3(n17635), .O(data_out_10__3__N_163));   // coms.v(174[15:122])
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [0]), .I2(\data_out_frame2[15] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18606));
    defparam byte_transmit_counter2_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1001 (.I0(tx_active), .I1(tx_transmit), .I2(tx_transmit_N_2239[3]), 
            .I3(n8550), .O(n113));
    defparam i1_2_lut_4_lut_adj_1001.LUT_INIT = 16'h1110;
    SB_LUT4 i7810_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[0][6] ), 
            .I3(\data_in_frame[0] [6]), .O(n10226));
    defparam i7810_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i2_3_lut_4_lut_adj_1002 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[4] [3]), 
            .I2(n9058), .I3(n9254), .O(n17522));   // coms.v(70[15:74])
    defparam i2_3_lut_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(data_out_7__7__N_519), .I1(\data_out[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17665));   // coms.v(116[16:91])
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i3 (.Q(\data_in[0][2] ), .C(CLK_c), .D(n9937));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_4_lut_4_lut_adj_1004 (.I0(n16468), .I1(n1396), .I2(\data_in[0][5] ), 
            .I3(\data_in_frame[0] [5]), .O(n10222));
    defparam i1_4_lut_4_lut_adj_1004.LUT_INIT = 16'h3210;
    SB_LUT4 i2_3_lut_4_lut_adj_1005 (.I0(n119), .I1(tx_active), .I2(tx_transmit), 
            .I3(n29), .O(\UART_TRANSMITTER.state_7__N_1749[2] ));   // coms.v(329[6] 341[9])
    defparam i2_3_lut_4_lut_adj_1005.LUT_INIT = 16'h0002;
    SB_LUT4 i7803_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[0][4] ), 
            .I3(\data_in_frame[0] [4]), .O(n10219));
    defparam i7803_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_DFF data_in_0___i4 (.Q(\data_in[0]_c [3]), .C(CLK_c), .D(n9936));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i5 (.Q(\data_in[0][4] ), .C(CLK_c), .D(n9935));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i6 (.Q(\data_in[0][5] ), .C(CLK_c), .D(n9934));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i7 (.Q(\data_in[0][6] ), .C(CLK_c), .D(n9932));   // coms.v(402[9] 410[5])
    SB_LUT4 i3_3_lut (.I0(n17668), .I1(n8812), .I2(n9195), .I3(GND_net), 
            .O(n8_adj_2511));   // coms.v(116[16:91])
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(n17623), .I1(n8926), .I2(n8_adj_2511), 
            .I3(n17665), .O(data_out_10__0__N_259));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1007 (.I0(n119), .I1(n13415), .I2(n29), 
            .I3(n8486), .O(n8488));   // coms.v(277[4] 373[11])
    defparam i1_2_lut_4_lut_adj_1007.LUT_INIT = 16'hfd00;
    SB_LUT4 i1_4_lut_4_lut_adj_1008 (.I0(n16468), .I1(n1396), .I2(\data_in[0]_c [3]), 
            .I3(\data_in_frame[0] [3]), .O(n10216));
    defparam i1_4_lut_4_lut_adj_1008.LUT_INIT = 16'h3210;
    SB_LUT4 n18606_bdd_4_lut (.I0(n18606), .I1(\data_out_frame2[13] [0]), 
            .I2(\data_out_frame2[12] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n17779));
    defparam n18606_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut (.I0(\data_out_frame2[8] [4]), 
            .I1(\data_out_frame2[9] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n8_c));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut (.I0(\data_out_frame2[10] [4]), 
            .I1(\data_out_frame2[11] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n9));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7797_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[0][2] ), 
            .I3(\data_in_frame[0] [2]), .O(n10213));
    defparam i7797_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i2_2_lut_3_lut_adj_1009 (.I0(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I1(n63), .I2(n63_adj_9), .I3(GND_net), .O(n16468));
    defparam i2_2_lut_3_lut_adj_1009.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16110 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [0]), .I2(\data_out_frame2[19][0] ), 
            .I3(byte_transmit_counter2[1]), .O(n18600));
    defparam byte_transmit_counter2_0__bdd_4_lut_16110.LUT_INIT = 16'he4aa;
    SB_LUT4 i9_4_lut_adj_1010 (.I0(n17_adj_2486), .I1(\data_in[0]_c [3]), 
            .I2(n16_adj_2485), .I3(n17745), .O(n63));   // coms.v(435[16:89])
    defparam i9_4_lut_adj_1010.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(n63), .I1(n63_adj_9), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2512));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1012 (.I0(\data_in[3][2] ), .I1(\data_in[2][3] ), 
            .I2(\data_in[0][5] ), .I3(\data_in[1][4] ), .O(n16_adj_2513));
    defparam i6_4_lut_adj_1012.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1013 (.I0(n8559), .I1(\data_in[3] [4]), .I2(n8556), 
            .I3(n8572), .O(n17_adj_2514));
    defparam i7_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 i7794_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[0][1] ), 
            .I3(\data_in_frame[0] [1]), .O(n10210));
    defparam i7794_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 n18600_bdd_4_lut (.I0(n18600), .I1(\data_out_frame2[17] [0]), 
            .I2(\data_out_frame2[16] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n18603));
    defparam n18600_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1014 (.I0(n17_adj_2514), .I1(\data_in[3] [0]), 
            .I2(n16_adj_2513), .I3(\data_in[0][6] ), .O(\FRAME_MATCHER.next_state_31__N_2026[1] ));
    defparam i9_4_lut_adj_1014.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_4_lut_adj_1015 (.I0(\data_in_frame[5] [5]), .I1(n25_adj_2491), 
            .I2(n9186), .I3(n22_adj_2508), .O(n8857));   // coms.v(452[9:67])
    defparam i1_2_lut_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i3947_3_lut (.I0(\data_in_frame[6] [0]), .I1(\data_in[6][0] ), 
            .I2(n16468), .I3(GND_net), .O(n2599));   // coms.v(435[13] 445[7])
    defparam i3947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15818_3_lut (.I0(\data_out_frame2[0] [6]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n18078));
    defparam i15818_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i3949_3_lut_4_lut (.I0(\data_in_frame[5] [7]), .I1(\data_in[5] [7]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2600));   // coms.v(435[13] 445[7])
    defparam i3949_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_4_lut_4_lut_adj_1016 (.I0(n16468), .I1(n1396), .I2(\data_in[0]_c [0]), 
            .I3(\data_in_frame[0] [0]), .O(n10188));
    defparam i1_4_lut_4_lut_adj_1016.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16105 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [7]), .I2(\data_out_frame2[11] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18588));
    defparam byte_transmit_counter2_0__bdd_4_lut_16105.LUT_INIT = 16'he4aa;
    SB_LUT4 i13613_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3] [4]), 
            .I3(\data_in_frame[3] [4]), .O(n10305));
    defparam i13613_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame2[6] [6]), 
            .I1(\data_out_frame2[7] [6]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2515));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(\FRAME_MATCHER.state [1]), .I1(n9606), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n81), .O(n1396));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hccce;
    SB_LUT4 i3951_3_lut_4_lut (.I0(\data_in_frame[5] [6]), .I1(\data_in[5] [6]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2601));   // coms.v(435[13] 445[7])
    defparam i3951_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n18588_bdd_4_lut (.I0(n18588), .I1(\data_out_frame2[9] [7]), 
            .I2(\data_out_frame2[8] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n17785));
    defparam n18588_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15843_2_lut (.I0(\data_out[10] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18016));   // coms.v(243[28:49])
    defparam i15843_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3959_3_lut_4_lut (.I0(\data_in_frame[5] [2]), .I1(\data_in[5] [2]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2605));   // coms.v(435[13] 445[7])
    defparam i3959_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut (.I0(\data_out_frame2[5] [6]), 
            .I1(n5_adj_2515), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2506));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i8206_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4][7] ), 
            .I3(\data_in_frame[4] [7]), .O(n10622));
    defparam i8206_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[5] [4]), .I1(n8674), .I2(GND_net), 
            .I3(GND_net), .O(n8062));   // coms.v(117[16:83])
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i15292_2_lut (.I0(\UART_TRANSMITTER.state[1] ), .I1(n149), .I2(GND_net), 
            .I3(GND_net), .O(n17741));   // coms.v(271[13:18])
    defparam i15292_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i8_3_lut (.I0(\data_out[8] [0]), 
            .I1(\data_out[9] [0]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2516));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1019 (.I0(n13415), .I1(n8550), .I2(n17741), .I3(tx_transmit_N_2239[3]), 
            .O(n93));   // coms.v(271[13:18])
    defparam i1_4_lut_adj_1019.LUT_INIT = 16'h5444;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16096 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [7]), .I2(\data_out_frame2[15] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18582));
    defparam byte_transmit_counter2_0__bdd_4_lut_16096.LUT_INIT = 16'he4aa;
    SB_LUT4 i15806_4_lut (.I0(n8_adj_2516), .I1(\byte_transmit_counter[2] ), 
            .I2(n18016), .I3(byte_transmit_counter[1]), .O(n18015));   // coms.v(243[28:49])
    defparam i15806_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i43_4_lut (.I0(n96), .I1(n93), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(\UART_TRANSMITTER.state[1] ), .O(n25_adj_2517));
    defparam i43_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 n18582_bdd_4_lut (.I0(n18582), .I1(\data_out_frame2[13] [7]), 
            .I2(\data_out_frame2[12] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n17788));
    defparam n18582_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11225_4_lut (.I0(n18501), .I1(\byte_transmit_counter[4] ), 
            .I2(n18015), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[0]));   // coms.v(243[28:49])
    defparam i11225_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i2_3_lut_adj_1020 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n9254));   // coms.v(70[15:74])
    defparam i2_3_lut_adj_1020.LUT_INIT = 16'h9696;
    SB_LUT4 i3957_3_lut_4_lut (.I0(\data_in_frame[5] [3]), .I1(\data_in[5] [3]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2604));   // coms.v(435[13] 445[7])
    defparam i3957_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_3_lut_adj_1021 (.I0(n9631), .I1(n25_adj_2517), .I2(\UART_TRANSMITTER.state[0] ), 
            .I3(GND_net), .O(n1314));
    defparam i1_3_lut_adj_1021.LUT_INIT = 16'h5d5d;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16091 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [7]), .I2(\data_out_frame2[19] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18576));
    defparam byte_transmit_counter2_0__bdd_4_lut_16091.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_4_lut_adj_1022 (.I0(n16468), .I1(n1396), .I2(\data_in[4]_c [6]), 
            .I3(\data_in_frame[4] [6]), .O(n10619));
    defparam i1_4_lut_4_lut_adj_1022.LUT_INIT = 16'h3210;
    SB_LUT4 i3955_3_lut_4_lut (.I0(\data_in_frame[5] [4]), .I1(\data_in[5] [4]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2603));   // coms.v(435[13] 445[7])
    defparam i3955_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n18360_bdd_4_lut (.I0(n18360), .I1(n6_adj_2504), .I2(n18086), 
            .I3(byte_transmit_counter2[3]), .O(n18363));
    defparam n18360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3961_3_lut_4_lut (.I0(\data_in_frame[5] [1]), .I1(\data_in[5] [1]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2606));   // coms.v(435[13] 445[7])
    defparam i3961_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i59_3_lut (.I0(\data_out[6] [1]), .I1(\data_out[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n45_adj_2518));   // coms.v(19[11:32])
    defparam i59_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n18576_bdd_4_lut (.I0(n18576), .I1(\data_out_frame2[17] [7]), 
            .I2(\data_out_frame2[16] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18579));
    defparam n18576_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8198_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4][5] ), 
            .I3(\data_in_frame[4] [5]), .O(n10614));
    defparam i8198_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i8195_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4]_c [4]), 
            .I3(\data_in_frame[4] [4]), .O(n10611));
    defparam i8195_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_4_lut_4_lut_adj_1023 (.I0(n16468), .I1(n1396), .I2(\data_in[4] [1]), 
            .I3(\data_in_frame[4] [1]), .O(n10608));
    defparam i1_4_lut_4_lut_adj_1023.LUT_INIT = 16'h3210;
    SB_LUT4 i15803_2_lut (.I0(\data_out[10] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18073));   // coms.v(243[28:49])
    defparam i15803_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i8_3_lut (.I0(\data_out[8] [1]), 
            .I1(\data_out[9] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2519));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_1_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut (.I0(n18579), .I1(\data_out_frame2[20] [7]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2520));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut (.I0(n18423), .I1(n22_adj_2520), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[7]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7934_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4][2] ), 
            .I3(\data_in_frame[4] [2]), .O(n10350));
    defparam i7934_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut (.I0(n18555), .I1(\data_out_frame2[20] [6]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2521));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i60_4_lut (.I0(\data_out[5] [1]), .I1(n45_adj_2518), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n46));   // coms.v(19[11:32])
    defparam i60_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut (.I0(n18411), .I1(n22_adj_2521), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[6]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7940_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4][3] ), 
            .I3(\data_in_frame[4] [3]), .O(n10356));
    defparam i7940_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9176));   // coms.v(70[15:74])
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut (.I0(n96), .I1(n113), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n17709));
    defparam i13_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i13941_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[4][0] ), 
            .I3(\data_in_frame[4] [0]), .O(n10663));
    defparam i13941_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16086 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [0]), .I2(\data_out_frame2[11] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18570));
    defparam byte_transmit_counter2_0__bdd_4_lut_16086.LUT_INIT = 16'he4aa;
    SB_LUT4 n18570_bdd_4_lut (.I0(n18570), .I1(\data_out_frame2[9] [0]), 
            .I2(\data_out_frame2[8] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n17773));
    defparam n18570_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i1_3_lut (.I0(\data_out[0][1] ), 
            .I1(\data_out[1] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n1_adj_2522));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i127 (.Q(\data_in[15] [6]), .C(CLK_c), .D(n10450));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15935 (.I0(byte_transmit_counter[1]), 
            .I1(n17936), .I2(n5_adj_2499), .I3(\byte_transmit_counter[2] ), 
            .O(n18378));
    defparam byte_transmit_counter_1__bdd_4_lut_15935.LUT_INIT = 16'he4aa;
    SB_LUT4 i13950_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][7] ), 
            .I3(\data_in_frame[3] [7]), .O(n10314));
    defparam i13950_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n13415), .I1(n8550), .I2(n97), .I3(tx_transmit_N_2239[3]), 
            .O(n96));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'h5554;
    SB_LUT4 i3945_3_lut (.I0(\data_in_frame[6] [1]), .I1(\data_in[6]_c [1]), 
            .I2(n16468), .I3(GND_net), .O(n2598));   // coms.v(435[13] 445[7])
    defparam i3945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15828_4_lut (.I0(n8_adj_2519), .I1(\byte_transmit_counter[2] ), 
            .I2(n18073), .I3(byte_transmit_counter[1]), .O(n18014));   // coms.v(19[11:32])
    defparam i15828_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 n18384_bdd_4_lut (.I0(n18384), .I1(n6_adj_2496), .I2(n18080), 
            .I3(byte_transmit_counter2[3]), .O(n18387));
    defparam n18384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7880_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][2] ), 
            .I3(\data_in_frame[3] [2]), .O(n10296));
    defparam i7880_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16081 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [6]), .I2(\data_out_frame2[11] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18564));
    defparam byte_transmit_counter2_0__bdd_4_lut_16081.LUT_INIT = 16'he4aa;
    SB_LUT4 i3963_3_lut_4_lut (.I0(\data_in_frame[5] [0]), .I1(\data_in[5] [0]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2607));   // coms.v(435[13] 445[7])
    defparam i3963_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i13947_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2]_c [0]), 
            .I3(\data_in_frame[2] [0]), .O(n10262));
    defparam i13947_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i7850_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2][1] ), 
            .I3(\data_in_frame[2] [1]), .O(n10266));
    defparam i7850_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_DFF data_in_0___i126 (.Q(\data_in[15] [5]), .C(CLK_c), .D(n10449));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i72 (.Q(\data_in[8] [7]), .C(CLK_c), .D(n10395));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17553));   // coms.v(452[9:67])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut (.I0(n18537), .I1(\data_out_frame2[20] [5]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2523));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut (.I0(n18387), .I1(n22_adj_2523), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[5]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i4518_2_lut (.I0(n29), .I1(n113), .I2(GND_net), .I3(GND_net), 
            .O(n6878));   // coms.v(362[16] 370[10])
    defparam i4518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i58_4_lut (.I0(n1_adj_2522), .I1(n46), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[1]), .O(n44_adj_2524));   // coms.v(19[11:32])
    defparam i58_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i7853_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2] [2]), 
            .I3(\data_in_frame[2] [2]), .O(n10269));
    defparam i7853_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i7856_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2][3] ), 
            .I3(\data_in_frame[2] [3]), .O(n10272));
    defparam i7856_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 n18564_bdd_4_lut (.I0(n18564), .I1(\data_out_frame2[9] [6]), 
            .I2(\data_out_frame2[8] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n17794));
    defparam n18564_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_1027 (.I0(\UART_TRANSMITTER.state[1] ), .I1(n4430), 
            .I2(n17709), .I3(n8488), .O(n16485));
    defparam i2_4_lut_adj_1027.LUT_INIT = 16'hffce;
    SB_LUT4 i7860_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2] [4]), 
            .I3(\data_in_frame[2] [4]), .O(n10276));
    defparam i7860_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i7863_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2][5] ), 
            .I3(\data_in_frame[2] [5]), .O(n10279));
    defparam i7863_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut (.I0(n18531), .I1(\data_out_frame2[20] [4]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2525));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_4_lut_adj_1028 (.I0(n16468), .I1(n1396), .I2(\data_in[2][6] ), 
            .I3(\data_in_frame[2] [6]), .O(n10333));
    defparam i1_4_lut_4_lut_adj_1028.LUT_INIT = 16'h3210;
    SB_LUT4 i11600217_i1_3_lut (.I0(n18459), .I1(n18447), .I2(byte_transmit_counter2[3]), 
            .I3(GND_net), .O(n15));
    defparam i11600217_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(\byte_transmit_counter[4] ), .I1(n44_adj_2524), 
            .I2(n18014), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[1]));   // coms.v(19[11:32])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'h5044;
    SB_LUT4 i7870_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[2][7] ), 
            .I3(\data_in_frame[2] [7]), .O(n10286));
    defparam i7870_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(\UART_TRANSMITTER.state[1] ), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(n17364), .I3(n6878), .O(n17672));
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'h57df;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17632));   // coms.v(452[9:67])
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut (.I0(n15), .I1(n22_adj_2525), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[4]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7883_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][3] ), 
            .I3(\data_in_frame[3] [3]), .O(n10299));
    defparam i7883_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 i13944_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3] [0]), 
            .I3(\data_in_frame[3] [0]), .O(n10289));
    defparam i13944_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16076 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [6]), .I2(\data_out_frame2[15] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18558));
    defparam byte_transmit_counter2_0__bdd_4_lut_16076.LUT_INIT = 16'he4aa;
    SB_LUT4 i7877_4_lut_4_lut (.I0(n16468), .I1(n1396), .I2(\data_in[3][1] ), 
            .I3(\data_in_frame[3] [1]), .O(n10293));
    defparam i7877_4_lut_4_lut.LUT_INIT = 16'h3210;
    SB_LUT4 n18558_bdd_4_lut (.I0(n18558), .I1(\data_out_frame2[13] [6]), 
            .I2(\data_out_frame2[12] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n17797));
    defparam n18558_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15800_2_lut (.I0(\data_out[10] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18071));   // coms.v(243[28:49])
    defparam i15800_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i8_3_lut (.I0(\data_out[8] [2]), 
            .I1(\data_out[9] [2]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2526));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i125 (.Q(\data_in[15] [4]), .C(CLK_c), .D(n10448));   // coms.v(402[9] 410[5])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut (.I0(n18513), .I1(\data_out_frame2[20] [3]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2527));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16071 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [6]), .I2(\data_out_frame2[19] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18552));
    defparam byte_transmit_counter2_0__bdd_4_lut_16071.LUT_INIT = 16'he4aa;
    SB_LUT4 n18552_bdd_4_lut (.I0(n18552), .I1(\data_out_frame2[17] [6]), 
            .I2(\data_out_frame2[16] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18555));
    defparam n18552_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3953_3_lut_4_lut (.I0(\data_in_frame[5] [5]), .I1(\data_in[5] [5]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2602));   // coms.v(435[13] 445[7])
    defparam i3953_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16066 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [5]), .I2(\data_out_frame2[11] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18546));
    defparam byte_transmit_counter2_0__bdd_4_lut_16066.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut (.I0(n18375), .I1(n22_adj_2527), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[3]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n18546_bdd_4_lut (.I0(n18546), .I1(\data_out_frame2[9] [5]), 
            .I2(\data_out_frame2[8] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n17803));
    defparam n18546_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1032 (.I0(data_out_7__7__N_519), .I1(\data_out[7] [5]), 
            .I2(\data_out[7] [6]), .I3(GND_net), .O(n17492));   // coms.v(168[15:28])
    defparam i1_2_lut_3_lut_adj_1032.LUT_INIT = 16'h9696;
    SB_LUT4 i15802_4_lut (.I0(n8_adj_2526), .I1(\byte_transmit_counter[2] ), 
            .I2(n18071), .I3(byte_transmit_counter[1]), .O(n18072));   // coms.v(243[28:49])
    defparam i15802_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11425_4_lut (.I0(n18381), .I1(\byte_transmit_counter[4] ), 
            .I2(n18072), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[2]));   // coms.v(243[28:49])
    defparam i11425_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1033 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[4] [0]), .O(n25_adj_2491));   // coms.v(383[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(data_out_7__7__N_519), .I1(\data_out[7] [5]), 
            .I2(n9087), .I3(n17668), .O(n8_adj_2528));   // coms.v(168[15:28])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16061 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [5]), .I2(\data_out_frame2[15] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18540));
    defparam byte_transmit_counter2_0__bdd_4_lut_16061.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut (.I0(n18489), .I1(\data_out_frame2[20] [2]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2529));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n18540_bdd_4_lut (.I0(n18540), .I1(\data_out_frame2[13] [5]), 
            .I2(\data_out_frame2[12] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n17806));
    defparam n18540_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9328));   // coms.v(517[9:65])
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut (.I0(n18369), .I1(n22_adj_2529), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[2]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16056 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [5]), .I2(\data_out_frame2[19] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n18534));
    defparam byte_transmit_counter2_0__bdd_4_lut_16056.LUT_INIT = 16'he4aa;
    SB_LUT4 n18534_bdd_4_lut (.I0(n18534), .I1(\data_out_frame2[17] [5]), 
            .I2(\data_out_frame2[16] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n18537));
    defparam n18534_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut (.I0(\data_out_frame2[14] [4]), 
            .I1(\data_out_frame2[15] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n12_c));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1035 (.I0(n9328), .I1(n17403), .I2(n30_adj_2489), 
            .I3(n17602), .O(n9345));   // coms.v(517[9:65])
    defparam i3_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15940 (.I0(byte_transmit_counter[1]), 
            .I1(n17937), .I2(n5_adj_2490), .I3(\byte_transmit_counter[2] ), 
            .O(n18390));
    defparam byte_transmit_counter_1__bdd_4_lut_15940.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut (.I0(\data_out_frame2[12] [4]), 
            .I1(\data_out_frame2[13] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n11));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16051 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [4]), .I2(\data_out_frame2[19] [4]), 
            .I3(byte_transmit_counter2[1]), .O(n18528));
    defparam byte_transmit_counter2_0__bdd_4_lut_16051.LUT_INIT = 16'he4aa;
    SB_LUT4 n18528_bdd_4_lut (.I0(n18528), .I1(\data_out_frame2[17] [4]), 
            .I2(\data_out_frame2[16] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n18531));
    defparam n18528_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15797_2_lut (.I0(\data_out[10] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18069));   // coms.v(243[28:49])
    defparam i15797_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut (.I0(n18471), .I1(\data_out_frame2[20] [1]), 
            .I2(byte_transmit_counter2[2]), .I3(n134), .O(n22_adj_2530));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16046 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [3]), .I2(\data_out_frame2[11] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18522));
    defparam byte_transmit_counter2_0__bdd_4_lut_16046.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut (.I0(n18363), .I1(n22_adj_2530), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[1]));   // coms.v(417[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i8_3_lut (.I0(\data_out[8] [3]), 
            .I1(\data_out[9] [3]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2531));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15799_4_lut (.I0(n8_adj_2531), .I1(\byte_transmit_counter[2] ), 
            .I2(n18069), .I3(byte_transmit_counter[1]), .O(n18070));   // coms.v(243[28:49])
    defparam i15799_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_2_lut_3_lut_adj_1036 (.I0(n9058), .I1(\data_in_frame[4] [3]), 
            .I2(n17467), .I3(GND_net), .O(n8751));   // coms.v(230[15:344])
    defparam i1_2_lut_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1037 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_2532));   // coms.v(300[11:30])
    defparam i2_2_lut_adj_1037.LUT_INIT = 16'heeee;
    SB_LUT4 n18522_bdd_4_lut (.I0(n18522), .I1(\data_out_frame2[9] [3]), 
            .I2(\data_out_frame2[8] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n17815));
    defparam n18522_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1038 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n31), .I3(\FRAME_MATCHER.state [0]), .O(n9606));
    defparam i1_3_lut_4_lut_adj_1038.LUT_INIT = 16'h0100;
    SB_LUT4 i11421_4_lut (.I0(n18393), .I1(\byte_transmit_counter[4] ), 
            .I2(n18070), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[3]));   // coms.v(243[28:49])
    defparam i11421_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16041 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [3]), .I2(\data_out_frame2[15] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18516));
    defparam byte_transmit_counter2_0__bdd_4_lut_16041.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1039 (.I0(delay_counter[10]), .I1(delay_counter[9]), 
            .I2(delay_counter[12]), .I3(delay_counter[6]), .O(n14_adj_2533));   // coms.v(300[11:30])
    defparam i6_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1040 (.I0(delay_counter[5]), .I1(n14_adj_2533), 
            .I2(n10_adj_2532), .I3(delay_counter[8]), .O(n17306));   // coms.v(300[11:30])
    defparam i7_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 n18516_bdd_4_lut (.I0(n18516), .I1(\data_out_frame2[13] [3]), 
            .I2(\data_out_frame2[12] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n17818));
    defparam n18516_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(n17306), .I1(n17387), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_2534));   // coms.v(300[11:30])
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1042 (.I0(\delay_counter[14] ), .I1(\delay_counter[0] ), 
            .I2(\delay_counter[13] ), .I3(n6_adj_2534), .O(n29));   // coms.v(300[11:30])
    defparam i4_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16036 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [3]), .I2(\data_out_frame2[19] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n18510));
    defparam byte_transmit_counter2_0__bdd_4_lut_16036.LUT_INIT = 16'he4aa;
    SB_LUT4 n18510_bdd_4_lut (.I0(n18510), .I1(\data_out_frame2[17] [3]), 
            .I2(\data_out_frame2[16] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n18513));
    defparam n18510_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1043 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(n10_adj_2493), .I3(n9039), .O(n17428));   // coms.v(76[16:93])
    defparam i5_3_lut_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i15822_2_lut (.I0(\data_out[10] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18067));   // coms.v(243[28:49])
    defparam i15822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i1_3_lut (.I0(\data_out[0] [6]), 
            .I1(\data_out[1][6] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n1_adj_2484));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15720_2_lut (.I0(\data_out[3][6] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18090));
    defparam i15720_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i8_3_lut (.I0(\data_out[8] [4]), 
            .I1(\data_out[9] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2535));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1044 (.I0(\data_out[7] [5]), .I1(\data_out[7] [4]), 
            .I2(n8953), .I3(GND_net), .O(n17626));   // coms.v(173[15:115])
    defparam i1_2_lut_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i15796_4_lut (.I0(n8_adj_2535), .I1(\byte_transmit_counter[2] ), 
            .I2(n18067), .I3(byte_transmit_counter[1]), .O(n18068));   // coms.v(243[28:49])
    defparam i15796_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i3_4_lut_adj_1045 (.I0(\data_in_frame[5] [4]), .I1(n8658), .I2(n9058), 
            .I3(n9163), .O(n17470));   // coms.v(517[9:65])
    defparam i3_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16031 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [2]), .I2(\data_out_frame2[11] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18504));
    defparam byte_transmit_counter2_0__bdd_4_lut_16031.LUT_INIT = 16'he4aa;
    SB_LUT4 i11416_4_lut (.I0(n18399), .I1(\byte_transmit_counter[4] ), 
            .I2(n18068), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[4]));   // coms.v(243[28:49])
    defparam i11416_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 n18504_bdd_4_lut (.I0(n18504), .I1(\data_out_frame2[9] [2]), 
            .I2(\data_out_frame2[8] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n17824));
    defparam n18504_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1046 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(n17614), .I3(n10_adj_2536), .O(n8666));   // coms.v(76[16:93])
    defparam i5_3_lut_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_2427));   // coms.v(383[12:25])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i15788_2_lut (.I0(\data_out[10] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18064));   // coms.v(243[28:49])
    defparam i15788_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i8_3_lut (.I0(\data_out[8] [5]), 
            .I1(\data_out[9] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2537));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n157));   // coms.v(428[12] 532[6])
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'h2222;
    SB_LUT4 i10637_3_lut (.I0(\data_in[3][6] ), .I1(\data_in[4]_c [6]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10330));   // coms.v(377[7:20])
    defparam i10637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15791_4_lut (.I0(n8_adj_2537), .I1(\byte_transmit_counter[2] ), 
            .I2(n18064), .I3(byte_transmit_counter[1]), .O(n18065));   // coms.v(243[28:49])
    defparam i15791_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11411_4_lut (.I0(n18405), .I1(\byte_transmit_counter[4] ), 
            .I2(n18065), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[5]));   // coms.v(243[28:49])
    defparam i11411_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i9090_3_lut (.I0(\data_in[7]_c [1]), .I1(\data_in[8] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10381));   // coms.v(377[7:20])
    defparam i9090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15746_2_lut (.I0(\data_out[10] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18060));   // coms.v(243[28:49])
    defparam i15746_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10536_3_lut (.I0(\data_out[8] [7]), .I1(\data_out[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n8_adj_2538));   // coms.v(19[11:32])
    defparam i10536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15781_4_lut (.I0(n8_adj_2538), .I1(\byte_transmit_counter[2] ), 
            .I2(n18060), .I3(byte_transmit_counter[1]), .O(n18061));   // coms.v(243[28:49])
    defparam i15781_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11402_4_lut (.I0(n18429), .I1(\byte_transmit_counter[4] ), 
            .I2(n18061), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[7]));   // coms.v(243[28:49])
    defparam i11402_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n17911), .I2(n5_adj_2488), .I3(\byte_transmit_counter[2] ), 
            .O(n18498));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i3935_3_lut_4_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in[6] [6]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2593));   // coms.v(435[13] 445[7])
    defparam i3935_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_adj_1049 (.I0(\data_in_frame[6] [7]), .I1(\data_in[6] [7]), 
            .I2(n16468), .I3(n8695), .O(n8867));   // coms.v(435[13] 445[7])
    defparam i1_2_lut_4_lut_adj_1049.LUT_INIT = 16'h53ac;
    SB_LUT4 i3943_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(\data_in[6][2] ), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2597));   // coms.v(435[13] 445[7])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n18498_bdd_4_lut (.I0(n18498), .I1(n2_adj_2487), .I2(n18088), 
            .I3(\byte_transmit_counter[2] ), .O(n18501));
    defparam n18498_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15782_2_lut (.I0(\data_out[10] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18062));   // coms.v(243[28:49])
    defparam i15782_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15705_2_lut (.I0(\rand_setpoint[24] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17957));   // coms.v(277[4] 373[11])
    defparam i15705_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1103_i1_4_lut (.I0(\data_out[0] [6]), .I1(n17957), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2579[0]));   // coms.v(277[4] 373[11])
    defparam mux_1103_i1_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n17442));   // coms.v(383[12:25])
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i8_3_lut (.I0(\data_out[8] [6]), 
            .I1(\data_out[9] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2539));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15787_4_lut (.I0(n8_adj_2539), .I1(\byte_transmit_counter[2] ), 
            .I2(n18062), .I3(byte_transmit_counter[1]), .O(n18063));   // coms.v(243[28:49])
    defparam i15787_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16026 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [2]), .I2(\data_out_frame2[15] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18492));
    defparam byte_transmit_counter2_0__bdd_4_lut_16026.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1051 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[5] [1]), .I3(GND_net), .O(n8976));   // coms.v(517[9:65])
    defparam i1_2_lut_3_lut_adj_1051.LUT_INIT = 16'h9696;
    SB_LUT4 i11407_4_lut (.I0(n18417), .I1(\byte_transmit_counter[4] ), 
            .I2(n18063), .I3(\byte_transmit_counter[3] ), .O(i_Tx_Byte[6]));   // coms.v(243[28:49])
    defparam i11407_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i15710_2_lut (.I0(\rand_setpoint[25] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17962));   // coms.v(277[4] 373[11])
    defparam i15710_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n18492_bdd_4_lut (.I0(n18492), .I1(\data_out_frame2[13] [2]), 
            .I2(\data_out_frame2[12] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n17827));
    defparam n18492_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16016 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [2]), .I2(\data_out_frame2[19] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n18486));
    defparam byte_transmit_counter2_0__bdd_4_lut_16016.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1052 (.I0(\data_out[5] [2]), .I1(n8634), 
            .I2(\data_out[5] [3]), .I3(n17389), .O(n17600));   // coms.v(114[16:245])
    defparam i2_3_lut_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 n18486_bdd_4_lut (.I0(n18486), .I1(\data_out_frame2[17] [2]), 
            .I2(\data_out_frame2[16] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n18489));
    defparam n18486_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1077_i1_4_lut (.I0(data_out_6__1__N_849), .I1(n17962), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2544[0]));   // coms.v(277[4] 373[11])
    defparam mux_1077_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i1_3_lut_4_lut_adj_1053 (.I0(\data_in_frame[5] [6]), .I1(n8687), 
            .I2(n17533), .I3(n2585), .O(n17));
    defparam i1_3_lut_4_lut_adj_1053.LUT_INIT = 16'hf6f9;
    SB_LUT4 i15712_2_lut (.I0(\rand_setpoint[26] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17964));   // coms.v(277[4] 373[11])
    defparam i15712_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16011 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [1]), .I2(\data_out_frame2[11] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18480));
    defparam byte_transmit_counter2_0__bdd_4_lut_16011.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1051_i1_4_lut (.I0(data_out_6__2__N_803), .I1(n17964), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2509[0]));   // coms.v(277[4] 373[11])
    defparam mux_1051_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1054 (.I0(\data_out[8] [5]), .I1(\data_out[8] [4]), 
            .I2(\data_out[6] [6]), .I3(n8953), .O(n8922));   // coms.v(181[16:29])
    defparam i1_2_lut_3_lut_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i15714_2_lut (.I0(\rand_setpoint[27] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17966));   // coms.v(277[4] 373[11])
    defparam i15714_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1055 (.I0(\UART_TRANSMITTER.state[0] ), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n8486));   // coms.v(277[4] 373[11])
    defparam i1_2_lut_3_lut_adj_1055.LUT_INIT = 16'h0404;
    SB_DFF data_in_0___i124 (.Q(\data_in[15] [3]), .C(CLK_c), .D(n10447));   // coms.v(402[9] 410[5])
    SB_LUT4 i3939_3_lut_4_lut (.I0(\data_in_frame[6] [4]), .I1(\data_in[6]_c [4]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2595));   // coms.v(435[13] 445[7])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n18480_bdd_4_lut (.I0(n18480), .I1(\data_out_frame2[9] [1]), 
            .I2(\data_out_frame2[8] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n17833));
    defparam n18480_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1025_i1_4_lut (.I0(data_out_5__3__N_964), .I1(n17966), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2474[0]));   // coms.v(277[4] 373[11])
    defparam mux_1025_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_DFF data_in_0___i123 (.Q(\data_in[15] [2]), .C(CLK_c), .D(n10446));   // coms.v(402[9] 410[5])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1056 (.I0(\data_out[5] [2]), .I1(data_out_5__5__N_950), 
            .I2(data_out_6__3__N_788), .I3(\data_out[5] [1]), .O(data_out_6__5__N_752));   // coms.v(113[16:37])
    defparam i1_2_lut_3_lut_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i15713_4_lut (.I0(data_out_6__2__N_804), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(data_out_5__4__N_959), .I3(\data_out[1][2] ), .O(n17967));   // coms.v(277[4] 373[11])
    defparam i15713_4_lut.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_2_lut_4_lut_adj_1057 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[1] [2]), .I3(n9306), .O(n9054));   // coms.v(71[16:29])
    defparam i1_2_lut_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1058 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [2]), 
            .I2(n17575), .I3(GND_net), .O(n9103));   // coms.v(452[9:67])
    defparam i1_2_lut_3_lut_adj_1058.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_2272_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[7]), .I3(n16411), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_2272_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[6]), .I3(n16410), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_16006 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [1]), .I2(\data_out_frame2[15] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n18474));
    defparam byte_transmit_counter2_0__bdd_4_lut_16006.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1059 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[3] [6]), .O(n10_adj_2536));   // coms.v(128[17:38])
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 mux_999_i1_4_lut (.I0(n17967), .I1(\rand_setpoint[28] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2439[0]));   // coms.v(277[4] 373[11])
    defparam mux_999_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY byte_transmit_counter2_2272_add_4_8 (.CI(n16410), .I0(GND_net), 
            .I1(byte_transmit_counter2[6]), .CO(n16411));
    SB_LUT4 byte_transmit_counter2_2272_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[5]), .I3(n16409), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5065_3_lut_4_lut (.I0(n17364), .I1(n29), .I2(n113), .I3(\UART_TRANSMITTER.state[2] ), 
            .O(n7428));   // coms.v(277[4] 373[11])
    defparam i5065_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 i15717_2_lut (.I0(\rand_setpoint[29] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17970));   // coms.v(277[4] 373[11])
    defparam i15717_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1207_i1_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n2719[0]));   // coms.v(277[4] 373[11])
    defparam mux_1207_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3777_5 (.CI(n16307), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n16308));
    SB_LUT4 i7604_2_lut_4_lut (.I0(\data_in_frame[6] [7]), .I1(\data_in[6] [7]), 
            .I2(n16468), .I3(n1396), .O(n10020));   // coms.v(435[13] 445[7])
    defparam i7604_2_lut_4_lut.LUT_INIT = 16'h00ac;
    SB_LUT4 i9041_3_lut (.I0(\data_in[1]_c [0]), .I1(\data_in[2]_c [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n10342));   // coms.v(377[7:20])
    defparam i9041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1060 (.I0(data_out_5__4__N_959), .I1(data_out_6__2__N_804), 
            .I2(n8634), .I3(\data_out[1][2] ), .O(n17398));   // coms.v(125[17:62])
    defparam i2_3_lut_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i3919_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7][6] ), .I3(\data_in_frame[7] [6]), .O(n2585));   // coms.v(435[13] 445[7])
    defparam i3919_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY byte_transmit_counter2_2272_add_4_7 (.CI(n16409), .I0(GND_net), 
            .I1(byte_transmit_counter2[5]), .CO(n16410));
    SB_LUT4 i3921_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7][5] ), .I3(\data_in_frame[7] [5]), .O(n2586));   // coms.v(435[13] 445[7])
    defparam i3921_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_973_i1_4_lut (.I0(data_out_5__5__N_950), .I1(n17970), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2404[0]));   // coms.v(277[4] 373[11])
    defparam mux_973_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 byte_transmit_counter2_2272_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[4]), .I3(n16408), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15722_2_lut (.I0(\rand_setpoint[30] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17972));   // coms.v(277[4] 373[11])
    defparam i15722_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3925_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7] [3]), .I3(\data_in_frame[7] [3]), .O(n2588));   // coms.v(435[13] 445[7])
    defparam i3925_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\data_out[8] [4]), .I1(\data_out[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n8970));   // coms.v(181[16:29])
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 mux_947_i1_4_lut (.I0(n17389), .I1(n17972), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2369[0]));   // coms.v(277[4] 373[11])
    defparam mux_947_i1_4_lut.LUT_INIT = 16'hcfc5;
    SB_CARRY byte_transmit_counter2_2272_add_4_6 (.CI(n16408), .I0(GND_net), 
            .I1(byte_transmit_counter2[4]), .CO(n16409));
    SB_LUT4 i10772_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7][0] ), .I3(\data_in_frame[7][0] ), .O(n2591));   // coms.v(435[13] 445[7])
    defparam i10772_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_1062 (.I0(\data_out[6] [2]), .I1(\data_out[8] [0]), 
            .I2(\data_out[8] [1]), .I3(GND_net), .O(n8953));   // coms.v(173[15:115])
    defparam i2_3_lut_adj_1062.LUT_INIT = 16'h9696;
    SB_LUT4 i3929_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7]_c [1]), .I3(\data_in_frame[7] [1]), .O(n2590));   // coms.v(435[13] 445[7])
    defparam i3929_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3923_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7]_c [4]), .I3(\data_in_frame[7] [4]), .O(n2587));   // coms.v(435[13] 445[7])
    defparam i3923_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3917_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7][7] ), .I3(\data_in_frame[7] [7]), .O(n2584));   // coms.v(435[13] 445[7])
    defparam i3917_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_0___i122 (.Q(\data_in[15] [1]), .C(CLK_c), .D(n10445));   // coms.v(402[9] 410[5])
    SB_LUT4 i15888_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(data_out_10__7__N_114));   // coms.v(310[5:21])
    defparam i15888_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 byte_transmit_counter2_2272_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[3]), .I3(n16407), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i121 (.Q(\data_in[15] [0]), .C(CLK_c), .D(n10444));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i120 (.Q(\data_in[14] [7]), .C(CLK_c), .D(n10443));   // coms.v(402[9] 410[5])
    SB_DFF data_in_0___i119 (.Q(\data_in[14] [6]), .C(CLK_c), .D(n10442));   // coms.v(402[9] 410[5])
    SB_LUT4 i3927_3_lut_4_lut (.I0(n4_adj_2512), .I1(\FRAME_MATCHER.next_state_31__N_2026[1] ), 
            .I2(\data_in[7] [2]), .I3(\data_in_frame[7] [2]), .O(n2589));   // coms.v(435[13] 445[7])
    defparam i3927_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY byte_transmit_counter2_2272_add_4_5 (.CI(n16407), .I0(GND_net), 
            .I1(byte_transmit_counter2[3]), .CO(n16408));
    SB_LUT4 i15723_2_lut (.I0(\rand_setpoint[31] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17974));   // coms.v(277[4] 373[11])
    defparam i15723_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_2272_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[2]), .I3(n16406), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15672_4_lut (.I0(data_out_5__5__N_950), .I1(n17438), .I2(data_out_6__3__N_781), 
            .I3(n17653), .O(n17976));   // coms.v(277[4] 373[11])
    defparam i15672_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1063 (.I0(\data_out[6] [4]), .I1(\data_out[8] [3]), 
            .I2(\data_out[8] [2]), .I3(GND_net), .O(n9091));   // coms.v(175[15:60])
    defparam i2_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(n9091), .I1(n8950), .I2(GND_net), .I3(GND_net), 
            .O(n17566));   // coms.v(175[15:60])
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_out[6] [5]), .I1(\data_out[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17510));   // coms.v(175[15:60])
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i118 (.Q(\data_in[14] [5]), .C(CLK_c), .D(n10441));   // coms.v(402[9] 410[5])
    SB_LUT4 i3_4_lut_adj_1066 (.I0(\data_out[6] [3]), .I1(n17510), .I2(data_out_7__6__N_530), 
            .I3(n17566), .O(n9195));   // coms.v(175[15:60])
    defparam i3_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i117 (.Q(\data_in[14] [4]), .C(CLK_c), .D(n10440));   // coms.v(402[9] 410[5])
    SB_LUT4 mux_921_i1_4_lut (.I0(n17976), .I1(n17974), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2334[0]));   // coms.v(277[4] 373[11])
    defparam mux_921_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_CARRY byte_transmit_counter2_2272_add_4_4 (.CI(n16406), .I0(GND_net), 
            .I1(byte_transmit_counter2[2]), .CO(n16407));
    SB_LUT4 i3_4_lut_adj_1067 (.I0(\data_out[2][0] ), .I1(data_out_6__6__N_729), 
            .I2(\data_out[2] [3]), .I3(n17578), .O(n17653));   // coms.v(76[16:213])
    defparam i3_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_2272_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[1]), .I3(n16405), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1068 (.I0(n17653), .I1(data_out_6__4__N_765), .I2(n17457), 
            .I3(GND_net), .O(n17654));   // coms.v(76[16:213])
    defparam i2_3_lut_adj_1068.LUT_INIT = 16'h9696;
    SB_CARRY byte_transmit_counter2_2272_add_4_3 (.CI(n16405), .I0(GND_net), 
            .I1(byte_transmit_counter2[1]), .CO(n16406));
    SB_LUT4 byte_transmit_counter2_2272_add_4_2_lut (.I0(GND_net), .I1(tx2_transmit_N_2287), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2272_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_884_i1_4_lut (.I0(n17654), .I1(\data_out[0] [6]), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(n8926), .O(n17693));   // coms.v(277[4] 373[11])
    defparam mux_884_i1_4_lut.LUT_INIT = 16'hc5ca;
    SB_CARRY byte_transmit_counter2_2272_add_4_2 (.CI(GND_net), .I0(tx2_transmit_N_2287), 
            .I1(byte_transmit_counter2[0]), .CO(n16405));
    SB_DFF data_in_0___i116 (.Q(\data_in[14] [3]), .C(CLK_c), .D(n10439));   // coms.v(402[9] 410[5])
    SB_LUT4 mux_895_i1_4_lut (.I0(n17693), .I1(\rand_setpoint[16] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2299[0]));   // coms.v(277[4] 373[11])
    defparam mux_895_i1_4_lut.LUT_INIT = 16'hc505;
    SB_LUT4 data_out_6__1__I_638_2_lut (.I0(data_out_6__1__N_850), .I1(data_out_6__7__N_678), 
            .I2(GND_net), .I3(GND_net), .O(data_out_6__1__N_849));   // coms.v(122[16:61])
    defparam data_out_6__1__I_638_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), 
           .D(n10044));   // coms.v(428[12] 532[6])
    SB_LUT4 mux_858_i1_4_lut (.I0(n17415), .I1(data_out_6__1__N_849), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(n8777), .O(n2250[0]));   // coms.v(277[4] 373[11])
    defparam mux_858_i1_4_lut.LUT_INIT = 16'hcac5;
    SB_LUT4 mux_869_i1_4_lut (.I0(n2250[0]), .I1(\rand_setpoint[17] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2264[0]));   // coms.v(277[4] 373[11])
    defparam mux_869_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 data_out_6__2__I_596_2_lut (.I0(data_out_6__2__N_804), .I1(\data_out[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(data_out_6__2__N_803));   // coms.v(123[17:69])
    defparam data_out_6__2__I_596_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_832_i1_4_lut (.I0(n17644), .I1(data_out_6__2__N_803), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(data_out_6__3__N_781), .O(n2215[0]));   // coms.v(277[4] 373[11])
    defparam mux_832_i1_4_lut.LUT_INIT = 16'h353a;
    SB_LUT4 mux_843_i1_4_lut (.I0(n2215[0]), .I1(\rand_setpoint[18] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2229[0]));   // coms.v(277[4] 373[11])
    defparam mux_843_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i3941_3_lut_4_lut (.I0(\data_in_frame[6] [3]), .I1(\data_in[6][3] ), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2596));   // coms.v(435[13] 445[7])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n18378_bdd_4_lut (.I0(n18378), .I1(n2_adj_2483), .I2(n18096), 
            .I3(\byte_transmit_counter[2] ), .O(n18381));
    defparam n18378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(data_out_6__3__N_788), .I1(data_out_5__3__N_964), 
            .I2(GND_net), .I3(GND_net), .O(data_out_6__3__N_785));   // coms.v(124[17:77])
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(data_out_7__4__N_556), .I1(n9195), .I2(GND_net), 
            .I3(GND_net), .O(n17608));   // coms.v(167[15:396])
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 mux_806_i1_4_lut (.I0(n8600), .I1(data_out_6__3__N_785), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(data_out_6__3__N_781), .O(n2180[0]));   // coms.v(277[4] 373[11])
    defparam mux_806_i1_4_lut.LUT_INIT = 16'hc5ca;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n67), .I1(n9606), .I2(n13530), .I3(n19_adj_2540), 
            .O(n4_adj_2480));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'hecee;
    SB_LUT4 i1_2_lut_3_lut_adj_1072 (.I0(\data_out[8] [5]), .I1(data_out_6__3__N_788), 
            .I2(data_out_5__3__N_964), .I3(GND_net), .O(n6_adj_2448));   // coms.v(174[15:122])
    defparam i1_2_lut_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_out[6] [7]), .I1(n8922), .I2(GND_net), 
            .I3(GND_net), .O(n17668));   // coms.v(167[15:396])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 mux_817_i1_4_lut (.I0(n2180[0]), .I1(\rand_setpoint[19] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2194[0]));   // coms.v(277[4] 373[11])
    defparam mux_817_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1074 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[7] [3]), .I3(\data_in_frame[7] [7]), .O(n9204));   // coms.v(226[15:362])
    defparam i1_2_lut_3_lut_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i15875_2_lut_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(n4430), .O(n9518));
    defparam i15875_2_lut_3_lut_4_lut.LUT_INIT = 16'h00e0;
    SB_LUT4 add_3777_16_lut (.I0(n29), .I1(\delay_counter[14] ), .I2(GND_net), 
            .I3(n16318), .O(n18105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1075 (.I0(\data_out[0] [6]), .I1(n9091), 
            .I2(n8950), .I3(GND_net), .O(data_out_9__0__N_475));   // coms.v(175[15:60])
    defparam i1_2_lut_3_lut_adj_1075.LUT_INIT = 16'h6969;
    SB_LUT4 data_out_6__4__I_567_2_lut (.I0(data_out_5__7__N_931), .I1(\data_out[3][6] ), 
            .I2(GND_net), .I3(GND_net), .O(data_out_6__4__N_765));   // coms.v(65[15:44])
    defparam data_out_6__4__I_567_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1076 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[6] [4]), .I3(\data_in_frame[8] [2]), .O(n17629));   // coms.v(226[15:362])
    defparam i1_2_lut_3_lut_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1077 (.I0(data_out_7__6__N_530), .I1(data_out_6__6__N_729), 
            .I2(\data_out[0][5] ), .I3(n17626), .O(data_out_10__6__N_118));   // coms.v(173[15:115])
    defparam i1_2_lut_4_lut_adj_1077.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(n17418), .I1(n17582), .I2(GND_net), 
            .I3(GND_net), .O(n17584));   // coms.v(229[15:344])
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i11502_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n4430));
    defparam i11502_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1079 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[1][1] ), .I3(\data_in_frame[1] [2]), .O(n8874));   // coms.v(452[9:67])
    defparam i1_2_lut_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1080 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[8] [7]), .I3(GND_net), .O(n9380));   // coms.v(230[15:344])
    defparam i1_2_lut_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 add_3777_15_lut (.I0(n29), .I1(\delay_counter[13] ), .I2(GND_net), 
            .I3(n16317), .O(n18008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1081 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[10] [2]), 
            .I2(\data_in_frame[10] [4]), .I3(GND_net), .O(n9051));   // coms.v(232[16:345])
    defparam i1_2_lut_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1082 (.I0(n17608), .I1(n8777), .I2(n8_adj_2528), 
            .I3(n17659), .O(data_out_10__1__N_196));
    defparam i1_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(n9131), .I1(n17544), .I2(GND_net), 
            .I3(GND_net), .O(n17545));   // coms.v(228[15:344])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1084 (.I0(data_out_7__4__N_556), .I1(data_out_7__7__N_519), 
            .I2(data_out_7__6__N_530), .I3(GND_net), .O(n17611));   // coms.v(114[16:245])
    defparam i1_2_lut_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15950 (.I0(byte_transmit_counter2[2]), 
            .I1(n17803), .I2(n17806), .I3(byte_transmit_counter2[3]), 
            .O(n18384));
    defparam byte_transmit_counter2_2__bdd_4_lut_15950.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), 
           .D(n10043));   // coms.v(428[12] 532[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15955 (.I0(byte_transmit_counter[1]), 
            .I1(n17943), .I2(n5_adj_2481), .I3(\byte_transmit_counter[2] ), 
            .O(n18402));
    defparam byte_transmit_counter_1__bdd_4_lut_15955.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), 
           .D(n10039));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_adj_1085 (.I0(n17541), .I1(n8989), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n17543));   // coms.v(227[15:353])
    defparam i2_3_lut_adj_1085.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1086 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n31), .O(n9900));
    defparam i2_3_lut_4_lut_adj_1086.LUT_INIT = 16'h0010;
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), 
           .D(n10038));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), 
           .D(n10034));   // coms.v(428[12] 532[6])
    SB_LUT4 i15860_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n31), .O(n9605));
    defparam i15860_3_lut_4_lut.LUT_INIT = 16'h0414;
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), 
           .D(n10033));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1087 (.I0(n25_adj_2491), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[2] [1]), .I3(n22_adj_2508), .O(n17569));   // coms.v(452[9:67])
    defparam i2_3_lut_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), 
           .D(n10032));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1088 (.I0(\data_out[1][2] ), .I1(\data_out[1] [1]), 
            .I2(data_out_6__1__N_850), .I3(GND_net), .O(data_out_5__3__N_964));   // coms.v(72[16:68])
    defparam i1_2_lut_3_lut_adj_1088.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), 
           .D(n10031));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), 
           .D(n10027));   // coms.v(428[12] 532[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1089 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[1] [5]), 
            .I2(n8645), .I3(n17485), .O(n30_adj_2489));   // coms.v(517[9:65])
    defparam i2_3_lut_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n3203[0]));
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i2_3_lut_4_lut_adj_1090 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[3] [4]), .O(n17516));   // coms.v(517[9:65])
    defparam i2_3_lut_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), 
           .D(n10026));   // coms.v(428[12] 532[6])
    SB_LUT4 mux_780_i1_4_lut (.I0(n17400), .I1(n17398), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(data_out_6__4__N_765), .O(n2145[0]));   // coms.v(277[4] 373[11])
    defparam mux_780_i1_4_lut.LUT_INIT = 16'h353a;
    SB_LUT4 n18402_bdd_4_lut (.I0(n18402), .I1(n2_adj_2476), .I2(n18091), 
            .I3(\byte_transmit_counter[2] ), .O(n18405));
    defparam n18402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_in_frame[9][6] ), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2541));   // coms.v(226[15:362])
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), 
           .D(n10025));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), 
           .D(n10024));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), 
           .D(n10023));   // coms.v(428[12] 532[6])
    SB_LUT4 mux_791_i1_4_lut (.I0(n2145[0]), .I1(\rand_setpoint[20] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2159[0]));   // coms.v(277[4] 373[11])
    defparam mux_791_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6][5] ), .C(CLK_c), 
           .D(n10022));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), 
           .D(n10021));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), 
           .D(n10020));   // coms.v(428[12] 532[6])
    SB_LUT4 i3937_3_lut_4_lut (.I0(\data_in_frame[6][5] ), .I1(\data_in[6] [5]), 
            .I2(\FRAME_MATCHER.next_state_31__N_2026[1] ), .I3(n4_adj_2512), 
            .O(n2594));   // coms.v(435[13] 445[7])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7][0] ), .C(CLK_c), 
           .D(n10019));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), 
           .D(n10018));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), 
           .D(n10017));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), 
           .D(n10016));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), 
           .D(n10009));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1092 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[5] [7]), 
            .I2(n8666), .I3(GND_net), .O(n8061));   // coms.v(116[16:91])
    defparam i1_2_lut_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1093 (.I0(\data_in_frame[5] [0]), .I1(n23_adj_2426), 
            .I2(\data_in_frame[4] [5]), .I3(n9368), .O(n12_adj_2542));   // coms.v(128[17:38])
    defparam i5_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1094 (.I0(n17488), .I1(n17591), .I2(n17504), 
            .I3(n6_adj_2541), .O(n17593));   // coms.v(226[15:362])
    defparam i4_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), 
           .D(n10005));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), 
           .D(n10004));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), 
           .D(n10003));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), 
           .D(n9993));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9028));   // coms.v(229[15:344])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1096 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[10][6] ), 
            .I2(\data_in_frame[7] [2]), .I3(GND_net), .O(n17504));   // coms.v(236[16:315])
    defparam i1_2_lut_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(data_out_5__7__N_931), .I1(\data_out[0][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2543));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1098 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n2839));   // coms.v(71[16:29])
    defparam i1_2_lut_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1099 (.I0(\data_in_frame[7] [2]), .I1(n8061), .I2(n9028), 
            .I3(n9148), .O(n17538));   // coms.v(225[15:370])
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1100 (.I0(byte_transmit_counter2[2]), .I1(byte_transmit_counter2[4]), 
            .I2(byte_transmit_counter2[3]), .I3(GND_net), .O(n18_adj_2544));   // coms.v(413[12:34])
    defparam i1_3_lut_adj_1100.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_754_i1_4_lut (.I0(n4_adj_2543), .I1(data_out_6__5__N_752), 
            .I2(\UART_TRANSMITTER.state[2] ), .I3(\data_out[2] [3]), .O(n9656));   // coms.v(277[4] 373[11])
    defparam mux_754_i1_4_lut.LUT_INIT = 16'hc5ca;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(\data_in_frame[10] [5]), .I1(n8989), 
            .I2(\data_in_frame[10][6] ), .I3(n17538), .O(n17540));   // coms.v(225[15:370])
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), 
           .D(n9989));   // coms.v(428[12] 532[6])
    SB_LUT4 i3_4_lut_adj_1102 (.I0(byte_transmit_counter2[7]), .I1(n18_adj_2544), 
            .I2(byte_transmit_counter2[6]), .I3(byte_transmit_counter2[5]), 
            .O(n19_adj_2540));   // coms.v(413[12:34])
    defparam i3_4_lut_adj_1102.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), 
           .D(n9988));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), 
           .D(n9987));   // coms.v(428[12] 532[6])
    SB_LUT4 i14_2_lut_3_lut_4_lut (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(n9365), .I3(\data_in_frame[3] [0]), .O(n9306));   // coms.v(71[16:29])
    defparam i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15867_2_lut (.I0(n19_adj_2540), .I1(n13530), .I2(GND_net), 
            .I3(GND_net), .O(tx2_transmit_N_2287));
    defparam i15867_2_lut.LUT_INIT = 16'h1111;
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), 
           .D(n9986));   // coms.v(428[12] 532[6])
    SB_CARRY add_3777_15 (.CI(n16317), .I0(\delay_counter[13] ), .I1(GND_net), 
            .CO(n16318));
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), 
           .D(n9985));   // coms.v(428[12] 532[6])
    SB_LUT4 mux_765_i1_4_lut (.I0(n9656), .I1(\rand_setpoint[21] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2124[0]));   // coms.v(277[4] 373[11])
    defparam mux_765_i1_4_lut.LUT_INIT = 16'hc505;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(\data_in_frame[7] [4]), .I1(n9103), .I2(\data_in_frame[7] [1]), 
            .I3(n9279), .O(n17412));   // coms.v(224[15:379])
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1104 (.I0(\data_out[3][4] ), .I1(data_out_5__5__N_950), 
            .I2(data_out_5__4__N_959), .I3(GND_net), .O(n17389));
    defparam i2_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1105 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n67));
    defparam i3_3_lut_adj_1105.LUT_INIT = 16'h1010;
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9][6] ), .C(CLK_c), 
           .D(n9984));   // coms.v(428[12] 532[6])
    SB_LUT4 add_3777_14_lut (.I0(n29), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n16316), .O(n18009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_14_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), 
           .D(n9983));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1106 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [0]), .O(n17403));   // coms.v(71[16:29])
    defparam i1_2_lut_3_lut_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n9982));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n9981));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n9980));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n9979));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n9978));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n9977));   // coms.v(428[12] 532[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10][6] ), .C(CLK_c), 
           .D(n9976));   // coms.v(428[12] 532[6])
    SB_LUT4 i149_2_lut_3_lut (.I0(tx_transmit_N_2239_c[1]), .I1(tx_transmit_N_2239_c[0]), 
            .I2(tx_transmit_N_2239[2]), .I3(GND_net), .O(n149));   // coms.v(25[6:17])
    defparam i149_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i4_4_lut_adj_1107 (.I0(n17412), .I1(n17488), .I2(n17482), 
            .I3(n6_adj_2502), .O(n17490));   // coms.v(226[15:362])
    defparam i4_4_lut_adj_1107.LUT_INIT = 16'h9669;
    SB_LUT4 mux_728_i1_4_lut (.I0(\data_out[0][5] ), .I1(n17600), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(data_out_6__6__N_729), .O(n9658));   // coms.v(277[4] 373[11])
    defparam mux_728_i1_4_lut.LUT_INIT = 16'hc5ca;
    SB_LUT4 mux_739_i1_4_lut (.I0(n9658), .I1(\rand_setpoint[22] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2089[0]));   // coms.v(277[4] 373[11])
    defparam mux_739_i1_4_lut.LUT_INIT = 16'hc505;
    SB_LUT4 i7_4_lut_adj_1108 (.I0(n30_adj_2489), .I1(n8976), .I2(n9279), 
            .I3(n9186), .O(n18_adj_2545));   // coms.v(230[15:344])
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(n17562), .I1(n17629), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_2546));   // coms.v(230[15:344])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1109 (.I0(\data_out[1][6] ), .I1(n8767), .I2(n8926), 
            .I3(GND_net), .O(n17438));   // coms.v(181[16:29])
    defparam i2_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1110 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9][6] ), .I3(\data_in_frame[10] [0]), .O(n9131));   // coms.v(228[15:344])
    defparam i1_2_lut_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1111 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_2542), 
            .I2(\data_in_frame[2] [2]), .I3(n22_adj_2508), .O(n17605));   // coms.v(128[17:38])
    defparam i6_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n9947));   // coms.v(428[12] 532[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1112 (.I0(tx_transmit_N_2239_c[1]), .I1(tx_transmit_N_2239_c[0]), 
            .I2(tx_transmit_N_2239[2]), .I3(GND_net), .O(n97));   // coms.v(25[6:17])
    defparam i1_2_lut_3_lut_adj_1112.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1113 (.I0(\data_in_frame[5] [2]), .I1(n9328), 
            .I2(\data_in_frame[4] [7]), .I3(n8645), .O(n9100));   // coms.v(74[16:53])
    defparam i1_2_lut_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1114 (.I0(data_out_6__3__N_788), .I1(n17438), .I2(n9276), 
            .I3(n6_adj_2467), .O(n17662));   // coms.v(113[16:37])
    defparam i4_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1115 (.I0(n17650), .I1(n18_adj_2545), .I2(n9283), 
            .I3(n8063), .O(n20_adj_2547));   // coms.v(230[15:344])
    defparam i9_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1116 (.I0(n9317), .I1(n20_adj_2547), .I2(n16_adj_2546), 
            .I3(n17470), .O(n8056));   // coms.v(230[15:344])
    defparam i10_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i15747_2_lut (.I0(\data_out[1][7] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18089));
    defparam i15747_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut_adj_1117 (.I0(n8056), .I1(n9240), .I2(n9131), .I3(\data_in_frame[9] [0]), 
            .O(n10_adj_2470));   // coms.v(235[16:323])
    defparam i4_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1118 (.I0(n9204), .I1(n8062), .I2(n2563), 
            .I3(\data_in_frame[7] [2]), .O(n17592));   // coms.v(226[15:362])
    defparam i2_3_lut_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i2_3_lut (.I0(data_out_6__1__N_850), 
            .I1(data_out_5__7__N_931), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2));   // coms.v(243[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2548));   // coms.v(178[16:29])
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 mux_702_i1_4_lut (.I0(data_out_6__7__N_675), .I1(n17611), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(n17662), .O(n2040[0]));   // coms.v(277[4] 373[11])
    defparam mux_702_i1_4_lut.LUT_INIT = 16'h3aca;
    SB_LUT4 i2_4_lut_adj_1120 (.I0(\data_in_frame[5] [7]), .I1(n9043), .I2(n4_adj_2548), 
            .I3(\data_in_frame[6] [3]), .O(n17562));   // coms.v(167[15:498])
    defparam i2_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 mux_713_i1_4_lut (.I0(n2040[0]), .I1(\rand_setpoint[23] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2054[0]));   // coms.v(277[4] 373[11])
    defparam mux_713_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17409));   // coms.v(225[15:370])
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 add_3777_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n16310), .O(n7260[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1122 (.I0(n9043), .I1(n8886), .I2(n15927), 
            .I3(\data_in_frame[7] [2]), .O(n17536));   // coms.v(177[16:29])
    defparam i2_3_lut_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_CARRY add_3777_14 (.CI(n16316), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n16317));
    SB_CARRY add_3777_8 (.CI(n16310), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n16311));
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_out[1][7] ), .I1(n8964), .I2(GND_net), 
            .I3(GND_net), .O(n17578));   // coms.v(62[15:196])
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 add_3777_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n16306), .O(n7260[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(\data_out[0][0] ), .I1(\data_out[0][1] ), 
            .I2(\data_out[0][3] ), .I3(GND_net), .O(n8926));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i61 (.Q(\data_in[7]_c [4]), .C(CLK_c), .D(n10384));   // coms.v(402[9] 410[5])
    SB_LUT4 i5_4_lut_adj_1125 (.I0(n9324), .I1(n9219), .I2(n9345), .I3(\data_in_frame[5] [6]), 
            .O(n12_adj_2549));   // coms.v(167[15:498])
    defparam i5_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 add_3777_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n16315), .O(n7260[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1126 (.I0(\UART_TRANSMITTER.state[0] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n17387), .I3(GND_net), .O(n8529));   // coms.v(277[4] 373[11])
    defparam i1_2_lut_3_lut_adj_1126.LUT_INIT = 16'h0404;
    SB_DFF data_in_0___i32 (.Q(\data_in[3][7] ), .C(CLK_c), .D(n9939));   // coms.v(402[9] 410[5])
    SB_LUT4 i6_4_lut_adj_1127 (.I0(n17562), .I1(n12_adj_2549), .I2(n9208), 
            .I3(\data_in_frame[8] [7]), .O(n17647));   // coms.v(167[15:498])
    defparam i6_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(n9135), .I1(n8989), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_2550));   // coms.v(233[16:338])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_CARRY add_3777_13 (.CI(n16315), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n16316));
    SB_LUT4 i4_4_lut_adj_1129 (.I0(n8995), .I1(n17647), .I2(n17433), .I3(n6_adj_2550), 
            .O(n17649));   // coms.v(233[16:338])
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    uart_tx tx (.r_SM_Main({r_SM_Main}), .CLK_N_keep(CLK_c), .n10638(n10638), 
            .r_Tx_Data({r_Tx_Data}), .r_Clock_Count({r_Clock_Count}), .GND_net(GND_net), 
            .n16998(n16998), .n18103(n18103), .n17366(n17366), .n10637(n10637), 
            .n10636(n10636), .n10635(n10635), .n10634(n10634), .n10633(n10633), 
            .n10632(n10632), .n18102(n18102), .n17054(n17054), .r_Bit_Index({r_Bit_Index}), 
            .n16932(n16932), .VCC_net(VCC_net), .n16954(n16954), .n16968(n16968), 
            .n17078(n17078), .n18101(n18101), .n17028(n17028), .n7364(n7364), 
            .n18104(n18104), .n9972(n9972), .n10702(n10702), .n17084(n17084), 
            .n17082(n17082), .n17080(n17080), .n17030(n17030), .\r_SM_Main_2__N_2323[1] (\r_SM_Main_2__N_2323[1] ), 
            .n18098(n18098), .\r_SM_Main_2__N_2326[0] (tx_transmit), .n4(n4_adj_11), 
            .n8517(n8517), .n12(n12), .n9390(n9390), .n16466(n16466), 
            .n10326(n10326), .n10325(n10325), .n10324(n10324), .tx_active(tx_active), 
            .n10323(n10323), .tx_o(tx_o_adj_8), .n7086(n7086), .n7734(n7734), 
            .tx_enable(tx_enable), .n13601(n13601), .n1(n1), .n3(n3), 
            .n17757(n17757), .n7080(n7080), .n9796(n9796), .n17950(n17950), 
            .n17356(n17356), .n17952(n17952), .n18010(n18010), .n18054(n18054), 
            .n18097(n18097)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1 */ ;   // coms.v(245[10:70])
    uart_tx_U0 tx2 (.n10245(n10245), .VCC_net(VCC_net), .r_Clock_Count({Open_39, 
            Open_40, Open_41, Open_42, Open_43, Open_44, Open_45, 
            Open_46, \r_Clock_Count[0]_adj_12 }), .CLK_c(CLK_c), .r_Bit_Index({r_Bit_Index_adj_35}), 
            .n10625(n10625), .n10346(n10346), .n10008(n10008), .\r_Clock_Count[5] (\r_Clock_Count[5]_adj_16 ), 
            .n10002(n10002), .\r_Clock_Count[4] (\r_Clock_Count[4]_adj_17 ), 
            .n9999(n9999), .\r_Clock_Count[3] (\r_Clock_Count[3]_adj_18 ), 
            .n9996(n9996), .\r_Clock_Count[2] (\r_Clock_Count[2]_adj_19 ), 
            .n9992(n9992), .\r_Clock_Count[1] (\r_Clock_Count[1]_adj_20 ), 
            .tx2_data({tx2_data}), .n10160(n10160), .\r_SM_Main[2] (\r_SM_Main[2]_adj_21 ), 
            .GND_net(GND_net), .n10244(n10244), .n316(n316), .n317(n317), 
            .tx2_o(tx2_o), .n318(n318), .n4980(n4980), .n9652(n9652), 
            .n319(n319), .n9922(n9922), .\r_SM_Main_2__N_2326[0] (r_SM_Main_2__N_2326[0]), 
            .n320(n320), .n321(n321), .n13530(n13530), .tx2_enable(tx2_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(418[10:77])
    uart_rx rx (.n10166(n10166), .r_Bit_Index({r_Bit_Index_adj_36}), .CLK_c(CLK_c), 
            .rx_data_ready(rx_data_ready), .n10194(n10194), .VCC_net(VCC_net), 
            .r_Clock_Count({Open_47, Open_48, \r_Clock_Count[5]_adj_26 , 
            \r_Clock_Count[4]_adj_27 , \r_Clock_Count[3]_adj_28 , \r_Clock_Count[2]_adj_29 , 
            \r_Clock_Count[1]_adj_30 , \r_Clock_Count[0]_adj_25 }), .n10170(n10170), 
            .rx_data({rx_data}), .n10628(n10628), .n10095(n10095), .n10092(n10092), 
            .n10089(n10089), .n10086(n10086), .n10083(n10083), .n10643(n10643), 
            .n10644(n10644), .n10645(n10645), .n10646(n10646), .n3(n3_adj_31), 
            .GND_net(GND_net), .n4(n4_adj_32), .n13597(n13597), .r_Rx_Data(r_Rx_Data), 
            .rx_i(rx_i), .n4_adj_1(n4_adj_33), .n4958(n4958), .n13880(n13880), 
            .n4_adj_2(n4_adj_34), .n9933(n9933), .n8567(n8567), .n8562(n8562), 
            .n9646(n9646), .n221(n221), .n222(n222), .n223(n223), .n224(n224), 
            .n225(n225), .n9920(n9920), .n226(n226), .n9942(n9942), 
            .n9941(n9941), .n9940(n9940)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(380[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_SM_Main, CLK_N_keep, n10638, r_Tx_Data, r_Clock_Count, 
            GND_net, n16998, n18103, n17366, n10637, n10636, n10635, 
            n10634, n10633, n10632, n18102, n17054, r_Bit_Index, 
            n16932, VCC_net, n16954, n16968, n17078, n18101, n17028, 
            n7364, n18104, n9972, n10702, n17084, n17082, n17080, 
            n17030, \r_SM_Main_2__N_2323[1] , n18098, \r_SM_Main_2__N_2326[0] , 
            n4, n8517, n12, n9390, n16466, n10326, n10325, n10324, 
            tx_active, n10323, tx_o, n7086, n7734, tx_enable, n13601, 
            n1, n3, n17757, n7080, n9796, n17950, n17356, n17952, 
            n18010, n18054, n18097) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    input CLK_N_keep;
    input n10638;
    output [7:0]r_Tx_Data;
    output [8:0]r_Clock_Count;
    input GND_net;
    input n16998;
    output n18103;
    input n17366;
    input n10637;
    input n10636;
    input n10635;
    input n10634;
    input n10633;
    input n10632;
    output n18102;
    input n17054;
    output [2:0]r_Bit_Index;
    input n16932;
    input VCC_net;
    input n16954;
    input n16968;
    input n17078;
    output n18101;
    input n17028;
    output n7364;
    output n18104;
    input n9972;
    input n10702;
    input n17084;
    input n17082;
    input n17080;
    input n17030;
    output \r_SM_Main_2__N_2323[1] ;
    output n18098;
    input \r_SM_Main_2__N_2326[0] ;
    output n4;
    output n8517;
    output n12;
    output n9390;
    output n16466;
    input n10326;
    input n10325;
    input n10324;
    output tx_active;
    input n10323;
    output tx_o;
    output n7086;
    output n7734;
    output tx_enable;
    output n13601;
    input n1;
    output n3;
    output n17757;
    output n7080;
    output n9796;
    output n17950;
    input n17356;
    output n17952;
    output n18010;
    output n18054;
    output n18097;
    
    
    wire n10639, n16360, n16361, n16359, n16358, n16357, n17, 
        n10, n17374, n16364, n16363, n16362;
    
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_N_keep), .D(n10639));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_N_keep), .D(n10638));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_6 (.CI(n16360), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n16361));
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_N_keep), .D(n16998));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_5_lut (.I0(n17366), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n16359), .O(n18103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_5 (.CI(n16359), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n16360));
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_N_keep), .D(n10637));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_N_keep), .D(n10636));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_N_keep), .D(n10635));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_N_keep), .D(n10634));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_N_keep), .D(n10633));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_N_keep), .D(n10632));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_4_lut (.I0(n17366), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n16358), .O(n18102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_4 (.CI(n16358), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n16359));
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_N_keep), .D(n17054));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(CLK_N_keep), .E(VCC_net), 
            .D(n16932));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_N_keep), .E(VCC_net), 
            .D(n16954));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_N_keep), .E(VCC_net), 
            .D(n16968));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_N_keep), .E(VCC_net), 
            .D(n17078));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_3_lut (.I0(n17366), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n16357), .O(n18101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'h8228;
    SB_DFFE r_Tx_Done_44 (.Q(n7364), .C(CLK_N_keep), .E(VCC_net), .D(n17028));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_3 (.CI(n16357), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n16358));
    SB_LUT4 add_59_2_lut (.I0(n17366), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n18104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n16357));
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_N_keep), .D(n9972));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_N_keep), .D(n10702));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_N_keep), .D(n17084));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_N_keep), .D(n17082));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n17));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_N_keep), .D(n17080));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_N_keep), .D(n17030));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i15809_2_lut_3_lut (.I0(\r_SM_Main_2__N_2323[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n18098));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i15809_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15852_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_2323[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_2326[0] ), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i15852_3_lut_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8517));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8223_3_lut_4_lut (.I0(\r_SM_Main_2__N_2323[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n10639));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8223_3_lut_4_lut.LUT_INIT = 16'h0078;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[8]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n12));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_2_lut_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[8]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n9390));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_826 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[8]), 
            .I2(r_Clock_Count[6]), .I3(n16466), .O(\r_SM_Main_2__N_2323[1] ));
    defparam i1_2_lut_4_lut_adj_826.LUT_INIT = 16'hfffe;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_N_keep), .D(n10326));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_N_keep), .D(n10325));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_N_keep), .D(n10324));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(CLK_N_keep), .D(n10323));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i4723_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7086));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i4723_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_2326[0] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n7734));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11216_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n13601));
    defparam i11216_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(n1), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[2]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15308_4_lut (.I0(\r_SM_Main_2__N_2323[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n17757));
    defparam i15308_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n16466));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4717_4_lut (.I0(\r_SM_Main_2__N_2326[0] ), .I1(n17), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2323[1] ), .O(n7080));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i4717_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_2323[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n17374));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i7381_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(r_SM_Main[1]), .O(n9796));
    defparam i7381_2_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 add_59_10_lut (.I0(n17356), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n16364), .O(n17950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_59_9_lut (.I0(n17356), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n16363), .O(n17952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_9 (.CI(n16363), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n16364));
    SB_LUT4 add_59_8_lut (.I0(n17356), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n16362), .O(n18010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_8 (.CI(n16362), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n16363));
    SB_LUT4 add_59_7_lut (.I0(n17366), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n16361), .O(n18054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_7 (.CI(n16361), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n16362));
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_N_keep), .D(n17374));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_6_lut (.I0(n17366), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n16360), .O(n18097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    
endmodule
//
// Verilog Description of module uart_tx_U0
//

module uart_tx_U0 (n10245, VCC_net, r_Clock_Count, CLK_c, r_Bit_Index, 
            n10625, n10346, n10008, \r_Clock_Count[5] , n10002, \r_Clock_Count[4] , 
            n9999, \r_Clock_Count[3] , n9996, \r_Clock_Count[2] , n9992, 
            \r_Clock_Count[1] , tx2_data, n10160, \r_SM_Main[2] , GND_net, 
            n10244, n316, n317, tx2_o, n318, n4980, n9652, n319, 
            n9922, \r_SM_Main_2__N_2326[0] , n320, n321, n13530, tx2_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n10245;
    input VCC_net;
    output [8:0]r_Clock_Count;
    input CLK_c;
    output [2:0]r_Bit_Index;
    input n10625;
    input n10346;
    input n10008;
    output \r_Clock_Count[5] ;
    input n10002;
    output \r_Clock_Count[4] ;
    input n9999;
    output \r_Clock_Count[3] ;
    input n9996;
    output \r_Clock_Count[2] ;
    input n9992;
    output \r_Clock_Count[1] ;
    input [7:0]tx2_data;
    input n10160;
    output \r_SM_Main[2] ;
    input GND_net;
    output n10244;
    output n316;
    output n317;
    output tx2_o;
    output n318;
    output n4980;
    output n9652;
    output n319;
    output n9922;
    input \r_SM_Main_2__N_2326[0] ;
    output n320;
    output n321;
    output n13530;
    output tx2_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n18450, n18453, n10656;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n16938;
    wire [8:0]r_Clock_Count_c;   // verilog/uart_tx.v(32[16:29])
    
    wire n16962, n16958, n7727, n18013, n17953, n17939, n10, n16452, 
        n16379, n16378;
    wire [2:0]r_SM_Main_2__N_2323;
    
    wire n16377, n16376, n16375, n23, n16454, n17052, n10331, 
        tx2_active, n10329, n16374, n6812, n16373, n18612, n4, 
        n17990, n18615, n16372, o_Tx_Serial_N_2354, n12306, n9568, 
        n12;
    
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(VCC_net), 
            .D(n10245));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_16115 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n18450));
    defparam r_Bit_Index_0__bdd_4_lut_16115.LUT_INIT = 16'he4aa;
    SB_LUT4 n18450_bdd_4_lut (.I0(n18450), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n18453));
    defparam n18450_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(VCC_net), 
            .D(n10625));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n10346));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n10656));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count_c[8]), .C(CLK_c), .D(n16938));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count_c[7]), .C(CLK_c), .D(n16962));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count_c[6]), .C(CLK_c), .D(n16958));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(\r_Clock_Count[5] ), .C(CLK_c), .D(n10008));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(\r_Clock_Count[4] ), .C(CLK_c), .D(n10002));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(\r_Clock_Count[3] ), .C(CLK_c), .D(n9999));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(\r_Clock_Count[2] ), .C(CLK_c), .D(n9996));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(\r_Clock_Count[1] ), .C(CLK_c), .D(n9992));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n7727), .D(tx2_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10160));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i17_3_lut (.I0(r_Clock_Count_c[6]), .I1(n18013), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n16958));
    defparam i17_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17_3_lut_adj_822 (.I0(r_Clock_Count_c[7]), .I1(n17953), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n16962));
    defparam i17_3_lut_adj_822.LUT_INIT = 16'hacac;
    SB_LUT4 i28_3_lut (.I0(r_Clock_Count_c[8]), .I1(n17939), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n16938));
    defparam i28_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(\r_Clock_Count[3] ), .I1(\r_Clock_Count[2] ), 
            .I2(r_Clock_Count[0]), .I3(\r_Clock_Count[4] ), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(\r_Clock_Count[1] ), .I1(n10), .I2(\r_Clock_Count[5] ), 
            .I3(GND_net), .O(n16452));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_59_10_lut (.I0(n10244), .I1(r_Clock_Count_c[8]), .I2(GND_net), 
            .I3(n16379), .O(n17939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_59_9_lut (.I0(n10244), .I1(r_Clock_Count_c[7]), .I2(GND_net), 
            .I3(n16378), .O(n17953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut (.I0(r_Clock_Count_c[8]), .I1(r_Clock_Count_c[7]), 
            .I2(n16452), .I3(r_Clock_Count_c[6]), .O(r_SM_Main_2__N_2323[1]));   // verilog/uart_tx.v(32[16:29])
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_59_9 (.CI(n16378), .I0(r_Clock_Count_c[7]), .I1(GND_net), 
            .CO(n16379));
    SB_LUT4 add_59_8_lut (.I0(n10244), .I1(r_Clock_Count_c[6]), .I2(GND_net), 
            .I3(n16377), .O(n18013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_8 (.CI(n16377), .I0(r_Clock_Count_c[6]), .I1(GND_net), 
            .CO(n16378));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(\r_Clock_Count[5] ), .I2(GND_net), 
            .I3(n16376), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n16376), .I0(\r_Clock_Count[5] ), .I1(GND_net), 
            .CO(n16377));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(\r_Clock_Count[4] ), .I2(GND_net), 
            .I3(n16375), .O(n317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n16375), .I0(\r_Clock_Count[4] ), .I1(GND_net), 
            .CO(n16376));
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2323[1]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(CLK_c), .D(n16454));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n17052));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx2_active), .C(CLK_c), .D(n10331));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx2_o), .C(CLK_c), .D(n10329));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(\r_Clock_Count[3] ), .I2(GND_net), 
            .I3(n16374), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n16374), .I0(\r_Clock_Count[3] ), .I1(GND_net), 
            .CO(n16375));
    SB_LUT4 i2450_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4980));   // verilog/uart_tx.v(98[36:51])
    defparam i2450_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n7727), .D(tx2_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n7727), .D(tx2_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n7727), .D(tx2_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n7727), .D(tx2_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n7727), .D(tx2_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n7727), .D(tx2_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n7727), .D(tx2_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_2323[1]), .O(n10244));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hccfe;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_2323[1]), .O(n16454));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i4452_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6812));   // verilog/uart_tx.v(96[21:36])
    defparam i4452_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_823 (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_2323[1]), .O(n9652));
    defparam i2_4_lut_adj_823.LUT_INIT = 16'h1101;
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(\r_Clock_Count[2] ), .I2(GND_net), 
            .I3(n16373), .O(n319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7506_4_lut (.I0(n9652), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(n6812), .O(n9922));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i7506_4_lut.LUT_INIT = 16'h8a0a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n18612));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_824 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2326[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_824.LUT_INIT = 16'h4444;
    SB_LUT4 i15730_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_SM_Main_2__N_2323[1]), .I3(GND_net), .O(n17990));   // verilog/uart_tx.v(33[16:27])
    defparam i15730_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n18612_bdd_4_lut (.I0(n18612), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n18615));
    defparam n18612_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_2326[0] ), 
            .I3(\r_SM_Main[2] ), .O(n7727));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_CARRY add_59_4 (.CI(n16373), .I0(\r_Clock_Count[2] ), .I1(GND_net), 
            .CO(n16374));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(\r_Clock_Count[1] ), .I2(GND_net), 
            .I3(n16372), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n16372), .I0(\r_Clock_Count[1] ), .I1(GND_net), 
            .CO(n16373));
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n16372));
    SB_LUT4 i11588211_i1_3_lut (.I0(n18615), .I1(n18453), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_2354));
    defparam i11588211_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9901_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2354), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12306));   // verilog/uart_tx.v(31[16:25])
    defparam i9901_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i9902_3_lut (.I0(tx2_o), .I1(n12306), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n10329));
    defparam i9902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_2323[1]), 
            .I3(r_SM_Main[1]), .O(n10656));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n4), .I2(n23), .I3(r_SM_Main[1]), 
            .O(n9568));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i9913_3_lut (.I0(n9568), .I1(r_SM_Main[1]), .I2(tx2_active), 
            .I3(GND_net), .O(n10331));   // verilog/uart_tx.v(31[16:25])
    defparam i9913_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i29_4_lut (.I0(\r_SM_Main_2__N_2326[0] ), .I1(n17990), .I2(r_SM_Main[1]), 
            .I3(r_Bit_Index[0]), .O(n12));   // verilog/uart_tx.v(33[16:27])
    defparam i29_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_825 (.I0(\r_SM_Main[2] ), .I1(n12), .I2(r_SM_Main_2__N_2323[1]), 
            .I3(r_SM_Main[0]), .O(n17052));   // verilog/uart_tx.v(33[16:27])
    defparam i1_4_lut_adj_825.LUT_INIT = 16'h0544;
    SB_LUT4 i11145_2_lut (.I0(tx2_active), .I1(\r_SM_Main_2__N_2326[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n13530));
    defparam i11145_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx2_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx2_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n10166, r_Bit_Index, CLK_c, rx_data_ready, n10194, 
            VCC_net, r_Clock_Count, n10170, rx_data, n10628, n10095, 
            n10092, n10089, n10086, n10083, n10643, n10644, n10645, 
            n10646, n3, GND_net, n4, n13597, r_Rx_Data, rx_i, 
            n4_adj_1, n4958, n13880, n4_adj_2, n9933, n8567, n8562, 
            n9646, n221, n222, n223, n224, n225, n9920, n226, 
            n9942, n9941, n9940) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n10166;
    output [2:0]r_Bit_Index;
    input CLK_c;
    output rx_data_ready;
    input n10194;
    input VCC_net;
    output [7:0]r_Clock_Count;
    input n10170;
    output [7:0]rx_data;
    input n10628;
    input n10095;
    input n10092;
    input n10089;
    input n10086;
    input n10083;
    input n10643;
    input n10644;
    input n10645;
    input n10646;
    output n3;
    input GND_net;
    output n4;
    output n13597;
    output r_Rx_Data;
    input rx_i;
    output n4_adj_1;
    output n4958;
    output n13880;
    output n4_adj_2;
    input n9933;
    output n8567;
    output n8562;
    output n9646;
    output n221;
    output n222;
    output n223;
    output n224;
    output n225;
    output n9920;
    output n226;
    input n9942;
    input n9941;
    input n9940;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_SM_Main_2__N_2380;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n17351, n16974, n10640, n10301;
    wire [7:0]r_Clock_Count_c;   // verilog/uart_rx.v(32[17:30])
    
    wire n17999, n79, n18066, r_Rx_Data_R, n18001, n10362, n10327, 
        n124, n97, n112, n17376, n10193, n18000, n17381, n13537;
    wire [2:0]r_SM_Main_2__N_2386;
    
    wire n17345, n2, n4_adj_2424, n18003, n16371, n16370, n18594, 
        n18597, n16369, n16368, n16367, n16366, n16365, n9553;
    
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10166));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(r_SM_Main_2__N_2380[2]), 
            .R(n17351));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n16974));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(VCC_net), 
            .D(n10194));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n10170));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(VCC_net), 
            .D(n10628));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n10095));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n10092));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n10089));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n10086));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n10083));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n10640));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(VCC_net), 
            .D(n10643));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n10644));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n10645));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n10646));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count_c[7]), .C(CLK_c), .D(n10301));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i9505_3_lut (.I0(r_Clock_Count_c[7]), .I1(n17999), .I2(n3), 
            .I3(GND_net), .O(n10301));
    defparam i9505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 equal_100_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_100_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i11212_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13597));
    defparam i11212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2380[2]), .I2(GND_net), 
            .I3(GND_net), .O(n79));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n18066), .I2(n79), .I3(r_SM_Main[1]), 
            .O(n10640));   // verilog/uart_rx.v(41[10] 45[8])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(rx_i));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i9493_3_lut (.I0(r_Clock_Count_c[6]), .I1(n18001), .I2(n3), 
            .I3(GND_net), .O(n10362));
    defparam i9493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 equal_102_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_102_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count_c[6]), .C(CLK_c), .D(n10362));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n10327));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2428_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4958));   // verilog/uart_rx.v(102[36:51])
    defparam i2428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n124));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_813 (.I0(r_Clock_Count[3]), .I1(n124), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(n97));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_3_lut_adj_813.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_814 (.I0(r_Clock_Count_c[6]), .I1(r_Clock_Count_c[7]), 
            .I2(GND_net), .I3(GND_net), .O(n112));
    defparam i1_2_lut_adj_814.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_815 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17376));   // verilog/uart_rx.v(36[17:26])
    defparam i1_2_lut_adj_815.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7678_1_lut (.I0(n13880), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n10193));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i7678_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15739_2_lut_3_lut_4_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[0]), .I3(r_SM_Main_2__N_2380[2]), .O(n18000));
    defparam i15739_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 equal_104_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_104_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n9933));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_adj_816 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n17381));   // verilog/uart_rx.v(36[17:26])
    defparam i1_2_lut_adj_816.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_4_lut (.I0(n13537), .I1(n112), .I2(n124), .I3(r_Clock_Count[5]), 
            .O(r_SM_Main_2__N_2386[0]));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i11152_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n13537));
    defparam i11152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_817 (.I0(n97), .I1(r_Clock_Count_c[6]), .I2(r_Clock_Count_c[7]), 
            .I3(r_Clock_Count[5]), .O(n17345));
    defparam i1_4_lut_adj_817.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_818 (.I0(r_SM_Main[2]), .I1(n2), .I2(n17345), 
            .I3(n17376), .O(n4_adj_2424));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_818.LUT_INIT = 16'h1110;
    SB_LUT4 i1_2_lut_adj_819 (.I0(r_SM_Main[2]), .I1(n2), .I2(GND_net), 
            .I3(GND_net), .O(n3));
    defparam i1_2_lut_adj_819.LUT_INIT = 16'heeee;
    SB_LUT4 i15740_4_lut (.I0(n4_adj_2424), .I1(n124), .I2(r_Clock_Count[5]), 
            .I3(n13537), .O(n18003));   // verilog/uart_rx.v(36[17:26])
    defparam i15740_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i57_4_lut (.I0(n18003), .I1(n4_adj_2424), .I2(n17381), .I3(n112), 
            .O(n13880));   // verilog/uart_rx.v(36[17:26])
    defparam i57_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15793_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2386[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n18066));
    defparam i15793_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2386[0]), 
            .I2(r_Rx_Data), .I3(r_SM_Main[1]), .O(n2));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 add_62_9_lut (.I0(n10193), .I1(r_Clock_Count_c[7]), .I2(GND_net), 
            .I3(n16371), .O(n17999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n10193), .I1(r_Clock_Count_c[6]), .I2(GND_net), 
            .I3(n16370), .O(n18001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut (.I0(n17381), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_2380[2]), 
            .I3(r_Bit_Index[0]), .O(n8567));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_4_lut_adj_820 (.I0(n17381), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_2380[2]), 
            .I3(r_Bit_Index[0]), .O(n8562));
    defparam i1_2_lut_4_lut_adj_820.LUT_INIT = 16'hffef;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(r_SM_Main_2__N_2380[2]), .I1(r_SM_Main[1]), 
            .I2(n18000), .I3(r_SM_Main[0]), .O(n18594));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 n18594_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_2386[0]), 
            .I3(n18594), .O(n18597));   // verilog/uart_rx.v(41[10] 45[8])
    defparam n18594_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i1_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_2380[2]), 
            .I3(r_SM_Main[1]), .O(n9646));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h1011;
    SB_LUT4 i130_3_lut_4_lut (.I0(r_Clock_Count_c[6]), .I1(r_Clock_Count_c[7]), 
            .I2(n97), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_2380[2]));   // verilog/uart_rx.v(32[17:30])
    defparam i130_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_adj_821 (.I0(r_SM_Main[2]), .I1(n18597), .I2(GND_net), 
            .I3(GND_net), .O(n10327));
    defparam i1_2_lut_adj_821.LUT_INIT = 16'h4444;
    SB_CARRY add_62_8 (.CI(n16370), .I0(r_Clock_Count_c[6]), .I1(GND_net), 
            .CO(n16371));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n16369), .O(n221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n16369), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n16370));
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n16368), .O(n222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_6 (.CI(n16368), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n16369));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n16367), .O(n223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n16367), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n16368));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n16366), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n16366), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n16367));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n16365), .O(n225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7504_3_lut_4_lut (.I0(r_Bit_Index[2]), .I1(n4958), .I2(r_SM_Main[1]), 
            .I3(n9646), .O(n9920));
    defparam i7504_3_lut_4_lut.LUT_INIT = 16'h8f00;
    SB_CARRY add_62_3 (.CI(n16365), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n16366));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n16365));
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_2380[2]), 
            .I3(r_SM_Main[0]), .O(n9553));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h4033;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n9553), 
            .I3(rx_data_ready), .O(n16974));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i15891_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n17351));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15891_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n9942));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n9941));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n9940));   // verilog/uart_rx.v(49[10] 144[8])
    
endmodule
